module in01s01 ();
  output o;
  input a;
endmodule

module in01s02 ();
  output o;
  input a;
endmodule

module in01s03 ();
  output o;
  input a;
endmodule

module in01s04 ();
  output o;
  input a;
endmodule

module in01s06 ();
  output o;
  input a;
endmodule

module in01s08 ();
  output o;
  input a;
endmodule

module in01s10 ();
  output o;
  input a;
endmodule

module in01s20 ();
  output o;
  input a;
endmodule

module in01s40 ();
  output o;
  input a;
endmodule

module in01s80 ();
  output o;
  input a;
endmodule

module in01m01 ();
  output o;
  input a;
endmodule

module in01m02 ();
  output o;
  input a;
endmodule

module in01m03 ();
  output o;
  input a;
endmodule

module in01m04 ();
  output o;
  input a;
endmodule

module in01m06 ();
  output o;
  input a;
endmodule

module in01m08 ();
  output o;
  input a;
endmodule

module in01m10 ();
  output o;
  input a;
endmodule

module in01m20 ();
  output o;
  input a;
endmodule

module in01m40 ();
  output o;
  input a;
endmodule

module in01m80 ();
  output o;
  input a;
endmodule

module in01f01 ();
  output o;
  input a;
endmodule

module in01f02 ();
  output o;
  input a;
endmodule

module in01f03 ();
  output o;
  input a;
endmodule

module in01f04 ();
  output o;
  input a;
endmodule

module in01f06 ();
  output o;
  input a;
endmodule

module in01f08 ();
  output o;
  input a;
endmodule

module in01f10 ();
  output o;
  input a;
endmodule

module in01f20 ();
  output o;
  input a;
endmodule

module in01f40 ();
  output o;
  input a;
endmodule

module in01f80 ();
  output o;
  input a;
endmodule

module na02s01 ();
  output o;
  input a;
  input b;
endmodule

module na02s02 ();
  output o;
  input a;
  input b;
endmodule

module na02s03 ();
  output o;
  input a;
  input b;
endmodule

module na02s04 ();
  output o;
  input a;
  input b;
endmodule

module na02s06 ();
  output o;
  input a;
  input b;
endmodule

module na02s08 ();
  output o;
  input a;
  input b;
endmodule

module na02s10 ();
  output o;
  input a;
  input b;
endmodule

module na02s20 ();
  output o;
  input a;
  input b;
endmodule

module na02s40 ();
  output o;
  input a;
  input b;
endmodule

module na02s80 ();
  output o;
  input a;
  input b;
endmodule

module na02m01 ();
  output o;
  input a;
  input b;
endmodule

module na02m02 ();
  output o;
  input a;
  input b;
endmodule

module na02m03 ();
  output o;
  input a;
  input b;
endmodule

module na02m04 ();
  output o;
  input a;
  input b;
endmodule

module na02m06 ();
  output o;
  input a;
  input b;
endmodule

module na02m08 ();
  output o;
  input a;
  input b;
endmodule

module na02m10 ();
  output o;
  input a;
  input b;
endmodule

module na02m20 ();
  output o;
  input a;
  input b;
endmodule

module na02m40 ();
  output o;
  input a;
  input b;
endmodule

module na02m80 ();
  output o;
  input a;
  input b;
endmodule

module na02f01 ();
  output o;
  input a;
  input b;
endmodule

module na02f02 ();
  output o;
  input a;
  input b;
endmodule

module na02f03 ();
  output o;
  input a;
  input b;
endmodule

module na02f04 ();
  output o;
  input a;
  input b;
endmodule

module na02f06 ();
  output o;
  input a;
  input b;
endmodule

module na02f08 ();
  output o;
  input a;
  input b;
endmodule

module na02f10 ();
  output o;
  input a;
  input b;
endmodule

module na02f20 ();
  output o;
  input a;
  input b;
endmodule

module na02f40 ();
  output o;
  input a;
  input b;
endmodule

module na02f80 ();
  output o;
  input a;
  input b;
endmodule

module na03s01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03s80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03m80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na03f80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module na04s01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04s80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04m80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module na04f80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no02s01 ();
  output o;
  input a;
  input b;
endmodule

module no02s02 ();
  output o;
  input a;
  input b;
endmodule

module no02s03 ();
  output o;
  input a;
  input b;
endmodule

module no02s04 ();
  output o;
  input a;
  input b;
endmodule

module no02s06 ();
  output o;
  input a;
  input b;
endmodule

module no02s08 ();
  output o;
  input a;
  input b;
endmodule

module no02s10 ();
  output o;
  input a;
  input b;
endmodule

module no02s20 ();
  output o;
  input a;
  input b;
endmodule

module no02s40 ();
  output o;
  input a;
  input b;
endmodule

module no02s80 ();
  output o;
  input a;
  input b;
endmodule

module no02m01 ();
  output o;
  input a;
  input b;
endmodule

module no02m02 ();
  output o;
  input a;
  input b;
endmodule

module no02m03 ();
  output o;
  input a;
  input b;
endmodule

module no02m04 ();
  output o;
  input a;
  input b;
endmodule

module no02m06 ();
  output o;
  input a;
  input b;
endmodule

module no02m08 ();
  output o;
  input a;
  input b;
endmodule

module no02m10 ();
  output o;
  input a;
  input b;
endmodule

module no02m20 ();
  output o;
  input a;
  input b;
endmodule

module no02m40 ();
  output o;
  input a;
  input b;
endmodule

module no02m80 ();
  output o;
  input a;
  input b;
endmodule

module no02f01 ();
  output o;
  input a;
  input b;
endmodule

module no02f02 ();
  output o;
  input a;
  input b;
endmodule

module no02f03 ();
  output o;
  input a;
  input b;
endmodule

module no02f04 ();
  output o;
  input a;
  input b;
endmodule

module no02f06 ();
  output o;
  input a;
  input b;
endmodule

module no02f08 ();
  output o;
  input a;
  input b;
endmodule

module no02f10 ();
  output o;
  input a;
  input b;
endmodule

module no02f20 ();
  output o;
  input a;
  input b;
endmodule

module no02f40 ();
  output o;
  input a;
  input b;
endmodule

module no02f80 ();
  output o;
  input a;
  input b;
endmodule

module no03s01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03s80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03m80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no03f80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module no04s01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04s80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04m80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module no04f80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao12s01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12s80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12m80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao12f80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module ao22s01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22s80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22m80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ao22f80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa12s01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12s80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12m80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f01 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f02 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f03 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f04 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f06 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f08 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa12f80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module oa22s01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22s80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22m80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f01 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f02 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f03 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f04 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f06 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f08 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module oa22f80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module ms00f10 ();
  input ck;
  input d;
  output q;
endmodule

module ms00f20 ();
  input ck;
  input d;
  output q;
endmodule

module ms00f40 ();
  input ck;
  input d;
  output q;
endmodule

module ms00f80 ();
  output o;
  input ck;
  input d;
endmodule

