`include <inter.v>

module top;

// Start PIs
input PI_AD_2;
input PI_AD_12;
input PI_AD_37;
input PI_AD_9;
input PI_AD_26;
input PI_AD_54;
input PI_AD_48;
input PI_AD_31;
input PI_AD_17;
input PI_AD_18;
input PI_AD_29;
input PI_AD_11;
input PI_FRAME_L;
input PI_AD_24;
input PI_AD_40;
input PI_AD_62;
input PI_AD_30;
input PI_AD_25;
input PI_CBE_L_4;
input PI_AD_46;
input PI_REQ64_L;
input PI_AD_6;
input PI_AD_19;
input PI_AD_47;
input PI_AD_59;
input PI_AD_60;
input PI_AD_32;
input PI_AD_3;
input PI_AD_1;
input PI_CBE_L_6;
input PI_AD_39;
input PI_AD_27;
input PI_AD_15;
input PI_AD_43;
input PI_PAR;
input PI_AD_42;
input PI_CBE_L_2;
input PI_AD_7;
input PI_AD_61;
input PI_AD_36;
input PI_CBE_L_7;
input PI_AD_16;
input PI_CBE_L_5;
input PI_AD_0;
input PI_AD_22;
input PI_PAR64;
input PI_AD_35;
input PI_AD_34;
input PI_IDSEL;
input PI_CBE_L_0;
input PI_AD_56;
input PI_AD_45;
input PI_AD_21;
input tau_clk;
input PI_AD_51;
input PI_CBE_L_3;
input PI_AD_10;
input PI_AD_52;
input PI_AD_5;
input PI_AD_23;
input PI_AD_63;
input PI_AD_20;
input PI_AD_13;
input PI_AD_55;
input PI_AD_58;
input PI_AD_4;
input PI_AD_28;
input PI_AD_38;
input PI_AD_33;
input PI_AD_41;
input PI_AD_44;
input PI_AD_8;
input PI_IRDY_L;
input PI_AD_50;
input PI_CBE_L_1;
input RESET;
input PI_AD_57;
input PI_AD_53;
input PI_AD_49;
input PI_AD_14;

// Start POs
output PO_AD_35;
output PO_AD_40;
output PO_AD_8;
output PO_AD_15;
output PO_AD_21;
output PO_AD_59;
output PO_AD_53;
output PO_AD_24;
output PO_PAR;
output PO_AD_52;
output PO_AD_9;
output PO_AD_57;
output PO_AD_48;
output PO_AD_14;
output PO_AD_39;
output PO_STOP_L;
output PO_AD_28;
output PO_AD_25;
output PO_AD_22;
output PO_AD_63;
output PO_AD_38;
output PO_AD_42;
output PO_AD_7;
output PO_AD_4;
output PO_PAR64;
output PO_AD_43;
output PO_AD_2;
output PO_AD_62;
output TAR_TRI_S;
output PO_AD_5;
output TAR_TRI_A;
output PO_AD_3;
output PO_AD_6;
output PO_AD_12;
output PO_AD_13;
output PO_AD_41;
output PO_ACK64_L;
output PO_TRDY_L;
output PO_AD_33;
output PO_AD_23;
output PO_AD_16;
output PO_AD_18;
output PO_AD_32;
output PO_AD_50;
output PO_AD_26;
output TAR_TRI_D;
output PO_AD_55;
output TAR_TRI_E;
output PO_SERR_L;
output TAR_TRI_T;
output PO_AD_54;
output PO_AD_49;
output PO_PERR_L;
output PO_AD_31;
output TAR_TRI_P;
output PO_AD_36;
output PO_AD_51;
output PO_DEVSEL_L;
output PO_AD_0;
output PO_AD_1;
output PO_AD_10;
output PO_AD_29;
output PO_AD_17;
output PO_AD_56;
output PO_AD_58;
output PO_AD_45;
output PO_AD_11;
output PO_AD_30;
output PO_AD_46;
output PO_AD_47;
output PO_AD_60;
output PO_AD_20;
output PO_AD_44;
output PO_AD_61;
output PO_AD_37;
output PO_AD_34;
output PO_AD_27;
output PO_AD_19;

// Start wires
wire n_356;
wire newNet_199;
wire n_707;
wire newNet_235;
wire cordic_Add0_MUX_0_n_14;
wire PO_AD_40;
wire newNet_10;
wire cordic_SH1_srl_35_26_n_73;
wire newNet_166;
wire cordic_SH2_srl_35_26_n_127;
wire cordic_AddX_MUX_1_n_17;
wire n_192;
wire n_685;
wire newNet_451;
wire n_75;
wire cordic_SH2_srl_35_26_n_33;
wire newNet_73;
wire cordic_Add0_MUX_0_n_16;
wire newNet_828;
wire newNet_342;
wire n_61;
wire n_502;
wire cordic_AddY_Atemp_15_;
wire n_98;
wire newNet_1073;
wire cordic_Add0_Compl_n_12;
wire cordic_AddX_MUX_1_n_18;
wire cordic_AddX_MUX_0_n_22;
wire n_750;
wire cordic_SH1_srl_35_26_n_109;
wire cordic_AddX_Atemp_14_;
wire n_89;
wire newNet_862;
wire n_868;
wire n_25;
wire cordic_AddX_MUX_1_n_28;
wire cordic_iteration_3_;
wire n_701;
wire cordic_n_119;
wire cordic_AddY_Compl_n_15;
wire n_861;
wire newNet_83;
wire CoreOutputReg_20_;
wire System_Busy;
wire n_410;
wire cordic_iteration_1_;
wire n_114;
wire newNet_857;
wire newNet_623;
wire newNet_562;
wire newNet_731;
wire cordic_AddX_Atemp_11_;
wire n_1047;
wire cordic_n_19;
wire n_274;
wire PI_AD_16;
wire newNet_780;
wire newNet_575;
wire cordic_AddX_Stemp_7_;
wire n_326;
wire newNet_353;
wire n_1062;
wire cordic_SH2_srl_35_26_n_22;
wire newNet_1178;
wire n_682;
wire newNet_774;
wire newNet_546;
wire Core_Cnt_2_;
wire n_373;
wire cordic_AddX_Add_n_29;
wire cordic_AddX_Add_n_6;
wire newNet_727;
wire newNet_92;
wire cordic_AddY_MUX_1_n_29;
wire newNet_19;
wire n_68;
wire newNet_769;
wire n_601;
wire cordic_SH1_srl_35_26_n_38;
wire newNet_1199;
wire cordic_AddX_Add_n_15;
wire cordic_AddY_Compl_n_31;
wire newNet_995;
wire newNet_662;
wire newNet_1162;
wire newNet_1084;
wire cordic_AddY_Stemp_13_;
wire n_736;
wire newNet_674;
wire n_811;
wire n_629;
wire newNet_961;
wire newNet_433;
wire newNet_183;
wire n_249;
wire cordic_pla_n_19;
wire newNet_256;
wire cordic_X_15_;
wire n_332;
wire newNet_99;
wire cordic_SH2_srl_35_26_n_63;
wire n_165;
wire newNet_237;
wire newNet_1202;
wire newNet_346;
wire n_363;
wire cordic_AddX_Stemp_3_;
wire cordic_AddX_Atemp_10_;
wire State_0_;
wire newNet_339;
wire newNet_268;
wire cordic_AddX_Btemp_7_;
wire newNet_369;
wire newNet_627;
wire newNet_894;
wire newNet_319;
wire newNet_365;
wire cordic_AddX_Btemp_15_;
wire newNet_1110;
wire newNet_817;
wire newNet_689;
wire cordic_AddY_MUX_1_n_12;
wire n_372;
wire n_147;
wire CoreOutput_32_;
wire cordic_SH2_srl_35_26_n_106;
wire cordic_AddX_Add_n_73;
wire cordic_SH2_srl_35_26_n_66;
wire cordic_SH2_srl_35_26_n_111;
wire newNet_761;
wire CoreOutputReg_13_;
wire newNet_883;
wire newNet_927;
wire cordic_AddY_MUX_1_n_19;
wire n_324;
wire newNet_244;
wire n_486;
wire cordic_n_51;
wire n_800;
wire newNet_261;
wire cordic_Add0_Btemp_13_;
wire cordic_n_31;
wire newNet_594;
wire cordic_X_2_;
wire PI_AD_24;
wire cordic_n_53;
wire n_780;
wire newNet_29;
wire cordic_n_44;
wire newNet_1023;
wire newNet_5;
wire PI_AD_60;
wire newNet_660;
wire n_349;
wire cordic_SH2_srl_35_26_n_105;
wire newNet_521;
wire cordic_SH1_srl_35_26_n_104;
wire n_359;
wire newNet_757;
wire cordic_AddY_Add_n_1;
wire newNet_873;
wire newNet_260;
wire n_485;
wire n_44;
wire cordic_AddY_MUX_0_n_8;
wire cordic_Angle_9_;
wire n_222;
wire n_537;
wire n_884;
wire newNet_821;
wire n_796;
wire cordic_Angle_6_;
wire cordic_BS2_10_;
wire n_506;
wire newNet_695;
wire newNet_1013;
wire newNet_848;
wire newNet_271;
wire cordic_AddY_Atemp_11_;
wire cordic_SH2_srl_35_26_n_80;
wire newNet_390;
wire cordic_AddX_Atemp_1_;
wire n_578;
wire newNet_721;
wire cordic_SH2_srl_35_26_n_90;
wire cordic_pla_n_8;
wire n_383;
wire newNet_335;
wire cordic_Add0_Add_n_0;
wire PI_AD_56;
wire n_606;
wire n_158;
wire n_152;
wire CoreOutputReg_19_;
wire newNet_967;
wire newNet_138;
wire newNet_293;
wire newNet_936;
wire newNet_867;
wire n_838;
wire cordic_AddY_Btemp_1_;
wire n_624;
wire cordic_Y_4_;
wire newNet_882;
wire Burst_Trans;
wire newNet_913;
wire n_727;
wire newNet_788;
wire newNet_385;
wire cordic_Add0_MUX_0_n_21;
wire newNet_607;
wire cordic_SH1_srl_35_26_n_22;
wire newNet_504;
wire n_298;
wire newNet_790;
wire newNet_285;
wire newNet_177;
wire cordic_AddY_Btemp_3_;
wire CoreCnt_En;
wire n_296;
wire newNet_1102;
wire cordic_SH2_srl_35_26_n_1;
wire cordic_Add0_MUX_0_n_29;
wire cordic_pla_n_14;
wire cordic_AddY_Add_n_5;
wire cordic_SH1_srl_35_26_n_64;
wire CoreOutputReg_17_;
wire cordic_Add0_MUX_0_n_8;
wire newNet_648;
wire cordic_Add0_Add_n_11;
wire cordic_Add0_Add_n_74;
wire cordic_pla_n_30;
wire newNet_879;
wire newNet_509;
wire newNet_705;
wire cordic_AddX_MUX_0_n_13;
wire newNet_811;
wire newNet_312;
wire n_200;
wire newNet_691;
wire cordic_AddY_Add_n_52;
wire cordic_pla_n_22;
wire cordic_tanangle_9_;
wire CoreOutput_14_;
wire cordic_SH2_srl_35_26_n_97;
wire PO_AD_53;
wire CoreInput_15_;
wire cordic_Add0_Add_n_33;
wire n_334;
wire cordic_Add0_Add_n_5;
wire n_303;
wire cordic_AddY_Add_n_23;
wire n_257;
wire Core_Cnt_1_;
wire cordic_AddY_MUX_1_n_28;
wire cordic_AddX_MUX_1_n_6;
wire cordic_SH1_srl_35_26_n_45;
wire newNet_1004;
wire cordic_BS2_2_;
wire n_35;
wire n_513;
wire newNet_975;
wire cordic_Angle_0_;
wire PI_AD_11;
wire n_718;
wire cordic_AddX_Add_n_26;
wire cordic_Add0_n_16;
wire n_735;
wire newNet_1063;
wire newNet_479;
wire n_2;
wire n_817;
wire cordic_n_8;
wire cordic_Add0_Compl_n_25;
wire cordic_AddY_Add_n_43;
wire cordic_AddY_Add_n_59;
wire n_20;
wire n_621;
wire cordic_Add0_Compl_n_29;
wire n_437;
wire n_431;
wire PO_AD_7;
wire n_104;
wire PI_AD_39;
wire n_477;
wire PI_AD_43;
wire cordic_pla_n_4;
wire newNet_779;
wire newNet_669;
wire newNet_388;
wire n_175;
wire n_531;
wire newNet_485;
wire CoreOutputReg_18_;
wire newNet_878;
wire cordic_SH2_srl_35_26_n_59;
wire newNet_1135;
wire newNet_983;
wire newNet_424;
wire n_692;
wire Trdy_Cnt_En;
wire cordic_AddX_Add_n_12;
wire cordic_AddX_Compl_n_2;
wire cordic_AddY_Btemp1_13_;
wire cordic_Add0_Add_n_48;
wire cordic_Y_8_;
wire n_597;
wire newNet_1175;
wire cordic_Add0_Add_n_14;
wire newNet_1144;
wire newNet_205;
wire newNet_316;
wire cordic_iteration_2_;
wire newNet_588;
wire newNet_743;
wire n_1063;
wire newNet_922;
wire cordic_SH2_srl_35_26_n_7;
wire cordic_AddX_Btemp_8_;
wire n_124;
wire cordic_n_20;
wire n_95;
wire newNet_376;
wire cordic_Add0_Add_n_30;
wire n_658;
wire cordic_AddY_Stemp_9_;
wire n_4;
wire cordic_SH1_srl_35_26_n_111;
wire cordic_n_47;
wire n_552;
wire cordic_AddX_n_0;
wire n_264;
wire cordic_AddX_MUX_1_n_25;
wire cordic_SH2_srl_35_26_n_56;
wire cordic_Add0_Btemp_2_;
wire newNet_591;
wire cordic_AddY_Btemp_11_;
wire newNet_748;
wire Access_Address_1_27_;
wire n_269;
wire n_651;
wire newNet_797;
wire cordic_AddY_Add_n_64;
wire n_9;
wire n_590;
wire Config_Reg_6_;
wire newNet_106;
wire CoreOutput_30_;
wire Core_Cnt_0_;
wire newNet_941;
wire cordic_AddY_Btemp_6_;
wire newNet_899;
wire cordic_SH1_srl_35_26_n_55;
wire newNet_1117;
wire PI_IRDY_L;
wire n_217;
wire n_618;
wire cordic_AddX_MUX_1_n_5;
wire cordic_Add0_MUX_0_n_4;
wire newNet_152;
wire n_57;
wire cordic_SH2_srl_35_26_n_122;
wire cordic_Add0_MUX_1_n_28;
wire cordic_Add0_MUX_0_n_31;
wire n_236;
wire n_743;
wire n_445;
wire newNet_482;
wire newNet_836;
wire n_522;
wire n_587;
wire n_787;
wire n_255;
wire n_639;
wire newNet_35;
wire n_452;
wire newNet_304;
wire cordic_AddY_MUX_1_n_24;
wire cordic_SH1_srl_35_26_n_60;
wire cordic_Add0_Btemp_1_;
wire cordic_Add0_Btemp_5_;
wire cordic_AddX_Btemp_3_;
wire cordic_Y_10_;
wire cordic_SH1_srl_35_26_n_6;
wire newNet_834;
wire cordic_SH1_srl_35_26_n_118;
wire Access_Address_1_25_;
wire newNet_1068;
wire cordic_n_27;
wire newNet_240;
wire newNet_543;
wire n_848;
wire newNet_396;
wire cordic_AddY_Btemp1_15_;
wire n_779;
wire newNet_444;
wire n_78;
wire newNet_902;
wire newNet_1042;
wire newNet_412;
wire newNet_598;
wire cordic_AddY_Atemp_14_;
wire newNet_49;
wire PI_AD_7;
wire newNet_870;
wire CoreInput_8_;
wire cordic_SH2_srl_35_26_n_101;
wire cordic_SH1_srl_35_26_n_98;
wire cordic_n_39;
wire n_28;
wire cordic_X_3_;
wire cordic_AddY_n_0;
wire n_499;
wire n_765;
wire newNet_1190;
wire n_245;
wire newNet_602;
wire newNet_96;
wire n_181;
wire newNet_1040;
wire newNet_1031;
wire cordic_AddY_MUX_0_n_21;
wire cordic_Add0_MUX_1_n_16;
wire newNet_307;
wire cordic_Add0_n_13;
wire cordic_n_75;
wire n_422;
wire newNet_806;
wire n_348;
wire PO_AD_32;
wire newNet_407;
wire newNet_1037;
wire cordic_Add0_MUX_0_n_24;
wire newNet_141;
wire cordic_SH1_srl_35_26_n_29;
wire cordic_SH1_srl_35_26_n_76;
wire newNet_1055;
wire cordic_n_73;
wire cordic_n_26;
wire n_967;
wire cordic_AddY_Stemp_7_;
wire n_419;
wire newNet_356;
wire n_833;
wire newNet_87;
wire cordic_SH1_srl_35_26_n_51;
wire n_666;
wire n_86;
wire cordic_AddY_Atemp_8_;
wire Issue_Rst;
wire cordic_AddY_MUX_0_n_15;
wire cordic_Add0_Atemp_2_;
wire n_496;
wire newNet_202;
wire n_133;
wire newNet_187;
wire Config_Reg_8_;
wire CoreInput_0_;
wire CoreOutput_12_;
wire newNet_1089;
wire newNet_448;
wire newNet_259;
wire n_50;
wire cordic_AddY_MUX_1_n_6;
wire newNet_68;
wire cordic_BS2_9_;
wire cordic_AddY_Compl_n_41;
wire n_131;
wire newNet_134;
wire n_482;
wire newNet_558;
wire cordic_AddY_MUX_1_n_2;
wire n_865;
wire cordic_SH1_srl_35_26_n_5;
wire PO_AD_21;
wire newNet_315;
wire n_722;
wire newNet_678;
wire cordic_Angle_10_;
wire newNet_7;
wire newNet_437;
wire newNet_752;
wire n_814;
wire newNet_526;
wire newNet_243;
wire cordic_Add0_MUX_0_n_7;
wire n_574;
wire n_729;
wire newNet_571;
wire cordic_AddX_Compl_n_43;
wire DevSel_Cnt_En;
wire cordic_AddX_MUX_1_n_14;
wire cordic_Angle_3_;
wire newNet_281;
wire newNet_443;
wire n_188;
wire newNet_637;
wire cordic_Angle_11_;
wire cordic_SH1_srl_35_26_n_67;
wire cordic_Add0_Add_n_22;
wire cordic_n_83;
wire n_843;
wire newNet_145;
wire newNet_1126;
wire n_292;
wire newNet_61;
wire newNet_162;
wire cordic_AddY_Add_n_17;
wire PI_CBE_L_6;
wire newNet_155;
wire cordic_AddY_Add_n_70;
wire n_676;
wire newNet_895;
wire newNet_1065;
wire cordic_n_102;
wire CoreOutputReg_7_;
wire n_471;
wire n_879;
wire n_754;
wire cordic_AddX_MUX_1_n_13;
wire cordic_SumAngle_14_;
wire cordic_Add0_Compl_n_5;
wire n_148;
wire newNet_765;
wire cordic_SH2_srl_35_26_n_26;
wire cordic_n_96;
wire n_474;
wire cordic_Add0_Atemp_3_;
wire cordic_tanangle_1_;
wire newNet_952;
wire n_898;
wire cordic_Add0_MUX_1_n_19;
wire cordic_SH2_srl_35_26_n_73;
wire cordic_Add0_Stemp_8_;
wire cordic_AddX_Y_2;
wire newNet_577;
wire n_74;
wire Access_Address_1_20_;
wire cordic_SH2_srl_35_26_n_126;
wire PI_CBE_L_0;
wire cordic_SH2_srl_35_26_n_19;
wire n_120;
wire n_376;
wire cordic_AddY_Y_1;
wire newNet_276;
wire newNet_95;
wire cordic_Add0_MUX_1_n_8;
wire n_455;
wire n_841;
wire newNet_1120;
wire newNet_784;
wire newNet_766;
wire cordic_Add0_MUX_0_n_25;
wire cordic_n_9;
wire cordic_AddX_MUX_0_n_20;
wire cordic_Add0_MUX_1_n_31;
wire cordic_SH2_srl_35_26_n_132;
wire cordic_Add0_n_10;
wire newNet_805;
wire cordic_AddY_Add_n_44;
wire n_851;
wire cordic_n_70;
wire newNet_459;
wire n_568;
wire newNet_30;
wire cordic_AddX_MUX_0_n_25;
wire newNet_21;
wire newNet_666;
wire cordic_tanangle_3_;
wire cordic_SH1_srl_35_26_n_100;
wire cordic_AddY_Add_n_32;
wire cordic_tanangle_5_;
wire newNet_823;
wire cordic_AddX_Add_n_56;
wire n_193;
wire n_39;
wire cordic_AddY_MUX_1_n_9;
wire cordic_n_35;
wire PO_AD_58;
wire n_201;
wire n_143;
wire cordic_SH1_srl_35_26_n_105;
wire n_377;
wire newNet_195;
wire cordic_AddY_Compl_n_11;
wire cordic_Add0_Atemp_12_;
wire cordic_AddY_Add_n_12;
wire cordic_AddX_MUX_1_n_20;
wire cordic_n_65;
wire cordic_X_8_;
wire newNet_1195;
wire newNet_712;
wire n_71;
wire newNet_123;
wire Access_Address_1_17_;
wire cordic_AddX_Add_n_43;
wire cordic_AddX_Stemp_14_;
wire newNet_249;
wire newNet_324;
wire newNet_222;
wire n_386;
wire newNet_171;
wire newNet_672;
wire cordic_pla_n_10;
wire newNet_963;
wire cordic_AddX_Y_3;
wire newNet_675;
wire newNet_326;
wire n_271;
wire newNet_360;
wire cordic_n_68;
wire cordic_AddX_Add_n_64;
wire cordic_n_16;
wire cordic_Add0_Atemp_6_;
wire newNet_701;
wire newNet_1016;
wire n_65;
wire n_41;
wire newNet_70;
wire newNet_289;
wire cordic_Add0_Atemp_0_;
wire cordic_AddY_Btemp_12_;
wire newNet_476;
wire cordic_SH2_srl_35_26_n_109;
wire n_304;
wire newNet_462;
wire n_100;
wire cordic_AddY_Add_n_68;
wire cordic_n_79;
wire PI_AD_47;
wire n_655;
wire n_719;
wire newNet_428;
wire cordic_Add0_Stemp_4_;
wire cordic_Add0_Add_n_54;
wire newNet_735;
wire cordic_AddY_MUX_0_n_20;
wire n_347;
wire n_620;
wire newNet_251;
wire newNet_886;
wire cordic_n_2;
wire n_793;
wire newNet_1045;
wire newNet_18;
wire n_542;
wire newNet_890;
wire cordic_AddY_Atemp_0_;
wire n_783;
wire newNet_15;
wire n_320;
wire Access_Type_1_1_;
wire newNet_77;
wire cordic_AddX_Btemp1_3_;
wire newNet_34;
wire PAR_Int_d;
wire newNet_530;
wire newNet_687;
wire n_117;
wire newNet_1166;
wire newNet_1155;
wire PO_AD_16;
wire cordic_AddX_Btemp1_0_;
wire newNet_887;
wire newNet_772;
wire cordic_Add0_Add_n_51;
wire n_880;
wire newNet_1096;
wire cordic_Add0_MUX_1_n_12;
wire newNet_655;
wire newNet_290;
wire cordic_AddX_Compl_n_33;
wire cordic_n_93;
wire n_469;
wire newNet_907;
wire newNet_1017;
wire cordic_AddX_MUX_0_n_3;
wire cordic_AddX_MUX_0_n_31;
wire newNet_943;
wire cordic_pla_n_36;
wire n_402;
wire newNet_184;
wire cordic_AddX_Add_n_22;
wire cordic_BS1_12_;
wire cordic_AddY_Compl_n_6;
wire PO_DEVSEL_L;
wire n_834;
wire cordic_Add0_MUX_0_n_13;
wire PI_AD_4;
wire newNet_590;
wire newNet_381;
wire n_615;
wire CoreOutputReg_9_;
wire newNet_849;
wire cordic_SH2_srl_35_26_n_72;
wire n_642;
wire n_48;
wire cordic_SH2_srl_35_26_n_37;
wire cordic_AddX_Add_n_58;
wire n_516;
wire newNet_709;
wire cordic_n_88;
wire n_859;
wire cordic_Add0_Atemp_5_;
wire CoreOutput_10_;
wire cordic_AddY_Compl_n_1;
wire newNet_40;
wire PO_AD_60;
wire n_858;
wire n_367;
wire PO_AD_44;
wire cordic_SH2_srl_35_26_n_91;
wire n_440;
wire newNet_1028;
wire n_204;
wire n_774;
wire n_726;
wire n_481;
wire cordic_SH2_srl_35_26_n_117;
wire n_198;
wire cordic_AddX_Stemp_11_;
wire cordic_AddY_Btemp1_11_;
wire cordic_n_45;
wire n_891;
wire n_226;
wire cordic_SH1_srl_35_26_n_88;
wire n_563;
wire newNet_1139;
wire newNet_632;
wire cordic_SH1_srl_35_26_n_42;
wire cordic_Add0_Atemp_14_;
wire newNet_103;
wire cordic_n_48;
wire cordic_SH1_srl_35_26_n_127;
wire cordic_BS1_10_;
wire n_465;
wire newNet_161;
wire newNet_493;
wire n_230;
wire n_449;
wire cordic_AddX_Add_n_16;
wire cordic_Ysign;
wire newNet_1106;
wire newNet_926;
wire cordic_SH2_srl_35_26_n_49;
wire n_696;
wire n_661;
wire cordic_Add0_Stemp_2_;
wire newNet_844;
wire cordic_AddX_Compl_n_11;
wire PI_AD_15;
wire cordic_Add0_MUX_1_n_20;
wire newNet_1130;
wire cordic_SH1_srl_35_26_n_59;
wire cordic_Angle_1_;
wire cordic_SH1_srl_35_26_n_115;
wire newNet_866;
wire cordic_Add0_MUX_0_n_1;
wire cordic_SumAngle_2_;
wire n_371;
wire newNet_159;
wire PO_AD_3;
wire PI_AD_61;
wire newNet_583;
wire newNet_842;
wire cordic_Angle_7_;
wire PO_AD_13;
wire newNet_1090;
wire newNet_371;
wire DevSel_Wait_Cnt_2_;
wire newNet_471;
wire n_770;
wire n_417;
wire newNet_775;
wire newNet_387;
wire newNet_229;
wire newNet_217;
wire newNet_696;
wire PI_IDSEL;
wire n_673;
wire newNet_947;
wire n_213;
wire newNet_516;
wire cordic_AddX_MUX_0_n_29;
wire n_171;
wire n_649;
wire newNet_875;
wire PO_AD_26;
wire newNet_1058;
wire n_495;
wire cordic_n_6;
wire n_288;
wire n_398;
wire cordic_SH1_srl_35_26_n_10;
wire cordic_Add0_MUX_0_n_19;
wire n_555;
wire newNet_203;
wire TAR_TRI_P;
wire newNet_333;
wire n_29;
wire newNet_127;
wire n_99;
wire PI_AD_28;
wire cordic_Angle_2_;
wire CoreOutputReg_10_;
wire n_706;
wire n_344;
wire cordic_Add0_Compl_n_2;
wire cordic_AddX_MUX_1_n_32;
wire cordic_SH1_srl_35_26_n_17;
wire PO_AD_56;
wire CoreOutputReg_25_;
wire Config_Reg_30_;
wire newNet_1101;
wire cordic_SH1_srl_35_26_n_40;
wire CoreOutput_5_;
wire n_10;
wire newNet_971;
wire n_432;
wire cordic_n_23;
wire newNet_1022;
wire newNet_20;
wire newNet_682;
wire n_18;
wire newNet_212;
wire n_173;
wire n_876;
wire cordic_SH2_srl_35_26_n_143;
wire n_239;
wire newNet_1180;
wire newNet_986;
wire newNet_501;
wire cordic_SH1_srl_35_26_n_72;
wire cordic_AddX_Btemp1_8_;
wire cordic_SH1_srl_35_26_n_145;
wire n_824;
wire newNet_717;
wire newNet_744;
wire cordic_SH1_srl_35_26_n_16;
wire n_309;
wire cordic_AddY_Compl_n_23;
wire n_337;
wire CoreOutputReg_29_;
wire n_251;
wire newNet_931;
wire cordic_AddX_Btemp_2_;
wire cordic_AddX_MUX_1_n_29;
wire PO_AD_28;
wire Dual_Cycle;
wire cordic_SH2_srl_35_26_n_42;
wire cordic_n_115;
wire n_492;
wire Config_Reg_3_;
wire newNet_991;
wire cordic_SH2_srl_35_26_n_87;
wire n_14;
wire n_594;
wire newNet_622;
wire cordic_AddY_MUX_0_n_3;
wire n_314;
wire PI_AD_32;
wire cordic_SH2_srl_35_26_n_83;
wire newNet_45;
wire PI_AD_3;
wire cordic_AddY_Btemp1_14_;
wire newNet_633;
wire cordic_AddX_Compl_n_6;
wire newNet_456;
wire cordic_Add0_MUX_1_n_24;
wire n_585;
wire n_761;
wire cordic_AddY_MUX_0_n_25;
wire cordic_Y_12_;
wire cordic_AddY_Add_n_22;
wire cordic_AddY_Btemp1_8_;
wire n_591;
wire newNet_402;
wire PO_AD_41;
wire newNet_43;
wire cordic_Add0_Compl_n_37;
wire newNet_1187;
wire n_307;
wire cordic_Add0_Atemp_15_;
wire n_327;
wire newNet_756;
wire newNet_58;
wire cordic_BS2_7_;
wire newNet_148;
wire cordic_SH2_srl_35_26_n_48;
wire newNet_1147;
wire CoreOutput_11_;
wire n_8;
wire newNet_1035;
wire cordic_Add0_Add_n_10;
wire n_600;
wire PIO_PAR_Value_Hold;
wire newNet_440;
wire newNet_1008;
wire newNet_1150;
wire newNet_920;
wire cordic_AddY_MUX_1_n_16;
wire cordic_SH1_srl_35_26_n_119;
wire n_746;
wire cordic_pla_n_28;
wire n_380;
wire newNet_1163;
wire n_442;
wire PO_PERR_L;
wire newNet_1205;
wire cordic_SH2_srl_35_26_n_10;
wire n_900;
wire newNet_1088;
wire newNet_231;
wire cordic_SumAngle_6_;
wire CoreOutputReg_8_;
wire newNet_347;
wire cordic_Add0_Add_n_66;
wire newNet_916;
wire n_137;
wire newNet_608;
wire n_129;
wire cordic_AddY_Add_n_29;
wire cordic_AddX_Add_n_31;
wire n_241;
wire PO_AD_37;
wire cordic_AddY_Add_n_56;
wire cordic_Add0_n_9;
wire cordic_SH2_srl_35_26_n_107;
wire newNet_912;
wire cordic_AddY_MUX_0_n_24;
wire CoreInput_11_;
wire CoreInput_1_;
wire cordic_SH1_srl_35_26_n_101;
wire cordic_SH2_srl_35_26_n_88;
wire n_297;
wire newNet_79;
wire n_520;
wire PI_AD_9;
wire cordic_AddX_Stemp_6_;
wire n_184;
wire cordic_X_10_;
wire PO_AD_48;
wire newNet_25;
wire cordic_n_54;
wire CoreOutput_25_;
wire n_331;
wire cordic_AddY_MUX_1_n_18;
wire n_189;
wire newNet_413;
wire cordic_AddX_MUX_0_n_16;
wire newNet_578;
wire cordic_SH1_srl_35_26_n_80;
wire cordic_n_32;
wire n_647;
wire cordic_Add0_MUX_1_n_3;
wire n_484;
wire newNet_940;
wire newNet_818;
wire n_353;
wire n_854;
wire newNet_292;
wire newNet_874;
wire cordic_AddY_MUX_0_n_29;
wire cordic_AddX_Btemp_10_;
wire n_157;
wire n_877;
wire newNet_494;
wire n_125;
wire n_323;
wire cordic_Add0_Stemp_1_;
wire cordic_AddX_Add_n_44;
wire newNet_336;
wire newNet_160;
wire Check_Add_Parity;
wire cordic_AddX_Add_n_53;
wire cordic_Add0_Atemp_9_;
wire n_724;
wire CoreOutput_18_;
wire cordic_AddX_Compl_n_37;
wire n_395;
wire n_883;
wire newNet_1034;
wire cordic_AddY_Add_n_24;
wire cordic_AddX_Add_n_74;
wire cordic_n_105;
wire n_763;
wire newNet_1014;
wire newNet_604;
wire cordic_AddX_MUX_1_n_2;
wire cordic_Add0_MUX_0_n_32;
wire cordic_SH1_srl_35_26_n_30;
wire cordic_AddX_Atemp_12_;
wire Access_Address_1_30_;
wire cordic_pla_n_9;
wire n_478;
wire newNet_297;
wire PI_AD_52;
wire n_227;
wire cordic_pla_n_13;
wire newNet_845;
wire cordic_AddY_Compl_n_14;
wire cordic_AddY_Btemp_5_;
wire n_507;
wire newNet_214;
wire cordic_AddX_Compl_n_0;
wire cordic_SH1_srl_35_26_n_124;
wire newNet_279;
wire cordic_AddY_MUX_1_n_5;
wire newNet_201;
wire n_223;
wire n_151;
wire newNet_286;
wire newNet_139;
wire PAR_Int;
wire newNet_140;
wire newNet_789;
wire PO_AD_36;
wire newNet_1186;
wire Access_Type_1_0_;
wire n_527;
wire newNet_881;
wire cordic_Add0_MUX_0_n_28;
wire PI_AD_41;
wire cordic_Add0_Add_n_1;
wire newNet_868;
wire cordic_Add0_Compl_n_4;
wire cordic_SH2_srl_35_26_n_77;
wire cordic_Add0_Compl_n_19;
wire cordic_AddY_Add_n_40;
wire newNet_722;
wire newNet_309;
wire newNet_791;
wire cordic_Y_9_;
wire cordic_n_113;
wire cordic_n_123;
wire PI_AD_57;
wire newNet_226;
wire cordic_SH2_srl_35_26_n_0;
wire cordic_Add0_MUX_0_n_20;
wire cordic_SH2_srl_35_26_n_128;
wire cordic_AddX_Compl_n_19;
wire newNet_984;
wire n_300;
wire cordic_AddX_Stemp_4_;
wire cordic_AddX_MUX_1_n_16;
wire n_97;
wire newNet_343;
wire cordic_AddY_Compl_n_33;
wire cordic_SH1_srl_35_26_n_139;
wire newNet_771;
wire n_561;
wire cordic_pla_n_18;
wire cordic_Add0_MUX_1_n_26;
wire newNet_572;
wire newNet_534;
wire Config_Reg_22_;
wire cordic_SH1_srl_35_26_n_79;
wire cordic_AddX_Add_n_27;
wire n_418;
wire newNet_234;
wire cordic_Add0_Compl_n_21;
wire n_809;
wire n_115;
wire n_70;
wire newNet_582;
wire newNet_188;
wire cordic_n_118;
wire n_190;
wire n_665;
wire CoreInput_5_;
wire newNet_732;
wire n_170;
wire CoreOutputReg_15_;
wire n_246;
wire newNet_777;
wire n_835;
wire newNet_357;
wire newNet_726;
wire cordic_AddY_Y_3;
wire cordic_SH1_srl_35_26_n_84;
wire cordic_Angle_8_;
wire cordic_SH2_srl_35_26_n_100;
wire cordic_AddY_Btemp_9_;
wire n_675;
wire n_693;
wire newNet_423;
wire cordic_Add0_MUX_1_n_15;
wire cordic_SumAngle_4_;
wire cordic_AddX_Add_n_7;
wire n_503;
wire cordic_SH1_srl_35_26_n_97;
wire newNet_958;
wire newNet_798;
wire n_867;
wire n_166;
wire n_195;
wire n_500;
wire newNet_1159;
wire cordic_AddX_MUX_0_n_32;
wire cordic_AddX_Atemp_5_;
wire cordic_AddX_Compl_n_35;
wire newNet_320;
wire newNet_522;
wire cordic_SH1_srl_35_26_n_0;
wire n_77;
wire n_739;
wire newNet_599;
wire cordic_SH2_srl_35_26_n_15;
wire newNet_368;
wire cordic_Add0_Add_n_59;
wire n_287;
wire cordic_SH1_srl_35_26_n_132;
wire newNet_321;
wire newNet_112;
wire newNet_169;
wire cordic_AddY_Stemp_10_;
wire cordic_AddY_Btemp1_9_;
wire cordic_Add0_Btemp_12_;
wire newNet_1160;
wire n_683;
wire cordic_Add0_MUX_1_n_18;
wire newNet_856;
wire cordic_Add0_Add_n_27;
wire newNet_781;
wire cordic_SH2_srl_35_26_n_119;
wire n_406;
wire newNet_1048;
wire newNet_539;
wire cordic_AddX_Atemp_8_;
wire n_827;
wire newNet_893;
wire n_565;
wire newNet_364;
wire cordic_AddX_Add_n_14;
wire cordic_AddY_Compl_n_39;
wire cordic_AddX_Stemp_15_;
wire n_312;
wire n_325;
wire cordic_AddX_MUX_0_n_28;
wire newNet_619;
wire newNet_742;
wire n_69;
wire newNet_1071;
wire newNet_352;
wire Config_Reg_16_;
wire newNet_450;
wire newNet_1074;
wire newNet_236;
wire newNet_122;
wire n_146;
wire cordic_X_9_;
wire newNet_267;
wire n_364;
wire cordic_AddY_Add_n_8;
wire n_825;
wire cordic_n_28;
wire n_461;
wire newNet_274;
wire newNet_241;
wire newNet_901;
wire cordic_AddY_MUX_0_n_0;
wire newNet_1067;
wire newNet_542;
wire cordic_Add0_MUX_1_n_29;
wire cordic_n_57;
wire newNet_545;
wire cordic_SH2_srl_35_26_n_45;
wire newNet_245;
wire newNet_65;
wire newNet_330;
wire newNet_48;
wire newNet_42;
wire n_58;
wire newNet_903;
wire PO_AD_14;
wire newNet_819;
wire cordic_Y_5_;
wire newNet_36;
wire cordic_tanangle_4_;
wire newNet_143;
wire cordic_AddY_Atemp_6_;
wire cordic_SH1_srl_35_26_n_117;
wire newNet_639;
wire newNet_107;
wire n_631;
wire cordic_AddX_Stemp_13_;
wire newNet_434;
wire PI_AD_6;
wire n_764;
wire newNet_915;
wire n_453;
wire n_543;
wire newNet_52;
wire cordic_tanangle_8_;
wire newNet_89;
wire PI_AD_27;
wire CoreInput_16_;
wire cordic_AddY_Add_n_49;
wire newNet_393;
wire cordic_AddY_Btemp_13_;
wire n_235;
wire newNet_835;
wire cordic_AddX_Compl_n_16;
wire CoreOutput_28_;
wire cordic_Add0_Add_n_69;
wire cordic_SH2_srl_35_26_n_74;
wire n_219;
wire cordic_AddY_Stemp_2_;
wire State_2_;
wire n_51;
wire newNet_1121;
wire n_607;
wire newNet_466;
wire newNet_258;
wire n_751;
wire cordic_Angle_5_;
wire cordic_SH1_srl_35_26_n_25;
wire newNet_833;
wire cordic_SH1_srl_35_26_n_68;
wire n_643;
wire newNet_408;
wire cordic_Add0_Add_n_60;
wire cordic_Add0_Btemp_14_;
wire cordic_Angle_4_;
wire cordic_SH1_srl_35_26_n_61;
wire n_85;
wire newNet_1191;
wire newNet_192;
wire newNet_1114;
wire newNet_656;
wire PI_AD_10;
wire n_279;
wire newNet_822;
wire newNet_563;
wire newNet_829;
wire newNet_1148;
wire newNet_643;
wire cordic_SH1_srl_35_26_n_143;
wire cordic_n_12;
wire TAR_TRI_T;
wire n_636;
wire newNet_603;
wire newNet_303;
wire newNet_1105;
wire cordic_Add0_Stemp_6_;
wire PO_AD_31;
wire newNet_93;
wire n_712;
wire cordic_Add0_n_14;
wire cordic_n_72;
wire newNet_636;
wire cordic_SH1_srl_35_26_n_7;
wire newNet_296;
wire cordic_SH1_srl_35_26_n_50;
wire newNet_82;
wire cordic_n_74;
wire n_132;
wire newNet_118;
wire cordic_AddY_MUX_0_n_32;
wire n_207;
wire n_632;
wire newNet_1041;
wire n_130;
wire newNet_308;
wire cordic_BS1_8_;
wire newNet_176;
wire Config_Reg_14_;
wire cordic_Add0_Add_n_56;
wire n_413;
wire newNet_1184;
wire n_690;
wire cordic_AddY_Compl_n_3;
wire cordic_SH1_srl_35_26_n_49;
wire newNet_704;
wire newNet_812;
wire cordic_n_97;
wire newNet_508;
wire newNet_668;
wire cordic_Add0_Compl_n_33;
wire n_32;
wire n_536;
wire PI_AD_31;
wire newNet_949;
wire cordic_SH1_srl_35_26_n_35;
wire CoreOutputReg_12_;
wire n_263;
wire cordic_AddX_Btemp1_12_;
wire newNet_925;
wire cordic_SH1_srl_35_26_n_44;
wire cordic_AddX_MUX_1_n_22;
wire newNet_531;
wire cordic_Add0_Add_n_42;
wire n_795;
wire newNet_1201;
wire cordic_AddX_Add_n_2;
wire n_818;
wire Access_Address_1_21_;
wire First_Entry;
wire newNet_100;
wire cordic_SumAngle_15_;
wire n_758;
wire n_176;
wire newNet_1018;
wire n_436;
wire cordic_AddY_Add_n_53;
wire cordic_AddX_Compl_n_1;
wire n_1;
wire newNet_1003;
wire newNet_778;
wire newNet_555;
wire cordic_n_86;
wire n_105;
wire Config_Reg_10_;
wire cordic_AddX_Stemp_10_;
wire newNet_54;
wire cordic_pla_n_6;
wire PI_AD_42;
wire n_801;
wire newNet_478;
wire newNet_1167;
wire newNet_389;
wire newNet_1197;
wire PO_AD_5;
wire n_497;
wire newNet_683;
wire cordic_AddX_MUX_0_n_14;
wire cordic_X_0_;
wire n_530;
wire newNet_1129;
wire cordic_pla_n_5;
wire newNet_1179;
wire cordic_Add0_Add_n_2;
wire n_21;
wire newNet_473;
wire PO_AD_6;
wire CoreOutputReg_2_;
wire newNet_1176;
wire cordic_AddX_Stemp_8_;
wire n_27;
wire newNet_718;
wire Check_Attr_Parity;
wire newNet_417;
wire newNet_208;
wire n_333;
wire cordic_AddX_n_1;
wire n_657;
wire newNet_377;
wire n_548;
wire newNet_612;
wire cordic_AddY_Add_n_18;
wire cordic_SH1_srl_35_26_n_56;
wire n_849;
wire newNet_337;
wire newNet_22;
wire PO_AD_50;
wire newNet_1204;
wire n_820;
wire cordic_n_144;
wire cordic_SH2_srl_35_26_n_96;
wire cordic_Add0_Add_n_8;
wire cordic_Add0_Add_n_47;
wire n_94;
wire cordic_SH2_srl_35_26_n_64;
wire PI_AD_63;
wire cordic_AddY_Add_n_35;
wire newNet_680;
wire newNet_311;
wire n_216;
wire newNet_998;
wire newNet_851;
wire cordic_Add0_n_4;
wire cordic_pla_n_21;
wire newNet_713;
wire cordic_AddY_Compl_n_25;
wire n_572;
wire cordic_AddY_Add_n_0;
wire n_700;
wire cordic_AddY_MUX_1_n_11;
wire n_446;
wire n_598;
wire cordic_Add0_Add_n_13;
wire PAR64_Int_d;
wire n_430;
wire n_551;
wire newNet_976;
wire newNet_802;
wire newNet_455;
wire newNet_690;
wire cordic_AddY_MUX_1_n_14;
wire cordic_Add0_Add_n_19;
wire cordic_AddY_MUX_1_n_32;
wire newNet_151;
wire Config_Reg_19_;
wire cordic_SH1_srl_35_26_n_110;
wire CoreInput_9_;
wire n_3;
wire cordic_AddY_Compl_n_19;
wire n_533;
wire n_40;
wire cordic_n_120;
wire cordic_AddX_Btemp_14_;
wire CoreOutput_9_;
wire cordic_AddY_MUX_0_n_9;
wire newNet_170;
wire n_857;
wire n_259;
wire n_17;
wire cordic_n_4;
wire n_887;
wire cordic_n_109;
wire cordic_SH1_srl_35_26_n_19;
wire newNet_671;
wire cordic_SH1_srl_35_26_n_15;
wire cordic_SH1_srl_35_26_n_133;
wire newNet_885;
wire newNet_80;
wire newNet_223;
wire newNet_16;
wire cordic_AddX_Add_n_23;
wire n_43;
wire n_782;
wire cordic_SH1_srl_35_26_n_3;
wire newNet_957;
wire cordic_SH1_srl_35_26_n_39;
wire PI_AD_46;
wire n_650;
wire cordic_SH2_srl_35_26_n_67;
wire newNet_1081;
wire newNet_427;
wire newNet_264;
wire Core_Cnt_3_;
wire n_554;
wire n_627;
wire newNet_1095;
wire n_33;
wire cordic_pla_n_16;
wire cordic_Add0_Add_n_24;
wire cordic_SH2_srl_35_26_n_6;
wire n_270;
wire PI_PAR;
wire n_336;
wire cordic_AddX_Stemp_9_;
wire TAR_TRI_S;
wire cordic_Y_0_;
wire n_0;
wire newNet_908;
wire cordic_n_3;
wire n_873;
wire newNet_968;
wire newNet_629;
wire Config_Reg_13_;
wire n_163;
wire n_400;
wire cordic_SumAngle_10_;
wire newNet_230;
wire cordic_SH2_srl_35_26_n_139;
wire n_573;
wire n_7;
wire n_757;
wire n_831;
wire newNet_57;
wire newNet_76;
wire newNet_708;
wire n_187;
wire newNet_1007;
wire n_468;
wire n_358;
wire cordic_n_87;
wire n_145;
wire cordic_Add0_MUX_1_n_11;
wire newNet_62;
wire cordic_AddX_Atemp_6_;
wire OutputAvail;
wire newNet_418;
wire n_82;
wire cordic_AddX_Add_n_11;
wire n_368;
wire n_352;
wire cordic_AddX_MUX_0_n_30;
wire Config_Reg_28_;
wire newNet_935;
wire n_771;
wire newNet_253;
wire n_792;
wire PO_AD_17;
wire cordic_SH2_srl_35_26_n_16;
wire n_821;
wire cordic_AddX_Add_n_59;
wire PO_AD_45;
wire newNet_1000;
wire n_475;
wire newNet_977;
wire cordic_AddY_Compl_n_2;
wire cordic_Add0_Btemp_0_;
wire n_480;
wire n_423;
wire newNet_942;
wire newNet_327;
wire RESET;
wire newNet_688;
wire newNet_999;
wire newNet_252;
wire n_136;
wire PO_AD_61;
wire n_387;
wire newNet_1151;
wire newNet_751;
wire cordic_tanangle_6_;
wire n_394;
wire cordic_Add0_MUX_0_n_0;
wire CoreOutputReg_11_;
wire newNet_447;
wire cordic_SH2_srl_35_26_n_36;
wire newNet_517;
wire n_890;
wire newNet_852;
wire newNet_196;
wire cordic_n_82;
wire newNet_1070;
wire newNet_677;
wire PO_PAR;
wire cordic_AddY_Add_n_13;
wire newNet_1156;
wire cordic_AddY_MUX_1_n_8;
wire cordic_Add0_Add_n_21;
wire cordic_AddY_MUX_1_n_1;
wire n_755;
wire cordic_AddY_MUX_1_n_31;
wire newNet_282;
wire n_339;
wire newNet_609;
wire n_844;
wire newNet_144;
wire n_443;
wire newNet_185;
wire cordic_AddY_Stemp_3_;
wire n_63;
wire cordic_SH1_srl_35_26_n_26;
wire n_723;
wire newNet_270;
wire cordic_Add0_MUX_1_n_2;
wire cordic_AddX_Compl_n_4;
wire PI_AD_19;
wire cordic_AddX_Compl_n_21;
wire n_283;
wire n_697;
wire newNet_154;
wire cordic_SH2_srl_35_26_n_4;
wire Config_Reg_0_;
wire cordic_AddY_Add_n_9;
wire cordic_SH2_srl_35_26_n_29;
wire n_734;
wire cordic_AddX_n_5;
wire cordic_BS2_5_;
wire newNet_1080;
wire cordic_n_103;
wire cordic_Add0_Btemp_15_;
wire cordic_n_13;
wire newNet_1196;
wire newNet_824;
wire n_199;
wire cordic_Add0_Compl_n_0;
wire cordic_AddY_MUX_0_n_14;
wire newNet_420;
wire n_291;
wire n_194;
wire n_275;
wire newNet_953;
wire newNet_586;
wire cordic_Add0_MUX_1_n_9;
wire cordic_n_36;
wire n_842;
wire newNet_699;
wire n_504;
wire cordic_tanangle_0_;
wire n_870;
wire n_301;
wire newNet_785;
wire newNet_767;
wire cordic_Add0_MUX_1_n_14;
wire n_278;
wire newNet_126;
wire newNet_898;
wire PI_CBE_L_3;
wire newNet_275;
wire cordic_SH2_srl_35_26_n_84;
wire n_686;
wire n_593;
wire newNet_1143;
wire n_375;
wire newNet_600;
wire n_689;
wire cordic_Add0_Compl_n_13;
wire cordic_SH2_srl_35_26_n_94;
wire cordic_AddY_MUX_0_n_28;
wire n_108;
wire newNet_165;
wire n_111;
wire n_73;
wire n_142;
wire n_121;
wire n_569;
wire newNet_458;
wire n_399;
wire Access_Address_1_18_;
wire n_806;
wire cordic_AddX_MUX_1_n_21;
wire cordic_n_21;
wire n_679;
wire n_280;
wire newNet_557;
wire newNet_31;
wire n_118;
wire cordic_AddY_Compl_n_10;
wire cordic_AddY_Stemp_15_;
wire n_786;
wire n_897;
wire n_16;
wire cordic_Y_1_;
wire CoreInput_14_;
wire cordic_AddX_Add_n_50;
wire cordic_Add0_MUX_1_n_7;
wire newNet_863;
wire CoreOutput_8_;
wire cordic_AddY_Btemp1_0_;
wire PO_AD_20;
wire cordic_AddX_MUX_0_n_4;
wire n_489;
wire cordic_n_64;
wire n_523;
wire cordic_SH2_srl_35_26_n_110;
wire newNet_620;
wire cordic_SH1_srl_35_26_n_89;
wire Config_Reg_31_;
wire newNet_792;
wire newNet_616;
wire cordic_SH2_srl_35_26_n_60;
wire cordic_AddX_Btemp1_4_;
wire newNet_990;
wire newNet_6;
wire cordic_Add0_n_3;
wire newNet_358;
wire cordic_Add0_n_8;
wire cordic_n_114;
wire n_705;
wire cordic_AddX_Stemp_12_;
wire cordic_n_24;
wire newNet_500;
wire cordic_BS1_15_;
wire cordic_SH2_srl_35_26_n_11;
wire n_36;
wire newNet_640;
wire newNet_595;
wire cordic_Add0_MUX_1_n_25;
wire newNet_747;
wire cordic_AddY_MUX_1_n_20;
wire newNet_475;
wire newNet_987;
wire newNet_69;
wire n_260;
wire cordic_Add0_Atemp_11_;
wire n_66;
wire n_456;
wire newNet_1;
wire newNet_213;
wire newNet_1164;
wire cordic_AddY_Stemp_1_;
wire cordic_AddX_Compl_n_25;
wire cordic_AddY_MUX_0_n_10;
wire n_760;
wire newNet_266;
wire cordic_AddX_Btemp1_15_;
wire newNet_736;
wire cordic_AddY_Add_n_67;
wire newNet_1183;
wire newNet_1050;
wire Access_Address_1_26_;
wire Access_Address_1_16_;
wire newNet_994;
wire newNet_980;
wire newNet_552;
wire cordic_SH2_srl_35_26_n_71;
wire cordic_AddY_MUX_1_n_15;
wire newNet_541;
wire cordic_n_92;
wire cordic_AddX_MUX_1_n_12;
wire cordic_SH1_srl_35_26_n_93;
wire n_308;
wire newNet_147;
wire cordic_SH2_srl_35_26_n_43;
wire n_428;
wire newNet_300;
wire n_265;
wire cordic_Add0_Compl_n_6;
wire n_517;
wire cordic_AddY_MUX_1_n_25;
wire CoreOutputReg_22_;
wire newNet_566;
wire n_254;
wire newNet_1099;
wire n_13;
wire n_646;
wire newNet_382;
wire cordic_AddX_Compl_n_5;
wire cordic_AddY_Stemp_8_;
wire cordic_SH1_srl_35_26_n_75;
wire n_791;
wire n_238;
wire newNet_1062;
wire n_747;
wire newNet_1136;
wire n_635;
wire cordic_Add0_Add_n_65;
wire n_47;
wire cordic_Add0_Add_n_36;
wire n_242;
wire newNet_794;
wire newNet_700;
wire n_240;
wire cordic_AddX_Add_n_30;
wire CoreOutputReg_0_;
wire n_403;
wire cordic_AddX_Btemp1_9_;
wire Access_Type_1_3_;
wire cordic_AddY_Atemp_3_;
wire cordic_AddY_Stemp_11_;
wire PI_AD_14;
wire newNet_1200;
wire newNet_111;
wire cordic_X_13_;
wire newNet_114;
wire cordic_SH2_srl_35_26_n_53;
wire newNet_104;
wire n_669;
wire PI_AD_2;
wire newNet_1125;
wire newNet_647;
wire cordic_AddY_Btemp1_6_;
wire n_672;
wire newNet_179;
wire n_464;
wire cordic_Add0_MUX_1_n_32;
wire DevSel_Wait_Cnt_1_;
wire newNet_809;
wire n_660;
wire newNet_642;
wire cordic_AddY_Atemp_7_;
wire newNet_490;
wire PO_AD_57;
wire n_215;
wire n_319;
wire newNet_135;
wire n_860;
wire n_564;
wire cordic_AddY_Add_n_4;
wire cordic_AddX_MUX_0_n_10;
wire n_617;
wire n_441;
wire cordic_AddX_MUX_1_n_9;
wire cordic_AddY_Compl_n_29;
wire newNet_86;
wire n_740;
wire newNet_209;
wire cordic_AddY_MUX_0_n_19;
wire n_738;
wire cordic_SH1_srl_35_26_n_41;
wire cordic_AddY_Add_n_74;
wire newNet_131;
wire CoreOutputReg_5_;
wire cordic_AddX_Compl_n_12;
wire CBE_par_2_;
wire n_24;
wire n_295;
wire cordic_SH1_srl_35_26_n_21;
wire cordic_SH1_srl_35_26_n_114;
wire n_212;
wire newNet_37;
wire newNet_839;
wire cordic_SH2_srl_35_26_n_32;
wire n_582;
wire cordic_SH2_srl_35_26_n_116;
wire n_654;
wire n_416;
wire n_156;
wire newNet_649;
wire cordic_AddX_Btemp_12_;
wire n_614;
wire newNet_438;
wire cordic_Add0_Compl_n_41;
wire n_579;
wire PO_AD_2;
wire newNet_1131;
wire n_588;
wire n_101;
wire Trdy_Wait_Cnt_1_;
wire cordic_SH1_srl_35_26_n_128;
wire n_370;
wire newNet_512;
wire cordic_tanangle_7_;
wire newNet_945;
wire n_343;
wire cordic_SH2_srl_35_26_n_78;
wire cordic_pla_n_2;
wire n_54;
wire newNet_972;
wire cordic_Angle_14_;
wire newNet_403;
wire newNet_395;
wire PI_AD_35;
wire cordic_Add0_MUX_1_n_21;
wire cordic_AddY_Add_n_31;
wire newNet_815;
wire newNet_372;
wire cordic_Add0_MUX_0_n_18;
wire cordic_n_46;
wire newNet_1059;
wire cordic_n_7;
wire PI_AD_45;
wire cordic_n_78;
wire newNet_535;
wire n_172;
wire cordic_AddY_MUX_0_n_4;
wire n_703;
wire newNet_1171;
wire cordic_Y_6_;
wire newNet_1100;
wire newNet_1027;
wire newNet_470;
wire n_313;
wire cordic_tanangle_13_;
wire cordic_tanangle_11_;
wire newNet_723;
wire n_390;
wire newNet_663;
wire cordic_SH1_srl_35_26_n_48;
wire cordic_n_52;
wire n_493;
wire cordic_tanangle_2_;
wire newNet_568;
wire cordic_Y_7_;
wire n_775;
wire cordic_Add0_Btemp_10_;
wire PO_AD_10;
wire PO_AD_1;
wire n_346;
wire n_628;
wire newNet_946;
wire cordic_Add0_Compl_n_1;
wire cordic_SH2_srl_35_26_n_133;
wire cordic_AddX_Add_n_3;
wire cordic_n_40;
wire newNet_929;
wire PI_AD_53;
wire cordic_n_110;
wire newNet_1079;
wire newNet_1021;
wire newNet_298;
wire PO_AD_27;
wire newNet_218;
wire cordic_SH1_srl_35_26_n_78;
wire n_479;
wire n_664;
wire newNet_1039;
wire cordic_AddY_Stemp_5_;
wire PI_AD_37;
wire cordic_AddY_Atemp_1_;
wire newNet_745;
wire newNet_738;
wire cordic_AddY_Add_n_21;
wire n_160;
wire newNet_930;
wire newNet_483;
wire Idsel;
wire cordic_Add0_Compl_n_27;
wire n_232;
wire newNet_536;
wire newNet_193;
wire n_694;
wire newNet_684;
wire newNet_414;
wire cordic_AddX_MUX_0_n_15;
wire cordic_Add0_Add_n_3;
wire n_592;
wire cordic_SH1_srl_35_26_n_86;
wire n_611;
wire cordic_SH1_srl_35_26_n_47;
wire newNet_314;
wire cordic_Add0_Compl_n_39;
wire cordic_Add0_Add_n_35;
wire newNet_973;
wire cordic_BS2_15_;
wire n_616;
wire newNet_1137;
wire newNet_651;
wire CoreOutputReg_30_;
wire newNet_38;
wire newNet_804;
wire newNet_318;
wire newNet_653;
wire n_584;
wire PI_AD_1;
wire newNet_1002;
wire cordic_AddX_Compl_n_10;
wire n_815;
wire newNet_985;
wire newNet_101;
wire n_640;
wire cordic_SH1_srl_35_26_n_95;
wire cordic_AddY_Add_n_50;
wire PO_AD_4;
wire newNet_876;
wire newNet_846;
wire newNet_189;
wire n_305;
wire cordic_n_94;
wire n_179;
wire newNet_113;
wire n_550;
wire cordic_SH2_srl_35_26_n_113;
wire newNet_53;
wire cordic_Add0_Btemp_4_;
wire n_247;
wire cordic_SH2_srl_35_26_n_95;
wire n_549;
wire n_599;
wire cordic_AddY_Stemp_6_;
wire n_318;
wire newNet_1168;
wire newNet_611;
wire cordic_AddX_Compl_n_27;
wire newNet_799;
wire n_535;
wire cordic_SH1_srl_35_26_n_113;
wire newNet_26;
wire n_772;
wire n_808;
wire n_426;
wire newNet_374;
wire cordic_Add0_Add_n_32;
wire newNet_1085;
wire cordic_AddY_Add_n_62;
wire n_404;
wire n_789;
wire cordic_AddX_Add_n_38;
wire TAR_TRI_E;
wire cordic_n_90;
wire PI_AD_20;
wire newNet_1161;
wire newNet_1177;
wire newNet_157;
wire n_828;
wire Access_Type_1_2_;
wire n_391;
wire cordic_SH1_srl_35_26_n_12;
wire n_557;
wire cordic_AngleCin;
wire cordic_Add0_Add_n_9;
wire newNet_618;
wire cordic_Add0_Compl_n_23;
wire cordic_AddX_Stemp_2_;
wire n_435;
wire newNet_1115;
wire newNet_108;
wire cordic_Add0_Stemp_14_;
wire newNet_150;
wire cordic_AddY_Add_n_41;
wire n_262;
wire newNet_1109;
wire cordic_AddY_MUX_0_n_12;
wire newNet_220;
wire cordic_SH2_srl_35_26_n_9;
wire n_6;
wire newNet_331;
wire newNet_269;
wire n_159;
wire n_511;
wire CoreOutput_22_;
wire Trdy_Wait_Cnt_0_;
wire n_154;
wire n_37;
wire cordic_pla_n_1;
wire PO_AD_15;
wire newNet_119;
wire n_826;
wire newNet_1075;
wire newNet_801;
wire cordic_Add0_MUX_1_n_6;
wire cordic_Add0_Add_n_68;
wire newNet_3;
wire newNet_158;
wire cordic_AddY_MUX_0_n_23;
wire cordic_Angle_13_;
wire n_653;
wire cordic_Add0_MUX_1_n_30;
wire cordic_AddY_Btemp_0_;
wire n_141;
wire newNet_400;
wire newNet_914;
wire n_361;
wire cordic_SumAngle_11_;
wire cordic_SH2_srl_35_26_n_57;
wire n_748;
wire cordic_SH2_srl_35_26_n_89;
wire n_126;
wire n_183;
wire newNet_257;
wire newNet_116;
wire n_566;
wire newNet_51;
wire n_853;
wire n_528;
wire n_637;
wire cordic_AddX_Compl_n_8;
wire newNet_904;
wire n_447;
wire n_360;
wire cordic_AddX_MUX_1_n_3;
wire newNet_23;
wire CoreOutput_2_;
wire n_450;
wire n_234;
wire cordic_n_63;
wire newNet_47;
wire cordic_AddY_MUX_0_n_17;
wire CoreOutputReg_24_;
wire newNet_625;
wire newNet_1044;
wire newNet_624;
wire newNet_832;
wire cordic_Add0_n_7;
wire newNet_41;
wire cordic_AddY_Stemp_12_;
wire n_715;
wire n_644;
wire cordic_AddY_Compl_n_21;
wire newNet_474;
wire n_52;
wire cordic_AddY_MUX_0_n_1;
wire n_424;
wire newNet_66;
wire newNet_207;
wire newNet_121;
wire PI_CBE_L_5;
wire cordic_Add0_Add_n_39;
wire cordic_SH1_srl_35_26_n_144;
wire cordic_n_67;
wire newNet_964;
wire newNet_635;
wire CoreOutput_20_;
wire newNet_0;
wire cordic_tanangle_12_;
wire cordic_SH1_srl_35_26_n_90;
wire n_218;
wire cordic_Add0_Stemp_3_;
wire newNet_1053;
wire cordic_AddY_Compl_n_4;
wire newNet_392;
wire cordic_AddY_Atemp_5_;
wire cordic_SH1_srl_35_26_n_8;
wire n_716;
wire newNet_1049;
wire newNet_714;
wire PO_SERR_L;
wire cordic_SH2_srl_35_26_n_145;
wire newNet_503;
wire newNet_137;
wire n_630;
wire cordic_n_77;
wire n_731;
wire newNet_776;
wire newNet_544;
wire newNet_939;
wire newNet_204;
wire n_253;
wire newNet_461;
wire newNet_431;
wire cordic_AddX_MUX_1_n_8;
wire cordic_Y_2_;
wire n_459;
wire n_794;
wire PO_AD_30;
wire newNet_446;
wire newNet_762;
wire n_135;
wire newNet_94;
wire newNet_1189;
wire PI_AD_50;
wire newNet_467;
wire newNet_1077;
wire n_623;
wire cordic_AddY_Add_n_77;
wire cordic_Add0_Compl_n_7;
wire newNet_1005;
wire cordic_SH1_srl_35_26_n_36;
wire PO_AD_35;
wire newNet_1019;
wire cordic_SH2_srl_35_26_n_50;
wire n_680;
wire cordic_n_85;
wire cordic_SH2_srl_35_26_n_35;
wire cordic_AddX_Add_n_19;
wire n_812;
wire cordic_AddX_Add_n_47;
wire Config_Reg_24_;
wire n_161;
wire cordic_Add0_Add_n_41;
wire n_381;
wire n_315;
wire cordic_n_81;
wire cordic_Add0_Add_n_20;
wire cordic_SH1_srl_35_26_n_96;
wire n_720;
wire newNet_197;
wire cordic_AddX_Add_n_8;
wire newNet_959;
wire newNet_900;
wire newNet_1123;
wire newNet_864;
wire newNet_592;
wire cordic_BS2_13_;
wire PI_AD_18;
wire PO_AD_39;
wire cordic_AddX_Add_n_41;
wire cordic_Add0_Compl_n_10;
wire newNet_581;
wire n_896;
wire newNet_770;
wire n_878;
wire PI_AD_30;
wire cordic_SH2_srl_35_26_n_28;
wire cordic_AddY_Y_4;
wire cordic_BS1_5_;
wire newNet_439;
wire cordic_SH2_srl_35_26_n_61;
wire newNet_363;
wire newNet_453;
wire cordic_SH2_srl_35_26_n_70;
wire CoreOutput_4_;
wire cordic_AddY_Btemp1_3_;
wire newNet_1128;
wire PO_AD_42;
wire n_514;
wire newNet_1033;
wire cordic_X_12_;
wire cordic_AddX_Add_n_67;
wire cordic_AddY_Y_2;
wire cordic_AddY_Stemp_4_;
wire cordic_AddX_MUX_1_n_15;
wire n_167;
wire cordic_Add0_Btemp_8_;
wire PO_AD_62;
wire cordic_AddX_MUX_0_n_24;
wire n_886;
wire Access_Address_1_28_;
wire n_674;
wire n_560;
wire newNet_1203;
wire newNet_733;
wire cordic_SH2_srl_35_26_n_114;
wire n_369;
wire cordic_Add0_Compl_n_15;
wire newNet_698;
wire cordic_SH1_srl_35_26_n_85;
wire newNet_75;
wire cordic_AddX_Btemp_11_;
wire newNet_17;
wire PO_AD_23;
wire cordic_n_112;
wire n_691;
wire cordic_n_106;
wire newNet_344;
wire newNet_367;
wire newNet_897;
wire n_412;
wire cordic_n_84;
wire CoreOutput_19_;
wire newNet_495;
wire n_518;
wire CoreOutput_26_;
wire cordic_SH1_srl_35_26_n_71;
wire newNet_596;
wire cordic_AddY_Compl_n_7;
wire newNet_556;
wire n_138;
wire Access_Address_1_19_;
wire n_490;
wire n_769;
wire Config_Reg_7_;
wire Access_Address_1_22_;
wire n_759;
wire cordic_SH1_srl_35_26_n_1;
wire newNet_859;
wire cordic_n_17;
wire CBE_par_0_;
wire cordic_Add0_Add_n_28;
wire cordic_AddY_Add_n_38;
wire cordic_pla_n_17;
wire n_330;
wire PI_AD_49;
wire n_871;
wire cordic_AddY_Stemp_14_;
wire newNet_239;
wire newNet_142;
wire newNet_354;
wire cordic_AddY_n_3;
wire newNet_429;
wire newNet_506;
wire newNet_869;
wire n_354;
wire cordic_SH1_srl_35_26_n_129;
wire n_211;
wire newNet_667;
wire PI_AD_26;
wire cordic_SumAngle_9_;
wire cordic_Add0_Add_n_72;
wire cordic_SH1_srl_35_26_n_106;
wire CoreOutput_23_;
wire CoreOutput_7_;
wire newNet_969;
wire n_460;
wire newNet_527;
wire n_286;
wire CoreOutputReg_6_;
wire n_220;
wire PI_AD_40;
wire newNet_399;
wire cordic_SH2_srl_35_26_n_3;
wire cordic_Y_13_;
wire cordic_AddX_Compl_n_17;
wire PI_AD_62;
wire n_407;
wire n_521;
wire n_250;
wire newNet_755;
wire n_329;
wire newNet_614;
wire newNet_287;
wire n_209;
wire newNet_854;
wire newNet_128;
wire n_116;
wire n_42;
wire cordic_AddY_Btemp1_10_;
wire newNet_322;
wire n_322;
wire cordic_AddY_Add_n_3;
wire cordic_Add0_Add_n_25;
wire cordic_n_5;
wire n_342;
wire newNet_1026;
wire cordic_AddX_MUX_1_n_31;
wire cordic_SH2_srl_35_26_n_103;
wire PI_CBE_L_2;
wire TAR_TRI_A;
wire newNet_1119;
wire newNet_410;
wire Config_Reg_5_;
wire newNet_570;
wire newNet_180;
wire n_575;
wire cordic_AddX_Add_n_77;
wire newNet_254;
wire cordic_SH2_srl_35_26_n_12;
wire n_856;
wire newNet_295;
wire n_388;
wire cordic_Add0_MUX_0_n_12;
wire cordic_AddX_MUX_0_n_1;
wire cordic_AddX_Compl_n_9;
wire n_206;
wire cordic_SH1_srl_35_26_n_69;
wire n_396;
wire n_559;
wire cordic_SH2_srl_35_26_n_124;
wire cordic_SH1_srl_35_26_n_28;
wire n_709;
wire cordic_SH2_srl_35_26_n_129;
wire newNet_892;
wire n_540;
wire n_472;
wire newNet_227;
wire n_864;
wire cordic_n_55;
wire PI_AD_58;
wire cordic_SH2_srl_35_26_n_130;
wire Config_Reg_23_;
wire newNet_909;
wire n_744;
wire cordic_AddX_Compl_n_31;
wire n_725;
wire n_109;
wire cordic_AddX_MUX_0_n_17;
wire cordic_Add0_Add_n_53;
wire cordic_AddX_Btemp1_1_;
wire newNet_786;
wire newNet_468;
wire n_224;
wire newNet_871;
wire newNet_215;
wire n_762;
wire cordic_n_11;
wire CoreOutputReg_33_;
wire newNet_273;
wire newNet_646;
wire cordic_BS2_1_;
wire newNet_605;
wire cordic_SH2_srl_35_26_n_82;
wire cordic_BS2_14_;
wire cordic_SH1_srl_35_26_n_24;
wire n_282;
wire n_638;
wire n_340;
wire newNet_442;
wire newNet_305;
wire newNet_507;
wire PO_AD_59;
wire n_415;
wire cordic_AddX_MUX_1_n_30;
wire n_345;
wire n_338;
wire PO_AD_24;
wire newNet_694;
wire newNet_178;
wire PO_AD_9;
wire n_604;
wire newNet_585;
wire cordic_SH2_srl_35_26_n_99;
wire cordic_SH2_srl_35_26_n_54;
wire cordic_AddX_MUX_0_n_11;
wire n_102;
wire newNet_1098;
wire newNet_840;
wire newNet_630;
wire cordic_AddX_MUX_1_n_27;
wire n_444;
wire newNet_1104;
wire n_668;
wire cordic_AddY_Add_n_25;
wire CoreOutputReg_16_;
wire Config_Reg_9_;
wire cordic_pla_n_24;
wire n_570;
wire n_357;
wire n_408;
wire n_698;
wire n_613;
wire newNet_488;
wire n_733;
wire n_228;
wire newNet_601;
wire newNet_518;
wire cordic_n_41;
wire cordic_AddY_Atemp_9_;
wire newNet_850;
wire newNet_808;
wire n_268;
wire cordic_Add0_Add_n_62;
wire newNet_491;
wire cordic_SH1_srl_35_26_n_31;
wire cordic_AngleCout;
wire newNet_924;
wire n_819;
wire n_776;
wire newNet_657;
wire cordic_SH1_srl_35_26_n_62;
wire n_439;
wire n_237;
wire n_214;
wire cordic_pla_n_7;
wire PO_ACK64_L;
wire newNet_719;
wire newNet_454;
wire newNet_1172;
wire n_22;
wire cordic_AddY_Btemp1_5_;
wire cordic_SH2_srl_35_26_n_5;
wire newNet_200;
wire n_177;
wire cordic_n_22;
wire newNet_1142;
wire newNet_813;
wire cordic_SH1_srl_35_26_n_57;
wire n_663;
wire cordic_AddX_Compl_n_13;
wire cordic_Add0_MUX_1_n_22;
wire newNet_569;
wire n_316;
wire newNet_404;
wire cordic_X_5_;
wire n_850;
wire n_589;
wire n_741;
wire n_93;
wire cordic_Add0_Stemp_15_;
wire newNet_554;
wire cordic_AddY_MUX_0_n_13;
wire n_420;
wire cordic_AddX_n_2;
wire newNet_263;
wire n_785;
wire n_704;
wire n_602;
wire newNet_378;
wire newNet_746;
wire cordic_Y_11_;
wire newNet_1030;
wire newNet_13;
wire cordic_SH2_srl_35_26_n_93;
wire n_805;
wire PO_AD_0;
wire n_488;
wire cordic_SH1_srl_35_26_n_14;
wire PI_AD_38;
wire cordic_SH1_srl_35_26_n_125;
wire n_119;
wire cordic_n_58;
wire PI_AD_44;
wire newNet_638;
wire cordic_Add0_n_11;
wire cordic_AddX_Add_n_9;
wire newNet_11;
wire n_702;
wire cordic_AddX_MUX_1_n_23;
wire n_88;
wire Config_Reg_17_;
wire n_463;
wire newNet_1056;
wire cordic_AddY_Compl_n_0;
wire newNet_793;
wire newNet_219;
wire n_335;
wire newNet_1182;
wire cordic_Add0_n_2;
wire cordic_Add0_Compl_n_14;
wire newNet_1082;
wire cordic_Add0_MUX_1_n_0;
wire PI_AD_54;
wire Set_Data_Parity;
wire cordic_Add0_MUX_1_n_13;
wire newNet_265;
wire cordic_Add0_Btemp_9_;
wire cordic_AddX_Atemp_15_;
wire n_553;
wire newNet_838;
wire newNet_615;
wire newNet_1118;
wire PI_FRAME_L;
wire newNet_685;
wire cordic_AddY_Atemp_10_;
wire cordic_SH1_srl_35_26_n_33;
wire cordic_n_49;
wire newNet_373;
wire newNet_486;
wire newNet_498;
wire cordic_SH2_srl_35_26_n_81;
wire newNet_981;
wire newNet_954;
wire newNet_724;
wire newNet_349;
wire cordic_SH1_srl_35_26_n_120;
wire n_55;
wire cordic_n_107;
wire newNet_190;
wire Config_Reg_21_;
wire n_596;
wire cordic_SH2_srl_35_26_n_21;
wire cordic_Angle_12_;
wire n_874;
wire n_711;
wire cordic_Add0_Atemp_7_;
wire cordic_AddY_MUX_0_n_31;
wire newNet_997;
wire newNet_978;
wire newNet_409;
wire cordic_AddY_Add_n_20;
wire n_243;
wire newNet_1006;
wire newNet_210;
wire newNet_90;
wire PO_AD_33;
wire cordic_AddY_Compl_n_43;
wire CoreOutputReg_23_;
wire cordic_Add0_Compl_n_35;
wire n_401;
wire newNet_567;
wire newNet_1165;
wire newNet_641;
wire newNet_988;
wire newNet_115;
wire newNet_540;
wire newNet_146;
wire tau_clk;
wire cordic_AddX_Add_n_10;
wire newNet_233;
wire newNet_496;
wire n_634;
wire cordic_SH1_srl_35_26_n_74;
wire cordic_AddX_Compl_n_41;
wire newNet_1132;
wire newNet_302;
wire n_790;
wire newNet_1149;
wire newNet_27;
wire CoreOutputReg_3_;
wire cordic_AddY_Btemp1_7_;
wire newNet_933;
wire cordic_AddY_MUX_1_n_21;
wire cordic_AddY_Compl_n_27;
wire cordic_AddY_Atemp_12_;
wire n_139;
wire cordic_AddX_Add_n_35;
wire n_583;
wire CoreOutput_21_;
wire newNet_551;
wire newNet_415;
wire newNet_993;
wire newNet_105;
wire n_973;
wire n_580;
wire cordic_AddY_Btemp_14_;
wire cordic_SH2_srl_35_26_n_85;
wire PO_AD_11;
wire cordic_SH2_srl_35_26_n_115;
wire newNet_934;
wire newNet_795;
wire cordic_Y_15_;
wire cordic_AddX_Y_4;
wire n_767;
wire cordic_pla_n_26;
wire n_822;
wire cordic_Add0_Btemp_7_;
wire cordic_SH2_srl_35_26_n_46;
wire Trdy_Wait_Cnt_3_;
wire cordic_n_29;
wire cordic_AddX_Btemp_9_;
wire cordic_AddY_Add_n_27;
wire newNet_85;
wire cordic_AddY_Btemp_10_;
wire cordic_AddX_Compl_n_3;
wire n_544;
wire n_122;
wire newNet_750;
wire newNet_560;
wire cordic_Add0_Atemp_8_;
wire CoreInput_7_;
wire cordic_n_66;
wire newNet_524;
wire cordic_AddY_Add_n_46;
wire n_457;
wire newNet_1152;
wire newNet_129;
wire cordic_SH1_srl_35_26_n_107;
wire newNet_579;
wire cordic_SH2_srl_35_26_n_75;
wire n_546;
wire cordic_AddX_MUX_0_n_27;
wire cordic_AddY_MUX_1_n_30;
wire newNet_510;
wire n_23;
wire cordic_SH2_srl_35_26_n_118;
wire Par_Sgnl;
wire cordic_AddY_Add_n_14;
wire newNet_182;
wire newNet_4;
wire cordic_SH1_srl_35_26_n_65;
wire newNet_32;
wire cordic_SH2_srl_35_26_n_39;
wire newNet_1192;
wire newNet_1124;
wire cordic_X_14_;
wire cordic_AddX_Atemp_13_;
wire newNet_919;
wire newNet_1157;
wire cordic_AddY_Add_n_73;
wire PI_CBE_L_4;
wire cordic_AddY_Compl_n_37;
wire cordic_n_117;
wire n_203;
wire cordic_n_91;
wire CoreOutput_33_;
wire cordic_Add0_MUX_1_n_1;
wire n_90;
wire newNet_351;
wire CoreOutputReg_14_;
wire newNet_825;
wire cordic_AddY_MUX_0_n_18;
wire n_62;
wire n_155;
wire cordic_AddX_Add_n_71;
wire n_510;
wire cordic_SH1_srl_35_26_n_81;
wire n_311;
wire newNet_9;
wire newNet_283;
wire n_781;
wire cordic_Add0_MUX_1_n_17;
wire cordic_SH2_srl_35_26_n_31;
wire n_294;
wire n_671;
wire newNet_573;
wire cordic_SH2_srl_35_26_n_25;
wire n_687;
wire PO_TRDY_L;
wire newNet_394;
wire PI_AD_34;
wire cordic_AddX_MUX_0_n_5;
wire newNet_928;
wire n_30;
wire PO_AD_18;
wire cordic_n_61;
wire newNet_782;
wire cordic_AddY_Add_n_34;
wire newNet_523;
wire cordic_AddY_MUX_1_n_4;
wire cordic_Add0_Stemp_9_;
wire n_458;
wire n_524;
wire cordic_AddX_Compl_n_29;
wire n_799;
wire cordic_SumAngle_1_;
wire cordic_n_14;
wire cordic_n_98;
wire newNet_816;
wire PI_AD_23;
wire newNet_664;
wire newNet_136;
wire n_508;
wire n_196;
wire n_501;
wire n_532;
wire newNet_168;
wire cordic_AddY_Add_n_15;
wire newNet_125;
wire n_112;
wire cordic_X_1_;
wire newNet_741;
wire cordic_SH1_srl_35_26_n_4;
wire cordic_Add0_MUX_0_n_9;
wire cordic_AddX_MUX_1_n_0;
wire cordic_AddX_Stemp_1_;
wire cordic_BS1_4_;
wire newNet_1047;
wire n_379;
wire n_678;
wire newNet_855;
wire newNet_246;
wire cordic_AddY_MUX_1_n_10;
wire newNet_132;
wire cordic_AddX_Add_n_4;
wire n_882;
wire Check_Data_Parity;
wire n_276;
wire cordic_Add0_Add_n_45;
wire cordic_BS2_0_;
wire cordic_AddX_MUX_0_n_7;
wire n_816;
wire cordic_n_33;
wire n_752;
wire newNet_340;
wire newNet_528;
wire cordic_AddX_MUX_0_n_0;
wire cordic_AddX_Btemp1_7_;
wire cordic_Add0_Add_n_18;
wire newNet_737;
wire Config_Reg_12_;
wire cordic_pla_n_12;
wire newNet_950;
wire newNet_1009;
wire newNet_1010;
wire cordic_SumAngle_5_;
wire newNet_430;
wire n_60;
wire newNet_72;
wire n_164;
wire n_81;
wire newNet_965;
wire newNet_97;
wire cordic_BS2_6_;
wire newNet_650;
wire n_186;
wire n_248;
wire n_626;
wire newNet_1094;
wire newNet_173;
wire n_302;
wire cordic_AddX_Add_n_62;
wire cordic_SH1_srl_35_26_n_52;
wire n_289;
wire newNet_759;
wire Trdy_Wait_Cnt_2_;
wire cordic_SH1_srl_35_26_n_92;
wire Config_Reg_25_;
wire newNet_710;
wire newNet_224;
wire Config_Reg_26_;
wire newNet_383;
wire n_832;
wire cordic_AddY_Btemp_15_;
wire n_384;
wire n_144;
wire newNet_830;
wire n_67;
wire newNet_831;
wire cordic_AddX_MUX_1_n_11;
wire newNet_880;
wire cordic_Add0_MUX_1_n_10;
wire newNet_1113;
wire newNet_889;
wire cordic_Add0_Compl_n_31;
wire cordic_SH2_srl_35_26_n_68;
wire Config_Reg_11_;
wire newNet_1051;
wire n_365;
wire cordic_n_122;
wire newNet_1061;
wire PO_AD_54;
wire n_836;
wire n_150;
wire cordic_AddY_MUX_1_n_17;
wire n_695;
wire cordic_Add0_Y_3;
wire cordic_Add0_Add_n_29;
wire newNet_513;
wire newNet_84;
wire cordic_AddY_Btemp_2_;
wire PI_AD_13;
wire cordic_n_0;
wire n_845;
wire newNet_673;
wire newNet_328;
wire cordic_AddY_Add_n_7;
wire cordic_BS1_13_;
wire newNet_175;
wire newNet_532;
wire newNet_278;
wire n_429;
wire n_576;
wire cordic_AddY_MUX_1_n_26;
wire n_467;
wire cordic_Add0_MUX_0_n_27;
wire newNet_626;
wire newNet_426;
wire PO_AD_46;
wire PI_AD_8;
wire newNet_905;
wire newNet_703;
wire cordic_SH2_srl_35_26_n_17;
wire cordic_Add0_Atemp_4_;
wire cordic_AddX_Add_n_20;
wire newNet_707;
wire CoreInput_3_;
wire newNet_120;
wire n_46;
wire n_730;
wire cordic_Add0_MUX_0_n_10;
wire newNet_110;
wire CoreInput_6_;
wire cordic_AddX_Add_n_61;
wire newNet_1092;
wire newNet_1069;
wire cordic_SH1_srl_35_26_n_54;
wire newNet_130;
wire newNet_24;
wire cordic_AddY_Add_n_71;
wire n_745;
wire cordic_SH2_srl_35_26_n_144;
wire n_210;
wire newNet_1076;
wire CoreOutput_13_;
wire newNet_1086;
wire newNet_117;
wire newNet_63;
wire PI_AD_48;
wire newNet_1181;
wire n_362;
wire cordic_SH1_srl_35_26_n_9;
wire newNet_2;
wire cordic_BS2_8_;
wire newNet_247;
wire n_823;
wire newNet_739;
wire cordic_AddX_Btemp_13_;
wire n_341;
wire cordic_Add0_Btemp_3_;
wire n_541;
wire n_509;
wire newNet_593;
wire PI_AD_25;
wire cordic_SH2_srl_35_26_n_44;
wire Access_Address_1_29_;
wire n_652;
wire n_451;
wire n_737;
wire cordic_Add0_Btemp_11_;
wire cordic_SH1_srl_35_26_n_27;
wire cordic_AddY_MUX_1_n_23;
wire n_749;
wire State_1_;
wire newNet_124;
wire newNet_149;
wire newNet_375;
wire cordic_SumAngle_13_;
wire cordic_BS2_11_;
wire cordic_n_43;
wire newNet_730;
wire n_830;
wire newNet_715;
wire n_498;
wire cordic_AddY_MUX_0_n_2;
wire n_534;
wire cordic_AddX_Add_n_5;
wire PO_AD_12;
wire newNet_1043;
wire newNet_800;
wire newNet_529;
wire Access_Address_1_31_;
wire n_256;
wire newNet_1038;
wire newNet_460;
wire newNet_634;
wire newNet_272;
wire cordic_BS1_3_;
wire cordic_pla_n_3;
wire n_92;
wire cordic_Add0_Stemp_12_;
wire newNet_938;
wire newNet_670;
wire n_233;
wire cordic_Add0_n_6;
wire newNet_359;
wire n_53;
wire cordic_Add0_Add_n_38;
wire cordic_AddY_MUX_0_n_16;
wire PI_AD_51;
wire newNet_502;
wire newNet_46;
wire n_107;
wire cordic_AddX_MUX_1_n_10;
wire n_645;
wire cordic_AddX_Compl_n_7;
wire n_205;
wire n_797;
wire cordic_Add0_Atemp_1_;
wire cordic_SH1_srl_35_26_n_63;
wire PAR64_Int;
wire newNet_763;
wire cordic_AddY_MUX_0_n_22;
wire newNet_174;
wire n_231;
wire cordic_AddY_n_1;
wire newNet_277;
wire newNet_1103;
wire newNet_702;
wire newNet_492;
wire newNet_951;
wire cordic_Add0_MUX_0_n_17;
wire newNet_917;
wire newNet_891;
wire newNet_1078;
wire n_622;
wire cordic_AddY_Btemp1_12_;
wire newNet_406;
wire n_855;
wire newNet_1024;
wire cordic_Y_14_;
wire cordic_SH1_srl_35_26_n_20;
wire cordic_AddX_MUX_0_n_9;
wire n_609;
wire newNet_449;
wire cordic_AddY_MUX_0_n_11;
wire n_290;
wire n_26;
wire n_641;
wire CoreOutputReg_26_;
wire n_558;
wire cordic_AddX_MUX_1_n_24;
wire cordic_n_95;
wire newNet_464;
wire n_556;
wire PO_AD_52;
wire n_681;
wire cordic_SH2_srl_35_26_n_34;
wire CoreOutputReg_21_;
wire n_127;
wire cordic_AddY_Add_n_58;
wire newNet_313;
wire n_773;
wire cordic_Add0_n_1;
wire newNet_1193;
wire cordic_AddY_Btemp1_2_;
wire n_83;
wire newNet_8;
wire n_96;
wire newNet_645;
wire cordic_SH1_srl_35_26_n_46;
wire PI_REQ64_L;
wire PO_AD_63;
wire n_427;
wire CoreOutput_31_;
wire newNet_652;
wire cordic_SH1_srl_35_26_n_87;
wire newNet_317;
wire cordic_Add0_Compl_n_9;
wire n_519;
wire PO_AD_38;
wire cordic_AddX_MUX_0_n_2;
wire n_366;
wire newNet_74;
wire newNet_877;
wire n_208;
wire cordic_n_25;
wire newNet_1170;
wire newNet_610;
wire newNet_228;
wire cordic_SH1_srl_35_26_n_94;
wire newNet_1140;
wire PO_AD_43;
wire cordic_SH2_srl_35_26_n_112;
wire Config_Reg_29_;
wire cordic_BS1_2_;
wire n_434;
wire newNet_654;
wire cordic_AddX_Add_n_13;
wire cordic_Add0_n_15;
wire newNet_1064;
wire newNet_1052;
wire newNet_661;
wire n_405;
wire n_273;
wire newNet_1012;
wire n_258;
wire newNet_370;
wire newNet_109;
wire newNet_255;
wire cordic_Add0_Add_n_44;
wire newNet_432;
wire newNet_1169;
wire newNet_853;
wire newNet_754;
wire cordic_AddY_Add_n_30;
wire cordic_AddX_Btemp_6_;
wire newNet_50;
wire PI_AD_21;
wire newNet_56;
wire newNet_1111;
wire n_659;
wire cordic_AddX_Add_n_28;
wire newNet_681;
wire n_847;
wire PO_AD_55;
wire cordic_AddX_Atemp_2_;
wire n_810;
wire newNet_803;
wire cordic_Add0_Add_n_12;
wire n_807;
wire cordic_SH2_srl_35_26_n_51;
wire cordic_Add0_Add_n_6;
wire n_512;
wire newNet_1029;
wire cordic_AddY_Add_n_61;
wire cordic_AddX_Add_n_0;
wire n_491;
wire CoreInput_2_;
wire cordic_AddY_Btemp_8_;
wire cordic_SH1_srl_35_26_n_11;
wire n_881;
wire n_266;
wire n_34;
wire newNet_974;
wire cordic_SumAngle_12_;
wire n_976;
wire PI_AD_33;
wire cordic_AddY_MUX_1_n_0;
wire newNet_631;
wire n_389;
wire newNet_39;
wire cordic_SH1_srl_35_26_n_112;
wire newNet_1001;
wire cordic_AddX_MUX_1_n_4;
wire cordic_SH1_srl_35_26_n_18;
wire n_317;
wire newNet_1108;
wire newNet_923;
wire cordic_SH2_srl_35_26_n_69;
wire newNet_872;
wire cordic_AddY_Add_n_2;
wire newNet_549;
wire cordic_n_62;
wire cordic_SH2_srl_35_26_n_121;
wire cordic_AddY_MUX_1_n_7;
wire newNet_181;
wire cordic_n_30;
wire newNet_280;
wire cordic_n_104;
wire cordic_AddY_Compl_n_17;
wire newNet_659;
wire newNet_398;
wire newNet_216;
wire n_393;
wire cordic_SumAngle_7_;
wire newNet_1154;
wire n_299;
wire newNet_481;
wire newNet_411;
wire n_778;
wire cordic_Add0_MUX_1_n_5;
wire cordic_AddX_Add_n_76;
wire n_742;
wire cordic_SH2_srl_35_26_n_79;
wire n_310;
wire cordic_AddX_Atemp_7_;
wire n_285;
wire cordic_Add0_Stemp_11_;
wire cordic_AddX_MUX_0_n_18;
wire newNet_294;
wire n_140;
wire newNet_221;
wire n_221;
wire n_45;
wire newNet_597;
wire n_529;
wire cordic_SH2_srl_35_26_n_13;
wire newNet_435;
wire PI_AD_59;
wire cordic_AddY_n_2;
wire newNet_847;
wire n_284;
wire newNet_288;
wire cordic_Add0_Add_n_26;
wire newNet_937;
wire newNet_814;
wire newNet_628;
wire newNet_325;
wire newNet_1032;
wire newNet_565;
wire cordic_Add0_Stemp_5_;
wire cordic_n_38;
wire cordic_Add0_Add_n_71;
wire n_351;
wire cordic_SH2_srl_35_26_n_104;
wire newNet_720;
wire n_182;
wire cordic_AddX_Add_n_68;
wire newNet_768;
wire cordic_SH1_srl_35_26_n_103;
wire n_610;
wire newNet_1127;
wire n_225;
wire newNet_1054;
wire PI_AD_0;
wire cordic_AddY_Add_n_19;
wire cordic_Xsign;
wire cordic_Add0_Add_n_23;
wire n_374;
wire newNet_910;
wire newNet_299;
wire cordic_pla_n_15;
wire newNet_587;
wire cordic_AddX_Btemp1_5_;
wire n_862;
wire newNet_469;
wire newNet_164;
wire cordic_Add0_Stemp_13_;
wire cordic_SH1_srl_35_26_n_91;
wire cordic_AddY_MUX_0_n_27;
wire n_80;
wire cordic_n_56;
wire n_473;
wire n_885;
wire Par64_Sgnl;
wire cordic_AddX_Atemp_9_;
wire newNet_515;
wire n_425;
wire cordic_AddY_Add_n_26;
wire cordic_Add0_MUX_0_n_22;
wire n_581;
wire n_505;
wire newNet_729;
wire newNet_505;
wire cordic_n_59;
wire cordic_Add0_Compl_n_17;
wire n_76;
wire n_728;
wire newNet_966;
wire n_708;
wire Config_Reg_15_;
wire cordic_SH2_srl_35_26_n_2;
wire n_15;
wire newNet_445;
wire CoreOutput_6_;
wire newNet_384;
wire CoreOutput_27_;
wire n_863;
wire newNet_787;
wire PO_AD_34;
wire n_272;
wire newNet_956;
wire newNet_884;
wire n_619;
wire newNet_1122;
wire CoreInput_4_;
wire n_803;
wire cordic_AddX_Btemp_0_;
wire newNet_167;
wire n_837;
wire n_110;
wire Config_Reg_27_;
wire n_717;
wire n_382;
wire cordic_AddX_Add_n_25;
wire cordic_AddX_MUX_1_n_7;
wire n_168;
wire newNet_198;
wire PI_AD_17;
wire newNet_1198;
wire newNet_580;
wire newNet_519;
wire n_539;
wire newNet_537;
wire cordic_AddX_Compl_n_23;
wire cordic_AddX_Add_n_37;
wire cordic_AddX_MUX_0_n_23;
wire cordic_BS2_4_;
wire newNet_232;
wire cordic_AddX_Add_n_40;
wire n_244;
wire n_888;
wire newNet_679;
wire cordic_Add0_Compl_n_8;
wire n_191;
wire cordic_SH1_srl_35_26_n_122;
wire cordic_n_80;
wire cordic_AddY_Compl_n_8;
wire newNet_186;
wire cordic_AddY_MUX_0_n_5;
wire Access_Address_1_24_;
wire n_277;
wire newNet_1134;
wire n_721;
wire cordic_AddX_Compl_n_39;
wire cordic_AddY_Compl_n_35;
wire newNet_301;
wire cordic_BS2_3_;
wire n_840;
wire cordic_X_6_;
wire cordic_AddX_Add_n_49;
wire cordic_SH1_srl_35_26_n_2;
wire n_306;
wire newNet_366;
wire cordic_AddY_MUX_1_n_27;
wire n_162;
wire newNet_484;
wire n_149;
wire newNet_861;
wire n_12;
wire PI_AD_36;
wire n_169;
wire n_321;
wire n_688;
wire newNet_452;
wire cordic_X_7_;
wire cordic_n_18;
wire cordic_AddX_Add_n_55;
wire cordic_AddY_Atemp_13_;
wire n_595;
wire n_788;
wire cordic_SH1_srl_35_26_n_82;
wire cordic_AddY_Add_n_10;
wire cordic_SH2_srl_35_26_n_20;
wire cordic_AddY_Compl_n_9;
wire cordic_SH2_srl_35_26_n_8;
wire n_567;
wire newNet_613;
wire n_852;
wire cordic_Add0_Add_n_31;
wire cordic_SH2_srl_35_26_n_23;
wire newNet_734;
wire newNet_520;
wire n_411;
wire n_839;
wire newNet_1145;
wire cordic_SH1_srl_35_26_n_70;
wire cordic_SH2_srl_35_26_n_62;
wire cordic_n_111;
wire newNet_362;
wire newNet_156;
wire cordic_Add0_MUX_0_n_15;
wire n_677;
wire newNet_697;
wire n_261;
wire newNet_960;
wire newNet_574;
wire newNet_421;
wire newNet_345;
wire newNet_59;
wire n_756;
wire cordic_AddX_Add_n_46;
wire n_476;
wire cordic_AddY_Add_n_11;
wire newNet_310;
wire cordic_AddY_Atemp_2_;
wire n_869;
wire cordic_AddY_Compl_n_16;
wire cordic_AddX_Add_n_18;
wire cordic_SH1_srl_35_26_n_130;
wire n_768;
wire n_813;
wire n_872;
wire newNet_338;
wire newNet_1083;
wire newNet_749;
wire n_64;
wire cordic_Add0_MUX_0_n_5;
wire cordic_Add0_Compl_n_16;
wire newNet_1185;
wire newNet_992;
wire cordic_SH1_srl_35_26_n_121;
wire newNet_728;
wire newNet_725;
wire newNet_238;
wire n_804;
wire newNet_1046;
wire cordic_AddY_Btemp_4_;
wire newNet_1116;
wire cordic_Add0_Add_n_63;
wire cordic_Add0_MUX_0_n_23;
wire newNet_191;
wire newNet_499;
wire CoreOutputReg_28_;
wire newNet_1025;
wire cordic_AddX_Add_n_24;
wire n_438;
wire n_766;
wire newNet_361;
wire CoreOutputReg_31_;
wire cordic_n_15;
wire cordic_SH1_srl_35_26_n_99;
wire newNet_1133;
wire newNet_837;
wire newNet_711;
wire newNet_380;
wire newNet_477;
wire cordic_AddX_Add_n_1;
wire newNet_996;
wire PI_AD_29;
wire newNet_472;
wire newNet_1173;
wire newNet_397;
wire cordic_SH1_srl_35_26_n_34;
wire cordic_AddX_Stemp_0_;
wire cordic_AddX_Add_n_32;
wire newNet_323;
wire cordic_Add0_Atemp_10_;
wire PO_AD_22;
wire n_656;
wire cordic_n_108;
wire cordic_Add0_Stemp_0_;
wire newNet_211;
wire newNet_355;
wire cordic_AddY_MUX_0_n_6;
wire cordic_AddY_Add_n_65;
wire n_538;
wire newNet_1060;
wire newNet_589;
wire newNet_753;
wire cordic_AddX_Add_n_65;
wire cordic_AddY_Add_n_76;
wire cordic_AddY_Btemp1_1_;
wire n_802;
wire cordic_AddY_Atemp_4_;
wire CoreInput_12_;
wire cordic_Add0_Atemp_13_;
wire n_710;
wire newNet_911;
wire newNet_88;
wire n_11;
wire newNet_1146;
wire n_670;
wire n_667;
wire newNet_348;
wire n_662;
wire newNet_796;
wire n_515;
wire cordic_Add0_Btemp_6_;
wire newNet_550;
wire newNet_658;
wire newNet_564;
wire newNet_489;
wire n_180;
wire n_633;
wire cordic_AddY_MUX_1_n_13;
wire cordic_Add0_MUX_0_n_30;
wire newNet_773;
wire newNet_533;
wire cordic_BS1_11_;
wire cordic_AddY_Compl_n_5;
wire DWord_Trans;
wire n_612;
wire newNet_982;
wire cordic_SH1_srl_35_26_n_77;
wire n_699;
wire CoreOutputReg_27_;
wire cordic_Add0_Stemp_10_;
wire newNet_422;
wire PI_AD_55;
wire PO_AD_51;
wire cordic_Add0_n_5;
wire newNet_1036;
wire n_56;
wire newNet_1188;
wire cordic_AddX_Add_n_34;
wire cordic_Add0_Add_n_4;
wire Config_Reg_1_;
wire newNet_497;
wire cordic_Add0_MUX_0_n_2;
wire cordic_AddX_Btemp1_13_;
wire Config_Reg_2_;
wire newNet_487;
wire newNet_391;
wire cordic_Y_3_;
wire newNet_67;
wire cordic_SH2_srl_35_26_n_47;
wire cordic_AddY_MUX_1_n_22;
wire cordic_n_42;
wire newNet_841;
wire n_462;
wire cordic_SH1_srl_35_26_n_126;
wire n_103;
wire newNet_1097;
wire n_293;
wire PO_AD_8;
wire cordic_AddY_Btemp1_4_;
wire PI_AD_12;
wire n_605;
wire cordic_X_11_;
wire n_562;
wire cordic_AddY_Add_n_6;
wire newNet_441;
wire cordic_SH2_srl_35_26_n_98;
wire cordic_BS1_9_;
wire cordic_SH2_srl_35_26_n_76;
wire n_777;
wire newNet_665;
wire newNet_28;
wire n_889;
wire cordic_Angle_15_;
wire cordic_AddX_Btemp_1_;
wire newNet_693;
wire PO_STOP_L;
wire newNet_480;
wire cordic_BS2_12_;
wire newNet_548;
wire newNet_1138;
wire newNet_525;
wire cordic_n_37;
wire newNet_1020;
wire PO_AD_25;
wire newNet_514;
wire newNet_379;
wire n_414;
wire n_328;
wire cordic_SH1_srl_35_26_n_32;
wire newNet_1107;
wire CoreOutputReg_32_;
wire newNet_810;
wire newNet_921;
wire cordic_AddX_n_3;
wire newNet_553;
wire cordic_BS1_0_;
wire n_409;
wire cordic_AddX_Add_n_17;
wire cordic_AddY_n_5;
wire newNet_692;
wire n_866;
wire cordic_AddX_Compl_n_15;
wire cordic_SH2_srl_35_26_n_18;
wire n_577;
wire cordic_SH1_srl_35_26_n_83;
wire newNet_843;
wire newNet_386;
wire n_252;
wire cordic_SH1_srl_35_26_n_23;
wire cordic_AddX_MUX_0_n_12;
wire n_470;
wire cordic_AddX_Atemp_3_;
wire n_448;
wire newNet_248;
wire newNet_12;
wire PI_PAR64;
wire newNet_948;
wire newNet_1194;
wire newNet_1057;
wire CoreInput_13_;
wire CBE_par_1_;
wire newNet_14;
wire cordic_SH2_srl_35_26_n_55;
wire cordic_AddX_MUX_1_n_26;
wire cordic_tanangle_10_;
wire newNet_419;
wire n_648;
wire newNet_970;
wire newNet_242;
wire n_421;
wire cordic_n_99;
wire cordic_BS1_14_;
wire cordic_pla_n_25;
wire cordic_AddX_Atemp_0_;
wire newNet_133;
wire cordic_AddY_Add_n_37;
wire newNet_163;
wire cordic_SH1_srl_35_26_n_43;
wire n_38;
wire cordic_pla_n_31;
wire newNet_98;
wire n_454;
wire newNet_206;
wire cordic_AddX_Compl_n_14;
wire CoreOutput_16_;
wire cordic_n_71;
wire cordic_SH1_srl_35_26_n_116;
wire cordic_Add0_Add_n_17;
wire n_494;
wire n_433;
wire newNet_644;
wire n_267;
wire cordic_Add0_Add_n_75;
wire newNet_1174;
wire cordic_SH1_srl_35_26_n_13;
wire cordic_AddX_Atemp_4_;
wire cordic_pla_n_23;
wire cordic_Add0_Add_n_15;
wire cordic_Add0_Stemp_7_;
wire PO_AD_29;
wire n_603;
wire n_178;
wire cordic_SH2_srl_35_26_n_131;
wire n_586;
wire cordic_AddX_MUX_0_n_19;
wire n_87;
wire newNet_807;
wire newNet_153;
wire cordic_Add0_Compl_n_3;
wire cordic_SH2_srl_35_26_n_40;
wire cordic_iteration_0_;
wire n_174;
wire newNet_436;
wire newNet_979;
wire newNet_760;
wire cordic_AddY_MUX_0_n_30;
wire n_875;
wire n_5;
wire cordic_Add0_Add_n_7;
wire CoreOutput_29_;
wire newNet_262;
wire newNet_71;
wire newNet_405;
wire newNet_463;
wire newNet_401;
wire n_385;
wire cordic_n_50;
wire newNet_676;
wire n_487;
wire newNet_617;
wire newNet_686;
wire newNet_1015;
wire newNet_225;
wire cordic_AddX_Btemp1_11_;
wire newNet_758;
wire n_84;
wire n_892;
wire newNet_172;
wire cordic_n_69;
wire newNet_906;
wire cordic_n_1;
wire newNet_576;
wire newNet_465;
wire cordic_SumAngle_3_;
wire cordic_AddY_Compl_n_12;
wire cordic_Add0_Compl_n_43;
wire cordic_SH2_srl_35_26_n_65;
wire n_899;
wire newNet_81;
wire n_185;
wire CBE_par_3_;
wire newNet_457;
wire newNet_820;
wire cordic_AddY_Add_n_55;
wire newNet_1093;
wire newNet_888;
wire n_113;
wire newNet_944;
wire cordic_SH1_srl_35_26_n_131;
wire cordic_n_89;
wire cordic_AddX_Btemp_5_;
wire newNet_621;
wire n_571;
wire newNet_547;
wire n_153;
wire cordic_pla_n_11;
wire newNet_250;
wire cordic_AddX_Btemp1_14_;
wire cordic_AddY_MUX_0_n_7;
wire cordic_SH1_srl_35_26_n_53;
wire n_59;
wire cordic_SH2_srl_35_26_n_86;
wire CoreOutput_1_;
wire newNet_1066;
wire newNet_55;
wire n_128;
wire cordic_AddY_Btemp_7_;
wire Access_Address_1_23_;
wire newNet_1011;
wire cordic_AddY_MUX_0_n_26;
wire n_355;
wire newNet_858;
wire cordic_AddY_Add_n_28;
wire n_229;
wire n_350;
wire cordic_AddX_Btemp1_2_;
wire n_846;
wire Config_Reg_4_;
wire cordic_AddX_Btemp1_10_;
wire cordic_Add0_MUX_0_n_26;
wire PI_AD_5;
wire newNet_606;
wire CoreOutputReg_4_;
wire cordic_SH2_srl_35_26_n_24;
wire n_392;
wire newNet_284;
wire newNet_102;
wire cordic_n_121;
wire newNet_1112;
wire newNet_334;
wire cordic_X_4_;
wire cordic_AddX_Add_n_21;
wire newNet_1072;
wire PO_AD_49;
wire newNet_706;
wire cordic_BS1_7_;
wire newNet_538;
wire CoreInput_10_;
wire CoreOutput_3_;
wire newNet_33;
wire cordic_SH2_srl_35_26_n_14;
wire newNet_291;
wire newNet_1153;
wire n_625;
wire PO_AD_47;
wire cordic_SumAngle_8_;
wire newNet_827;
wire CoreOutput_15_;
wire n_466;
wire newNet_425;
wire cordic_Add0_Add_n_50;
wire PO_AD_19;
wire newNet_764;
wire n_684;
wire n_753;
wire newNet_740;
wire n_547;
wire newNet_329;
wire n_134;
wire cordic_Add0_n_12;
wire newNet_350;
wire cordic_SH2_srl_35_26_n_41;
wire n_281;
wire n_49;
wire newNet_896;
wire n_545;
wire cordic_AddY_Add_n_47;
wire n_483;
wire newNet_416;
wire newNet_561;
wire cordic_AddX_Btemp1_6_;
wire cordic_n_76;
wire cordic_n_10;
wire newNet_1087;
wire cordic_AddX_MUX_0_n_21;
wire cordic_AddY_Stemp_0_;
wire cordic_AddX_MUX_0_n_8;
wire CoreOutputReg_1_;
wire cordic_AddX_Stemp_5_;
wire newNet_1158;
wire newNet_60;
wire cordic_SH2_srl_35_26_n_38;
wire newNet_826;
wire newNet_716;
wire newNet_44;
wire cordic_AddX_MUX_1_n_19;
wire newNet_932;
wire newNet_306;
wire cordic_SH2_srl_35_26_n_52;
wire n_106;
wire newNet_584;
wire cordic_BS1_6_;
wire n_197;
wire newNet_918;
wire cordic_Add0_Compl_n_11;
wire newNet_511;
wire newNet_1141;
wire newNet_64;
wire PO_PAR64;
wire n_123;
wire newNet_78;
wire cordic_SH1_srl_35_26_n_66;
wire newNet_1091;
wire newNet_989;
wire cordic_SH2_srl_35_26_n_30;
wire PI_CBE_L_7;
wire cordic_SH2_srl_35_26_n_120;
wire cordic_n_116;
wire cordic_BS1_1_;
wire newNet_860;
wire cordic_AddX_Btemp_4_;
wire cordic_AddX_Y_1;
wire PI_AD_22;
wire Config_Reg_20_;
wire cordic_SH1_srl_35_26_n_37;
wire cordic_n_60;
wire newNet_865;
wire newNet_91;
wire n_31;
wire newNet_332;
wire n_91;
wire cordic_AddX_Add_n_70;
wire n_397;
wire n_202;
wire n_525;
wire TAR_TRI_D;
wire newNet_955;
wire n_72;
wire cordic_AddX_MUX_1_n_1;
wire cordic_SH2_srl_35_26_n_27;
wire CoreOutput_24_;
wire cordic_AddY_Compl_n_13;
wire n_79;
wire cordic_AddX_Add_n_52;
wire DevSel_Wait_Cnt_0_;
wire n_19;
wire cordic_n_34;
wire newNet_194;
wire cordic_SH2_srl_35_26_n_92;
wire cordic_Add0_Add_n_57;
wire cordic_Add0_MUX_1_n_4;
wire cordic_AddX_MUX_0_n_26;
wire cordic_AddY_MUX_1_n_3;
wire newNet_962;
wire n_829;
wire cordic_AddY_Add_n_16;
wire newNet_783;
wire n_378;
wire newNet_559;
wire cordic_Add0_MUX_0_n_6;
wire cordic_n_101;
wire cordic_AddX_MUX_0_n_6;
wire n_608;
wire PI_CBE_L_1;
wire n_798;
wire cordic_n_100;
wire n_784;
wire n_526;
wire n_732;
wire Config_Reg_18_;
wire newNet_341;
wire cordic_SH2_srl_35_26_n_125;

// Start cells
BUF_X2 newInst_312 ( .a(newNet_311), .o(newNet_312) );
NOR2_Z1 g15431 ( .a(n_210), .b(n_135), .o(n_273) );
NAND2_Z01 cordic_AddX_MUX_0_g281 ( .a(cordic_AddX_MUX_0_n_24), .b(cordic_AddX_MUX_0_n_8), .o(cordic_AddX_Atemp_7_) );
BUF_X2 newInst_1154 ( .a(newNet_423), .o(newNet_1154) );
AND2_X1 cordic_AddX_Compl_g349 ( .a(cordic_AddX_Compl_n_31), .b(cordic_AddX_Compl_n_15), .o(cordic_AddX_Compl_n_33) );
INV_X1 g15651 ( .a(PO_SERR_L), .o(n_14) );
NAND2_Z01 g15249 ( .a(n_313), .b(n_314), .o(n_411) );
NAND2_Z01 g14930 ( .a(n_591), .b(n_521), .o(n_644) );
NAND2_Z01 cordic_SH1_srl_35_26_g1113 ( .a(cordic_SH1_srl_35_26_n_126), .b(cordic_iteration_3_), .o(cordic_SH1_srl_35_26_n_139) );
NAND2_Z01 cordic_Add0_Add_g675 ( .a(cordic_Add0_Stemp_0_), .b(cordic_Add0_Add_n_0), .o(cordic_Add0_Add_n_32) );
BUF_X2 newInst_540 ( .a(newNet_539), .o(newNet_540) );
NAND2_Z01 g14897 ( .a(n_624), .b(n_553), .o(n_677) );
BUF_X2 newInst_1096 ( .a(newNet_848), .o(newNet_1096) );
BUF_X2 newInst_224 ( .a(newNet_223), .o(newNet_224) );
NOR2_Z1 g13447 ( .a(n_802), .b(n_710), .o(n_835) );
BUF_X2 newInst_378 ( .a(newNet_377), .o(newNet_378) );
NAND2_Z01 cordic_Add0_MUX_0_g272 ( .a(cordic_tanangle_8_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_31) );
NAND2_Z01 g15378 ( .a(n_214), .b(CoreOutputReg_25_), .o(n_283) );
BUF_X2 newInst_785 ( .a(newNet_784), .o(newNet_785) );
BUF_X2 newInst_569 ( .a(newNet_568), .o(newNet_569) );
fflopd cordic_X_reg_8_ ( .CK(newNet_16), .D(cordic_n_30), .Q(cordic_X_8_) );
NAND2_Z01 g14939 ( .a(n_582), .b(n_510), .o(n_635) );
NAND3_Z1 g14819 ( .a(n_689), .b(n_691), .c(n_155), .o(n_700) );
NOR2_Z1 g15311 ( .a(n_271), .b(n_127), .o(n_382) );
XOR2_X1 cordic_AddY_Compl_g364 ( .a(cordic_AddY_Compl_n_11), .b(cordic_AddY_Compl_n_1), .o(CoreOutput_1_) );
NAND2_Z01 cordic_AddY_MUX_0_g281 ( .a(cordic_AddY_MUX_0_n_24), .b(cordic_AddY_MUX_0_n_8), .o(cordic_AddY_Atemp_7_) );
NAND2_Z01 cordic_Add0_Add_g650 ( .a(cordic_Add0_Add_n_56), .b(cordic_Add0_Add_n_21), .o(cordic_Add0_Add_n_57) );
fflopd CoreInput_reg_1_ ( .CK(newNet_775), .D(n_648), .Q(CoreInput_1_) );
BUF_X2 newInst_369 ( .a(newNet_368), .o(newNet_369) );
AND2_X1 cordic_Add0_Compl_g345 ( .a(cordic_Add0_Compl_n_35), .b(cordic_Add0_Compl_n_3), .o(cordic_Add0_Compl_n_37) );
BUF_X2 newInst_1068 ( .a(newNet_1067), .o(newNet_1068) );
NAND2_Z01 g14922 ( .a(n_599), .b(n_529), .o(n_652) );
NAND2_Z01 g13491 ( .a(n_724), .b(n_763), .o(n_793) );
BUF_X2 newInst_410 ( .a(newNet_409), .o(newNet_410) );
XOR2_X1 cordic_AddY_Add_g705 ( .a(cordic_AddY_Btemp1_11_), .b(cordic_AddY_Atemp_11_), .o(cordic_AddY_Add_n_29) );
NAND3_Z1 g15441 ( .a(n_106), .b(n_6), .c(n_116), .o(n_268) );
NAND2_Z01 g14978 ( .a(n_571), .b(CoreInput_13_), .o(n_599) );
NAND2_Z01 cordic_AddX_Add_g702 ( .a(cordic_AddX_Add_n_16), .b(cordic_AddX_Y_2), .o(cordic_AddX_Add_n_32) );
NAND2_Z01 cordic_pla_g297 ( .a(cordic_iteration_1_), .b(cordic_iteration_0_), .o(cordic_pla_n_14) );
BUF_X2 newInst_667 ( .a(newNet_666), .o(newNet_667) );
INV_X1 cordic_g490 ( .a(CoreOutput_9_), .o(cordic_n_17) );
NOR2_Z1 cordic_g447 ( .a(cordic_n_27), .b(Issue_Rst), .o(cordic_n_60) );
NAND2_Z01 cordic_SH2_srl_35_26_g1133 ( .a(cordic_SH2_srl_35_26_n_98), .b(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_119) );
NAND2_Z01 cordic_AddX_Add_g679 ( .a(cordic_AddX_Add_n_53), .b(cordic_AddX_Add_n_15), .o(cordic_AddX_Add_n_55) );
XNOR2_X1 cordic_AddX_Compl_g379 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_6_), .o(cordic_AddX_Compl_n_4) );
NAND2_Z01 cordic_Add0_MUX_0_g298 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_12_), .o(cordic_Add0_MUX_0_n_5) );
NAND2_Z01 cordic_SH2_srl_35_26_g1137 ( .a(cordic_SH2_srl_35_26_n_97), .b(cordic_SH2_srl_35_26_n_18), .o(cordic_SH2_srl_35_26_n_115) );
NAND2_Z01 g14971 ( .a(n_572), .b(Config_Reg_7_), .o(n_606) );
NAND2_Z01 g15265 ( .a(n_264), .b(n_265), .o(n_395) );
BUF_X2 newInst_1107 ( .a(newNet_1106), .o(newNet_1107) );
BUF_X2 newInst_1048 ( .a(newNet_104), .o(newNet_1048) );
BUF_X2 newInst_143 ( .a(newNet_142), .o(newNet_143) );
NOR2_Z1 g13431 ( .a(n_782), .b(n_710), .o(n_851) );
BUF_X2 newInst_1168 ( .a(newNet_1167), .o(newNet_1168) );
NAND2_Z01 g15267 ( .a(n_260), .b(n_261), .o(n_393) );
INV_X1 cordic_SH1_srl_35_26_g1250 ( .a(cordic_iteration_2_), .o(cordic_SH1_srl_35_26_n_2) );
NAND2_Z01 cordic_Add0_MUX_0_g282 ( .a(cordic_tanangle_9_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_21) );
NAND2_Z01 cordic_AddY_MUX_0_g286 ( .a(cordic_AddY_MUX_0_n_21), .b(cordic_AddY_MUX_0_n_4), .o(cordic_AddY_Atemp_5_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1120 ( .a(cordic_SH2_srl_35_26_n_125), .b(cordic_SH2_srl_35_26_n_121), .o(cordic_SH2_srl_35_26_n_132) );
NAND2_Z01 cordic_AddX_MUX_0_g313 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_7_), .o(cordic_AddX_MUX_0_n_8) );
BUF_X2 newInst_693 ( .a(newNet_692), .o(newNet_693) );
NAND2_Z01 cordic_AddY_MUX_1_g298 ( .a(cordic_AddY_Y_1), .b(cordic_Y_11_), .o(cordic_AddY_MUX_1_n_23) );
NAND2_Z01 g13473 ( .a(n_747), .b(n_775), .o(n_811) );
NAND2_Z01 cordic_SH1_srl_35_26_g1224 ( .a(cordic_iteration_0_), .b(cordic_Y_9_), .o(cordic_SH1_srl_35_26_n_28) );
AND2_X1 cordic_g473 ( .a(CoreOutput_28_), .b(Issue_Rst), .o(cordic_n_34) );
BUF_X2 newInst_7 ( .a(newNet_6), .o(newNet_7) );
fflopd Config_Reg_reg_23_ ( .CK(newNet_952), .D(n_673), .Q(Config_Reg_23_) );
NAND2_Z01 cordic_AddY_Add_g694 ( .a(cordic_AddY_Add_n_38), .b(cordic_AddY_Add_n_3), .o(cordic_AddY_Add_n_40) );
NAND2_Z01 g15072 ( .a(n_473), .b(PI_AD_4), .o(n_536) );
BUF_X2 newInst_509 ( .a(newNet_508), .o(newNet_509) );
BUF_X2 newInst_173 ( .a(newNet_44), .o(newNet_173) );
BUF_X2 newInst_839 ( .a(newNet_838), .o(newNet_839) );
BUF_X2 newInst_108 ( .a(newNet_107), .o(newNet_108) );
NAND2_Z01 g15326 ( .a(n_184), .b(PI_AD_19), .o(n_335) );
INV_X1 g13576 ( .a(Par_Sgnl), .o(n_711) );
NOR2_Z1 g13454 ( .a(n_791), .b(n_710), .o(n_828) );
AND2_X1 g60 ( .a(n_831), .b(n_856), .o(PO_AD_4) );
NOR2_Z1 g15428 ( .a(n_189), .b(n_8), .o(n_226) );
NAND2_Z01 g13528 ( .a(Idsel), .b(Config_Reg_25_), .o(n_758) );
NAND2_Z01 cordic_SH2_srl_35_26_g1168 ( .a(cordic_SH2_srl_35_26_n_51), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_84) );
NAND2_Z01 g14983 ( .a(n_571), .b(CoreInput_2_), .o(n_594) );
fflopd Access_Address_1_reg_25_ ( .CK(newNet_1151), .D(n_483), .Q(Access_Address_1_25_) );
BUF_X2 newInst_1147 ( .a(newNet_1146), .o(newNet_1147) );
fflopd cordic_iteration_reg_3_ ( .CK(newNet_300), .D(cordic_n_123), .Q(cordic_iteration_3_) );
BUF_X2 newInst_754 ( .a(newNet_753), .o(newNet_754) );
XOR2_X1 g15587 ( .a(PI_AD_21), .b(PI_AD_9), .o(n_78) );
BUF_X2 newInst_519 ( .a(newNet_518), .o(newNet_519) );
fflopd CoreInput_reg_12_ ( .CK(newNet_804), .D(n_653), .Q(CoreInput_12_) );
NAND2_Z01 g15099 ( .a(n_473), .b(PI_AD_9), .o(n_509) );
BUF_X2 newInst_762 ( .a(newNet_761), .o(newNet_762) );
AND3_X1 g14833 ( .a(n_139), .b(n_685), .c(n_131), .o(n_687) );
XOR2_X1 cordic_AddY_Compl_g348 ( .a(cordic_AddY_Compl_n_31), .b(cordic_AddY_Compl_n_15), .o(CoreOutput_9_) );
NAND2_Z01 g15342 ( .a(cordic_AddY_Stemp_0_), .b(n_2), .o(n_319) );
BUF_X2 newInst_1190 ( .a(newNet_1189), .o(newNet_1190) );
AND2_X1 g15568 ( .a(n_37), .b(State_1_), .o(n_108) );
BUF_X2 newInst_644 ( .a(newNet_643), .o(newNet_644) );
fflopd CoreOutputReg_reg_26_ ( .CK(newNet_623), .D(n_395), .Q(CoreOutputReg_26_) );
NAND2_Z01 g13495 ( .a(n_735), .b(n_754), .o(n_789) );
NAND2_Z01 cordic_AddY_MUX_0_g306 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_9_), .o(cordic_AddY_MUX_0_n_15) );
AND2_X1 g15439 ( .a(n_6), .b(n_133), .o(n_220) );
fflopd CoreOutputReg_reg_33_ ( .CK(newNet_589), .D(n_387), .Q(CoreOutputReg_33_) );
BUF_X2 newInst_434 ( .a(newNet_433), .o(newNet_434) );
INV_X2 newInst_892 ( .a(newNet_891), .o(newNet_892) );
NAND2_Z01 cordic_Add0_MUX_0_g285 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_2_), .o(cordic_Add0_MUX_0_n_18) );
INV_X1 g15384 ( .a(n_266), .o(n_267) );
XOR2_X1 cordic_Add0_Compl_g356 ( .a(cordic_Add0_Compl_n_23), .b(cordic_Add0_Compl_n_5), .o(cordic_SumAngle_5_) );
INV_X1 g15641 ( .a(Burst_Trans), .o(n_24) );
NAND2_Z01 g15360 ( .a(cordic_AddX_Stemp_0_), .b(n_2), .o(n_301) );
BUF_X2 newInst_702 ( .a(newNet_467), .o(newNet_702) );
NAND2_Z01 g15300 ( .a(n_266), .b(DevSel_Wait_Cnt_0_), .o(n_355) );
NOR2_Z1 cordic_SH2_srl_35_26_g1246 ( .a(cordic_SH2_srl_35_26_n_2), .b(cordic_iteration_3_), .o(cordic_SH2_srl_35_26_n_21) );
BUF_X2 newInst_690 ( .a(newNet_689), .o(newNet_690) );
INV_Z1 cordic_AddY_MUX_1_g321 ( .a(cordic_AddY_Y_1), .o(cordic_AddY_MUX_1_n_0) );
AND2_X1 cordic_pla_g287 ( .a(cordic_pla_n_9), .b(cordic_pla_n_4), .o(cordic_pla_n_24) );
fflopd CoreOutputReg_reg_17_ ( .CK(newNet_687), .D(n_405), .Q(CoreOutputReg_17_) );
BUF_X2 newInst_878 ( .a(newNet_877), .o(newNet_878) );
BUF_X2 newInst_1006 ( .a(newNet_1005), .o(newNet_1006) );
BUF_X2 newInst_20 ( .a(newNet_19), .o(newNet_20) );
XOR2_X1 cordic_Add0_Add_g667 ( .a(cordic_Add0_Add_n_38), .b(cordic_Add0_Add_n_23), .o(cordic_Add0_Stemp_3_) );
NAND2_Z01 g15270 ( .a(n_254), .b(n_255), .o(n_390) );
BUF_X2 newInst_944 ( .a(newNet_429), .o(newNet_944) );
BUF_X2 newInst_1166 ( .a(newNet_1165), .o(newNet_1166) );
BUF_X2 newInst_926 ( .a(newNet_925), .o(newNet_926) );
NAND2_Z01 cordic_AddX_MUX_1_g317 ( .a(cordic_BS1_5_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_4) );
AND2_X1 g361 ( .a(n_851), .b(n_856), .o(PO_AD_33) );
BUF_X2 newInst_1197 ( .a(newNet_1196), .o(newNet_1197) );
INV_X1 g15647 ( .a(Access_Type_1_1_), .o(n_18) );
NAND2_Z01 cordic_SH2_srl_35_26_g1191 ( .a(cordic_SH2_srl_35_26_n_56), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_61) );
XOR2_X1 cordic_AddX_Add_g711 ( .a(cordic_AddX_Btemp1_13_), .b(cordic_AddX_Atemp_13_), .o(cordic_AddX_Add_n_23) );
NAND2_Z01 cordic_SH1_srl_35_26_g1199 ( .a(cordic_SH1_srl_35_26_n_17), .b(cordic_SH1_srl_35_26_n_29), .o(cordic_SH1_srl_35_26_n_53) );
BUF_X2 newInst_584 ( .a(newNet_583), .o(newNet_584) );
BUF_X2 newInst_700 ( .a(newNet_699), .o(newNet_700) );
NOR2_Z1 cordic_SH1_srl_35_26_g1211 ( .a(cordic_SH1_srl_35_26_n_19), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_43) );
XOR2_X1 cordic_AddX_Add_g717 ( .a(cordic_AddX_Btemp1_8_), .b(cordic_AddX_Atemp_8_), .o(cordic_AddX_Add_n_17) );
BUF_X2 newInst_647 ( .a(newNet_646), .o(newNet_647) );
NAND2_Z01 g15348 ( .a(CoreOutput_12_), .b(n_2), .o(n_313) );
AND2_X1 g15567 ( .a(n_50), .b(DevSel_Wait_Cnt_0_), .o(n_109) );
BUF_X2 newInst_298 ( .a(newNet_297), .o(newNet_298) );
BUF_X2 newInst_402 ( .a(newNet_401), .o(newNet_402) );
NAND2_Z01 g15133 ( .a(n_435), .b(n_383), .o(n_478) );
NAND2_Z01 cordic_SH2_srl_35_26_g1245 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_14_), .o(cordic_SH2_srl_35_26_n_4) );
NOR2_Z1 g15482 ( .a(n_158), .b(n_46), .o(n_186) );
XOR2_X1 cordic_AddY_Add_g717 ( .a(cordic_AddY_Btemp1_8_), .b(cordic_AddY_Atemp_8_), .o(cordic_AddY_Add_n_17) );
NAND2_Z01 cordic_Add0_MUX_1_g255 ( .a(cordic_Add0_MUX_1_n_13), .b(cordic_Add0_MUX_1_n_18), .o(cordic_Add0_Btemp_13_) );
NAND2_Z01 cordic_AddX_MUX_1_g281 ( .a(cordic_AddX_MUX_1_n_8), .b(cordic_AddX_MUX_1_n_24), .o(cordic_AddX_Btemp_7_) );
BUF_X2 newInst_923 ( .a(newNet_922), .o(newNet_923) );
BUF_X2 newInst_1017 ( .a(newNet_1016), .o(newNet_1017) );
BUF_X2 newInst_10 ( .a(newNet_9), .o(newNet_10) );
BUF_X2 newInst_1057 ( .a(newNet_1056), .o(newNet_1057) );
BUF_X2 newInst_216 ( .a(newNet_215), .o(newNet_216) );
BUF_X2 newInst_168 ( .a(newNet_167), .o(newNet_168) );
NAND2_Z01 cordic_pla_g283 ( .a(cordic_pla_n_9), .b(cordic_pla_n_11), .o(cordic_pla_n_31) );
NAND2_Z01 cordic_AddY_MUX_0_g294 ( .a(cordic_BS2_1_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_27) );
NOR2_Z1 g13442 ( .a(n_808), .b(n_710), .o(n_840) );
NAND2_Z01 g15062 ( .a(n_473), .b(PI_AD_7), .o(n_546) );
fflopd Access_Address_1_reg_31_ ( .CK(newNet_1121), .D(n_471), .Q(Access_Address_1_31_) );
BUF_X2 newInst_1019 ( .a(newNet_1018), .o(newNet_1019) );
fflopd cordic_X_reg_5_ ( .CK(newNet_126), .D(cordic_n_49), .Q(cordic_X_5_) );
AND2_X1 g15106 ( .a(n_465), .b(n_497), .o(n_502) );
NAND2_Z01 cordic_SH1_srl_35_26_g1233 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_8_), .o(cordic_SH1_srl_35_26_n_16) );
NAND2_Z01 cordic_g398 ( .a(cordic_n_67), .b(cordic_n_89), .o(cordic_n_109) );
AND4_X1 g15021 ( .a(Access_Address_1_25_), .b(n_21), .c(n_437), .d(Access_Address_1_24_), .o(n_561) );
NAND2_Z01 g13480 ( .a(n_734), .b(n_770), .o(n_804) );
XOR2_X1 g13408 ( .a(n_871), .b(PO_AD_25), .o(n_872) );
BUF_X2 newInst_505 ( .a(newNet_504), .o(newNet_505) );
XNOR2_X1 cordic_Add0_Compl_g370 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_12_), .o(cordic_Add0_Compl_n_12) );
fflopd DevSel_Wait_Cnt_reg_1_ ( .CK(newNet_500), .D(n_487), .Q(DevSel_Wait_Cnt_1_) );
BUF_X2 newInst_681 ( .a(newNet_680), .o(newNet_681) );
BUF_X2 newInst_19 ( .a(newNet_18), .o(newNet_19) );
NAND2_Z01 cordic_AddY_MUX_0_g288 ( .a(cordic_AddY_MUX_0_n_17), .b(cordic_AddY_MUX_0_n_16), .o(cordic_AddY_Atemp_3_) );
AND2_X1 cordic_AddX_g64 ( .a(cordic_AddX_Y_3), .b(cordic_AddX_n_1), .o(cordic_AddX_n_3) );
NAND2_Z01 cordic_SH2_srl_35_26_g1171 ( .a(cordic_SH2_srl_35_26_n_46), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_81) );
BUF_X2 newInst_488 ( .a(newNet_487), .o(newNet_488) );
NAND2_Z01 cordic_AddY_Add_g697 ( .a(cordic_AddY_Add_n_35), .b(cordic_AddY_Add_n_2), .o(cordic_AddY_Add_n_37) );
BUF_X2 newInst_274 ( .a(newNet_273), .o(newNet_274) );
AND2_X1 g339 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_55) );
BUF_X2 newInst_197 ( .a(newNet_196), .o(newNet_197) );
BUF_X2 newInst_340 ( .a(newNet_339), .o(newNet_340) );
INV_X1 cordic_SH1_srl_35_26_g1125 ( .a(cordic_SH1_srl_35_26_n_126), .o(cordic_SH1_srl_35_26_n_127) );
NAND2_Z01 cordic_Add0_MUX_0_g275 ( .a(cordic_tanangle_0_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_28) );
NAND2_Z01 cordic_g393 ( .a(cordic_n_72), .b(cordic_n_94), .o(cordic_n_114) );
NAND2_Z01 g15119 ( .a(n_447), .b(PI_PAR64), .o(n_490) );
BUF_X2 newInst_933 ( .a(newNet_932), .o(newNet_933) );
NOR2_Z1 cordic_g460 ( .a(cordic_n_6), .b(Issue_Rst), .o(cordic_n_47) );
BUF_X2 newInst_843 ( .a(newNet_842), .o(newNet_843) );
NAND2_Z01 g15083 ( .a(n_494), .b(PI_AD_1), .o(n_525) );
BUF_X2 newInst_295 ( .a(newNet_294), .o(newNet_295) );
NAND2_Z01 cordic_SH2_srl_35_26_g1189 ( .a(cordic_SH2_srl_35_26_n_45), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_63) );
NAND2_Z01 g15053 ( .a(n_473), .b(PI_AD_18), .o(n_555) );
NAND2_Z01 cordic_Add0_MUX_1_g270 ( .a(cordic_AngleCin), .b(cordic_Angle_8_), .o(cordic_Add0_MUX_1_n_31) );
AND2_X1 g15221 ( .a(n_386), .b(RESET), .o(n_433) );
INV_X2 newInst_375 ( .a(newNet_374), .o(newNet_375) );
BUF_X2 newInst_997 ( .a(newNet_996), .o(newNet_997) );
NAND2_Z01 cordic_AddY_Add_g672 ( .a(cordic_AddY_Add_n_61), .b(cordic_AddY_Add_n_27), .o(cordic_AddY_Add_n_62) );
BUF_X2 newInst_652 ( .a(newNet_651), .o(newNet_652) );
NAND2_Z01 g15151 ( .a(n_445), .b(n_384), .o(n_461) );
NAND2_Z01 cordic_AddX_MUX_1_g302 ( .a(cordic_AddX_Y_1), .b(cordic_X_10_), .o(cordic_AddX_MUX_1_n_19) );
NAND2_Z01 cordic_SH2_srl_35_26_g1225 ( .a(cordic_iteration_0_), .b(cordic_X_7_), .o(cordic_SH2_srl_35_26_n_27) );
BUF_X2 newInst_42 ( .a(newNet_41), .o(newNet_42) );
BUF_X2 newInst_716 ( .a(newNet_715), .o(newNet_716) );
BUF_X2 newInst_4 ( .a(newNet_3), .o(newNet_4) );
fflopd cordic_Angle_reg_12_ ( .CK(newNet_254), .D(cordic_n_114), .Q(cordic_Angle_12_) );
NOR2_Z1 g15447 ( .a(n_157), .b(n_15), .o(n_207) );
fflopd cordic_X_reg_14_ ( .CK(newNet_153), .D(cordic_n_55), .Q(cordic_X_14_) );
NOR2_Z1 cordic_SH2_srl_35_26_g1144 ( .a(cordic_SH2_srl_35_26_n_94), .b(cordic_SH2_srl_35_26_n_19), .o(cordic_BS2_12_) );
BUF_X2 newInst_808 ( .a(newNet_807), .o(newNet_808) );
NAND2_Z01 cordic_Add0_Add_g674 ( .a(cordic_Add0_Add_n_32), .b(cordic_Add0_Add_n_18), .o(cordic_Add0_Add_n_33) );
BUF_X2 newInst_102 ( .a(newNet_101), .o(newNet_102) );
NAND2_Z01 cordic_AddX_Add_g682 ( .a(cordic_AddX_Add_n_50), .b(cordic_AddX_Add_n_0), .o(cordic_AddX_Add_n_52) );
XOR2_X1 g15606 ( .a(PI_AD_54), .b(PI_AD_36), .o(n_59) );
NAND2_Z01 g13555 ( .a(n_712), .b(CoreOutputReg_8_), .o(n_732) );
fflopd CoreOutputReg_reg_30_ ( .CK(newNet_606), .D(n_390), .Q(CoreOutputReg_30_) );
NAND2_Z01 cordic_AddY_MUX_1_g293 ( .a(cordic_AddY_Y_1), .b(cordic_Y_12_), .o(cordic_AddY_MUX_1_n_28) );
NAND2_Z01 g15387 ( .a(n_214), .b(CoreOutputReg_27_), .o(n_263) );
XNOR2_X1 cordic_Add0_Compl_g379 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_6_), .o(cordic_Add0_Compl_n_4) );
BUF_X2 newInst_1108 ( .a(newNet_1107), .o(newNet_1108) );
NAND2_Z01 cordic_Add0_MUX_1_g284 ( .a(cordic_AngleCin), .b(cordic_Angle_2_), .o(cordic_Add0_MUX_1_n_17) );
NAND3_Z1 g15312 ( .a(n_187), .b(n_276), .c(n_22), .o(n_347) );
NAND2_Z01 cordic_SH2_srl_35_26_g1155 ( .a(cordic_SH2_srl_35_26_n_85), .b(cordic_SH2_srl_35_26_n_71), .o(cordic_SH2_srl_35_26_n_98) );
NAND2_Z01 g13526 ( .a(Idsel), .b(Config_Reg_26_), .o(n_760) );
NAND2_Z01 g15077 ( .a(n_4), .b(PI_AD_11), .o(n_531) );
NAND2_Z01 g14809 ( .a(n_705), .b(n_104), .o(n_707) );
BUF_X2 newInst_233 ( .a(newNet_232), .o(newNet_233) );
NAND2_Z01 cordic_g418 ( .a(Issue_Rst), .b(CoreInput_3_), .o(cordic_n_89) );
NAND2_Z01 cordic_SH2_srl_35_26_g1227 ( .a(cordic_iteration_0_), .b(cordic_X_6_), .o(cordic_SH2_srl_35_26_n_25) );
AND2_X1 g346 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_48) );
BUF_X2 newInst_512 ( .a(newNet_511), .o(newNet_512) );
INV_X1 cordic_g506 ( .a(CoreOutput_21_), .o(cordic_n_1) );
NAND2_Z01 g15283 ( .a(n_237), .b(n_218), .o(n_372) );
BUF_X2 newInst_530 ( .a(newNet_529), .o(newNet_530) );
XOR2_X1 g15163 ( .a(n_338), .b(n_339), .o(n_449) );
XNOR2_X1 cordic_AddY_g2 ( .a(cordic_AngleCin), .b(cordic_Ysign), .o(cordic_AddY_n_0) );
BUF_X2 newInst_883 ( .a(newNet_882), .o(newNet_883) );
NAND2_Z01 cordic_SH1_srl_35_26_g1146 ( .a(cordic_SH1_srl_35_26_n_91), .b(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_106) );
fflopd cordic_Y_reg_7_ ( .CK(newNet_188), .D(cordic_n_77), .Q(cordic_Y_7_) );
NAND2_Z01 g15258 ( .a(n_295), .b(n_296), .o(n_402) );
fflopd PO_SERR_L_reg ( .CK(newNet_430), .D(n_432), .Q(PO_SERR_L) );
NAND2_Z01 cordic_AddX_MUX_1_g295 ( .a(cordic_AddX_Y_1), .b(cordic_X_8_), .o(cordic_AddX_MUX_1_n_26) );
XOR2_X1 g13413 ( .a(n_866), .b(PO_AD_17), .o(n_867) );
AND2_X1 g335 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_59) );
NAND2_Z01 cordic_AddY_MUX_1_g276 ( .a(cordic_AddY_MUX_1_n_14), .b(cordic_AddY_MUX_1_n_29), .o(cordic_AddY_Btemp_2_) );
XOR2_X1 cordic_AddX_Add_g689 ( .a(cordic_AddX_Add_n_43), .b(cordic_AddX_Add_n_26), .o(cordic_AddX_Stemp_4_) );
BUF_X2 newInst_241 ( .a(newNet_114), .o(newNet_241) );
NAND2_Z01 cordic_Add0_MUX_1_g261 ( .a(cordic_Add0_MUX_1_n_6), .b(cordic_Add0_MUX_1_n_25), .o(cordic_Add0_Btemp_10_) );
NAND2_Z01 g13563 ( .a(n_712), .b(CoreOutputReg_12_), .o(n_724) );
BUF_X2 newInst_901 ( .a(newNet_900), .o(newNet_901) );
XNOR2_X1 cordic_AddX_Compl_g375 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_4_), .o(cordic_AddX_Compl_n_7) );
NAND2_Z01 cordic_AddY_Add_g660 ( .a(cordic_AddY_Add_n_73), .b(cordic_AddY_Add_n_22), .o(cordic_AddY_Add_n_74) );
NAND2_Z01 g15090 ( .a(n_4), .b(PI_AD_8), .o(n_518) );
NAND2_Z01 g14942 ( .a(n_579), .b(n_503), .o(n_632) );
NOR2_Z1 cordic_g467 ( .a(cordic_n_12), .b(Issue_Rst), .o(cordic_n_40) );
NOR2_Z1 g15520 ( .a(n_100), .b(RESET), .o(n_143) );
XOR2_X1 cordic_Add0_Add_g655 ( .a(cordic_Add0_Add_n_50), .b(cordic_Add0_Add_n_29), .o(cordic_Add0_Stemp_7_) );
NAND2_Z01 g15556 ( .a(n_31), .b(State_1_), .o(n_116) );
BUF_X2 newInst_1123 ( .a(newNet_1122), .o(newNet_1123) );
BUF_X2 newInst_688 ( .a(newNet_164), .o(newNet_688) );
XOR2_X1 cordic_Add0_Add_g634 ( .a(cordic_Add0_Add_n_71), .b(cordic_Add0_Add_n_22), .o(cordic_Add0_Stemp_14_) );
INV_Z1 cordic_Add0_g51 ( .a(cordic_Add0_Btemp_10_), .o(cordic_Add0_n_11) );
BUF_X2 newInst_23 ( .a(newNet_22), .o(newNet_23) );
NAND2_Z01 g15289 ( .a(n_232), .b(n_120), .o(n_366) );
NAND2_Z01 cordic_Add0_Add_g666 ( .a(cordic_Add0_Add_n_39), .b(cordic_Add0_Add_n_6), .o(cordic_Add0_Add_n_41) );
INV_X2 newInst_281 ( .a(newNet_280), .o(newNet_281) );
fflopd CoreInput_reg_10_ ( .CK(newNet_822), .D(n_655), .Q(CoreInput_10_) );
NAND2_Z01 g13562 ( .a(n_712), .b(CoreOutputReg_25_), .o(n_725) );
NAND3_Z1 g15303 ( .a(n_211), .b(n_199), .c(n_152), .o(n_352) );
AND2_X1 g44 ( .a(n_844), .b(n_856), .o(PO_AD_20) );
AND2_X1 g354 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_40) );
NAND2_Z01 g13554 ( .a(n_712), .b(CoreOutputReg_29_), .o(n_733) );
BUF_X2 newInst_415 ( .a(newNet_414), .o(newNet_415) );
XOR2_X1 cordic_AddX_Compl_g342 ( .a(cordic_AddX_Compl_n_37), .b(cordic_AddX_Compl_n_12), .o(CoreOutput_29_) );
BUF_X2 newInst_1043 ( .a(newNet_1042), .o(newNet_1043) );
AND2_X1 cordic_pla_g292 ( .a(cordic_pla_n_9), .b(cordic_iteration_1_), .o(cordic_pla_n_18) );
XOR2_X1 cordic_Add0_Add_g640 ( .a(cordic_Add0_Add_n_65), .b(cordic_Add0_Add_n_19), .o(cordic_Add0_Stemp_12_) );
BUF_X2 newInst_1170 ( .a(newNet_1169), .o(newNet_1170) );
AND2_X1 cordic_AddX_Compl_g345 ( .a(cordic_AddX_Compl_n_35), .b(cordic_AddX_Compl_n_3), .o(cordic_AddX_Compl_n_37) );
INV_X1 cordic_SH1_srl_35_26_g1151 ( .a(cordic_SH1_srl_35_26_n_101), .o(cordic_SH1_srl_35_26_n_100) );
INV_X1 g15615 ( .a(n_46), .o(n_45) );
AND2_X1 g356 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_38) );
NAND2_Z01 cordic_AddX_MUX_0_g296 ( .a(cordic_BS1_0_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_25) );
NAND2_Z01 cordic_SH1_srl_35_26_g1124 ( .a(cordic_SH1_srl_35_26_n_124), .b(cordic_SH1_srl_35_26_n_106), .o(cordic_SH1_srl_35_26_n_128) );
BUF_X2 newInst_71 ( .a(newNet_70), .o(newNet_71) );
BUF_X2 newInst_1124 ( .a(newNet_1123), .o(newNet_1124) );
BUF_X2 newInst_1113 ( .a(newNet_1112), .o(newNet_1113) );
NAND2_Z01 cordic_AddY_g65 ( .a(cordic_AngleCin), .b(cordic_Ysign), .o(cordic_AddY_n_2) );
BUF_X2 newInst_1034 ( .a(newNet_1033), .o(newNet_1034) );
BUF_X2 newInst_454 ( .a(newNet_453), .o(newNet_454) );
BUF_X2 newInst_1063 ( .a(newNet_1062), .o(newNet_1063) );
AND2_X1 cordic_AddY_Compl_g355 ( .a(cordic_AddY_Compl_n_25), .b(cordic_AddY_Compl_n_4), .o(cordic_AddY_Compl_n_27) );
INV_Z1 g8017 ( .a(CoreOutputReg_33_), .o(n_900) );
BUF_X2 newInst_1031 ( .a(newNet_1030), .o(newNet_1031) );
BUF_X2 newInst_473 ( .a(newNet_472), .o(newNet_473) );
BUF_X2 newInst_355 ( .a(newNet_354), .o(newNet_355) );
XOR2_X1 cordic_Add0_Add_g649 ( .a(cordic_Add0_Add_n_56), .b(cordic_Add0_Add_n_21), .o(cordic_Add0_Stemp_9_) );
NAND2_Z01 g14959 ( .a(n_572), .b(Config_Reg_25_), .o(n_618) );
BUF_X2 newInst_792 ( .a(newNet_791), .o(newNet_792) );
NOR2_Z1 cordic_Add0_MUX_1_g274 ( .a(cordic_Add0_MUX_1_n_2), .b(cordic_Add0_MUX_1_n_1), .o(cordic_Add0_Btemp_14_) );
NAND2_Z01 cordic_Add0_Add_g653 ( .a(cordic_Add0_Add_n_53), .b(cordic_Add0_Add_n_17), .o(cordic_Add0_Add_n_54) );
XOR2_X1 g15593 ( .a(PI_AD_57), .b(PI_AD_40), .o(n_72) );
BUF_X2 newInst_248 ( .a(newNet_247), .o(newNet_248) );
NAND2_Z01 cordic_AddX_MUX_1_g274 ( .a(cordic_AddX_MUX_1_n_11), .b(cordic_AddX_MUX_1_n_28), .o(cordic_AddX_Btemp_12_) );
BUF_X2 newInst_153 ( .a(newNet_152), .o(newNet_153) );
BUF_X2 newInst_395 ( .a(newNet_394), .o(newNet_395) );
BUF_X2 newInst_453 ( .a(newNet_452), .o(newNet_453) );
INV_X1 cordic_g495 ( .a(CoreOutput_1_), .o(cordic_n_12) );
AND2_X1 g15148 ( .a(n_444), .b(n_218), .o(n_464) );
BUF_X2 newInst_62 ( .a(newNet_46), .o(newNet_62) );
NAND2_Z01 cordic_SH1_srl_35_26_g1245 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_14_), .o(cordic_SH1_srl_35_26_n_4) );
NAND2_Z01 cordic_Add0_MUX_1_g264 ( .a(cordic_Add0_MUX_1_n_3), .b(cordic_Add0_MUX_1_n_20), .o(cordic_Add0_Btemp_9_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1176 ( .a(cordic_SH1_srl_35_26_n_43), .b(cordic_SH1_srl_35_26_n_52), .o(cordic_SH1_srl_35_26_n_76) );
NAND2_Z01 cordic_SH2_srl_35_26_g1235 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_5_), .o(cordic_SH2_srl_35_26_n_14) );
XOR2_X1 cordic_AddY_Add_g656 ( .a(cordic_AddY_Add_n_76), .b(cordic_AddY_Add_n_25), .o(cordic_AddY_Stemp_15_) );
BUF_X2 newInst_617 ( .a(newNet_616), .o(newNet_617) );
XNOR2_X1 g13423 ( .a(PO_AD_0), .b(CBE_par_1_), .o(n_858) );
BUF_X2 newInst_908 ( .a(newNet_907), .o(newNet_908) );
INV_X1 g15648 ( .a(OutputAvail), .o(n_17) );
NAND2_Z01 cordic_g409 ( .a(Issue_Rst), .b(CoreInput_1_), .o(cordic_n_97) );
BUF_X2 newInst_874 ( .a(newNet_873), .o(newNet_874) );
BUF_X2 newInst_1 ( .a(newNet_0), .o(newNet_1) );
BUF_X2 newInst_596 ( .a(newNet_595), .o(newNet_596) );
NOR2_Z1 cordic_g457 ( .a(cordic_n_21), .b(Issue_Rst), .o(cordic_n_50) );
NAND2_Z01 cordic_AddX_Add_g727 ( .a(cordic_AddX_Btemp1_4_), .b(cordic_AddX_Atemp_4_), .o(cordic_AddX_Add_n_7) );
NAND2_Z01 cordic_SH2_srl_35_26_g1147 ( .a(cordic_SH2_srl_35_26_n_99), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_105) );
BUF_X2 newInst_443 ( .a(newNet_442), .o(newNet_443) );
BUF_X2 newInst_314 ( .a(newNet_31), .o(newNet_314) );
NAND2_Z01 g15395 ( .a(n_214), .b(CoreOutputReg_30_), .o(n_255) );
BUF_X2 newInst_543 ( .a(newNet_542), .o(newNet_543) );
NAND2_Z01 cordic_SH2_srl_35_26_g1161 ( .a(cordic_SH2_srl_35_26_n_79), .b(cordic_SH2_srl_35_26_n_61), .o(cordic_SH2_srl_35_26_n_91) );
INV_X1 g15528 ( .a(n_127), .o(n_126) );
AND2_X1 cordic_Add0_Compl_g351 ( .a(cordic_Add0_Compl_n_29), .b(cordic_Add0_Compl_n_10), .o(cordic_Add0_Compl_n_31) );
NAND2_Z01 cordic_AddX_Add_g722 ( .a(cordic_AddX_Btemp1_13_), .b(cordic_AddX_Atemp_13_), .o(cordic_AddX_Add_n_12) );
NAND2_Z01 g14965 ( .a(n_572), .b(Config_Reg_30_), .o(n_612) );
XOR2_X1 cordic_AddX_Add_g671 ( .a(cordic_AddX_Add_n_61), .b(cordic_AddX_Add_n_27), .o(cordic_AddX_Stemp_10_) );
AND2_X1 cordic_g474 ( .a(CoreOutput_29_), .b(Issue_Rst), .o(cordic_n_33) );
BUF_X2 newInst_331 ( .a(newNet_330), .o(newNet_331) );
INV_X1 cordic_pla_g308 ( .a(cordic_iteration_1_), .o(cordic_pla_n_3) );
INV_X1 cordic_SH2_srl_35_26_g1123 ( .a(cordic_SH2_srl_35_26_n_128), .o(cordic_SH2_srl_35_26_n_129) );
XOR2_X1 cordic_AddX_Add_g701 ( .a(cordic_AddX_Add_n_16), .b(cordic_AddX_Y_2), .o(cordic_AddX_Stemp_0_) );
INV_X1 g15654 ( .a(PI_REQ64_L), .o(n_11) );
BUF_X2 newInst_629 ( .a(newNet_628), .o(newNet_629) );
BUF_X2 newInst_1070 ( .a(newNet_1069), .o(newNet_1070) );
BUF_X2 newInst_881 ( .a(newNet_880), .o(newNet_881) );
NAND2_Z01 g15210 ( .a(n_380), .b(PI_PAR), .o(n_442) );
BUF_X2 newInst_573 ( .a(newNet_275), .o(newNet_573) );
BUF_X2 newInst_1143 ( .a(newNet_1142), .o(newNet_1143) );
BUF_X2 newInst_828 ( .a(newNet_827), .o(newNet_828) );
NAND3_Z1 g14804 ( .a(n_474), .b(n_706), .c(n_227), .o(n_709) );
XOR2_X1 cordic_AddY_Add_g680 ( .a(cordic_AddY_Add_n_52), .b(cordic_AddY_Add_n_30), .o(cordic_AddY_Stemp_7_) );
NAND2_Z01 cordic_AddX_MUX_0_g306 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_9_), .o(cordic_AddX_MUX_0_n_15) );
BUF_X2 newInst_183 ( .a(newNet_182), .o(newNet_183) );
NOR2_Z1 g15638 ( .a(State_0_), .b(State_2_), .o(n_31) );
NAND2_Z01 cordic_Add0_Add_g700 ( .a(cordic_Add0_n_11), .b(cordic_Add0_Atemp_10_), .o(cordic_Add0_Add_n_7) );
fflopd Core_Cnt_reg_3_ ( .CK(newNet_531), .D(n_224), .Q(Core_Cnt_3_) );
BUF_X2 newInst_965 ( .a(newNet_964), .o(newNet_965) );
NAND2_Z01 g15356 ( .a(n_214), .b(CoreOutputReg_16_), .o(n_305) );
BUF_X2 newInst_383 ( .a(newNet_382), .o(newNet_383) );
BUF_X2 newInst_1134 ( .a(newNet_902), .o(newNet_1134) );
BUF_X2 newInst_148 ( .a(newNet_147), .o(newNet_148) );
fflopd CoreInput_reg_5_ ( .CK(newNet_756), .D(n_644), .Q(CoreInput_5_) );
BUF_X2 newInst_398 ( .a(newNet_358), .o(newNet_398) );
AND3_X1 g15542 ( .a(n_39), .b(n_48), .c(Trdy_Wait_Cnt_2_), .o(n_120) );
BUF_X2 newInst_953 ( .a(newNet_445), .o(newNet_953) );
NAND2_Z01 cordic_AddY_MUX_0_g316 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_6_), .o(cordic_AddY_MUX_0_n_5) );
NAND2_Z01 cordic_g419 ( .a(Issue_Rst), .b(CoreInput_4_), .o(cordic_n_88) );
BUF_X2 newInst_940 ( .a(newNet_939), .o(newNet_940) );
NAND2_Z01 g15256 ( .a(n_299), .b(n_300), .o(n_404) );
INV_X1 cordic_Add0_Add_g707 ( .a(cordic_Add0_n_1), .o(cordic_Add0_Add_n_0) );
AND2_X1 g15469 ( .a(n_137), .b(PI_FRAME_L), .o(n_209) );
BUF_X2 newInst_1195 ( .a(newNet_1194), .o(newNet_1195) );
BUF_X2 newInst_362 ( .a(newNet_361), .o(newNet_362) );
BUF_X2 newInst_133 ( .a(newNet_132), .o(newNet_133) );
BUF_X2 newInst_269 ( .a(newNet_215), .o(newNet_269) );
BUF_X2 newInst_308 ( .a(newNet_307), .o(newNet_308) );
fflopd cordic_Y_reg_6_ ( .CK(newNet_51), .D(cordic_n_36), .Q(cordic_Y_6_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1189 ( .a(cordic_SH1_srl_35_26_n_45), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_63) );
NAND2_Z01 cordic_Add0_MUX_1_g289 ( .a(cordic_tanangle_0_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_12) );
NAND2_Z01 cordic_AddX_MUX_0_g275 ( .a(cordic_AddX_MUX_0_n_30), .b(cordic_AddX_MUX_0_n_15), .o(cordic_AddX_Atemp_9_) );
NAND2_Z01 g15400 ( .a(CoreOutput_33_), .b(n_2), .o(n_250) );
BUF_X2 newInst_464 ( .a(newNet_463), .o(newNet_464) );
NAND2_Z01 g13487 ( .a(n_730), .b(n_768), .o(n_797) );
fflopd CBE_par_reg_3_ ( .CK(newNet_1071), .D(n_349), .Q(CBE_par_3_) );
NAND2_Z01 cordic_AddX_MUX_0_g307 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_2_), .o(cordic_AddX_MUX_0_n_14) );
NAND2_Z01 g15058 ( .a(n_473), .b(PI_AD_22), .o(n_550) );
NAND2_Z01 g13549 ( .a(n_712), .b(CoreOutputReg_4_), .o(n_737) );
NAND2_Z01 cordic_AddX_MUX_0_g289 ( .a(cordic_BS1_15_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_32) );
NOR2_Z1 cordic_SH2_srl_35_26_g1129 ( .a(cordic_SH2_srl_35_26_n_100), .b(cordic_SH2_srl_35_26_n_19), .o(cordic_BS2_13_) );
BUF_X2 newInst_1185 ( .a(newNet_1184), .o(newNet_1185) );
NAND2_Z01 cordic_SH2_srl_35_26_g1202 ( .a(cordic_SH2_srl_35_26_n_9), .b(cordic_SH2_srl_35_26_n_34), .o(cordic_SH2_srl_35_26_n_49) );
INV_Z1 cordic_AddX_MUX_1_g321 ( .a(cordic_AddX_Y_1), .o(cordic_AddX_MUX_1_n_0) );
AND2_X1 g341 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_53) );
BUF_X2 newInst_190 ( .a(newNet_189), .o(newNet_190) );
BUF_X2 newInst_94 ( .a(newNet_93), .o(newNet_94) );
NAND2_Z01 cordic_AddX_Add_g669 ( .a(cordic_AddX_Add_n_64), .b(cordic_AddX_Add_n_29), .o(cordic_AddX_Add_n_65) );
NAND2_Z01 cordic_SH1_srl_35_26_g1181 ( .a(cordic_SH1_srl_35_26_n_57), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_71) );
NAND2_Z01 cordic_AddY_Add_g658 ( .a(cordic_AddY_Add_n_74), .b(cordic_AddY_Add_n_10), .o(cordic_AddY_Add_n_76) );
AND2_X1 cordic_SH1_srl_35_26_g1192 ( .a(cordic_SH1_srl_35_26_n_41), .b(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_60) );
BUF_X2 newInst_35 ( .a(newNet_34), .o(newNet_35) );
NAND2_Z01 g13382 ( .a(n_896), .b(TAR_TRI_P), .o(PO_PAR) );
NAND2_Z01 g15331 ( .a(n_184), .b(PI_AD_26), .o(n_330) );
XNOR2_X1 cordic_AddY_Compl_g374 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_13_), .o(cordic_AddY_Compl_n_8) );
AND3_X1 g14842 ( .a(Access_Address_1_31_), .b(n_628), .c(Access_Address_1_30_), .o(n_681) );
AND2_X1 g15530 ( .a(n_99), .b(Core_Cnt_0_), .o(n_140) );
NAND2_Z01 g14824 ( .a(n_692), .b(PO_DEVSEL_L), .o(n_696) );
NAND2_Z01 cordic_g435 ( .a(cordic_SumAngle_12_), .b(cordic_n_7), .o(cordic_n_72) );
XOR2_X1 g13403 ( .a(n_876), .b(PO_AD_18), .o(n_877) );
NAND2_Z01 cordic_SH1_srl_35_26_g1201 ( .a(cordic_SH1_srl_35_26_n_16), .b(cordic_SH1_srl_35_26_n_28), .o(cordic_SH1_srl_35_26_n_51) );
NOR2_Z1 g13462 ( .a(n_785), .b(n_710), .o(n_820) );
XNOR2_X1 cordic_AddX_Compl_g367 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_9_), .o(cordic_AddX_Compl_n_15) );
INV_Z1 cordic_Add0_g58 ( .a(cordic_Add0_Btemp_3_), .o(cordic_Add0_n_4) );
NAND2_Z01 g15412 ( .a(n_3), .b(PI_AD_29), .o(n_238) );
NAND2_Z01 cordic_AddY_MUX_0_g279 ( .a(cordic_AddY_MUX_0_n_25), .b(cordic_AddY_MUX_0_n_12), .o(cordic_AddY_Atemp_0_) );
BUF_X2 newInst_1024 ( .a(newNet_1023), .o(newNet_1024) );
NAND2_Z01 g15095 ( .a(n_473), .b(PI_AD_10), .o(n_513) );
XOR2_X1 g13389 ( .a(n_890), .b(PO_AD_14), .o(n_891) );
fflopd TAR_TRI_D_reg ( .CK(newNet_363), .D(n_699), .Q(TAR_TRI_D) );
BUF_X2 newInst_862 ( .a(newNet_861), .o(newNet_862) );
NAND2_Z01 cordic_AddY_MUX_1_g286 ( .a(cordic_AddY_MUX_1_n_4), .b(cordic_AddY_MUX_1_n_21), .o(cordic_AddY_Btemp_5_) );
NAND2_Z01 g13517 ( .a(Idsel), .b(Config_Reg_2_), .o(n_769) );
fflopd CoreOutputReg_reg_20_ ( .CK(newNet_665), .D(n_401), .Q(CoreOutputReg_20_) );
BUF_X2 newInst_1085 ( .a(newNet_1084), .o(newNet_1085) );
NAND3_Z1 cordic_SH2_srl_35_26_g1116 ( .a(cordic_SH2_srl_35_26_n_114), .b(cordic_SH2_srl_35_26_n_103), .c(cordic_SH2_srl_35_26_n_112), .o(cordic_BS2_6_) );
AND2_X1 g15633 ( .a(n_973), .b(n_19), .o(n_35) );
BUF_X2 newInst_621 ( .a(newNet_620), .o(newNet_621) );
NAND2_Z01 cordic_AddY_Add_g702 ( .a(cordic_AddY_Add_n_16), .b(cordic_AddY_Y_2), .o(cordic_AddY_Add_n_32) );
NAND2_Z01 cordic_AddX_MUX_1_g286 ( .a(cordic_AddX_MUX_1_n_4), .b(cordic_AddX_MUX_1_n_21), .o(cordic_AddX_Btemp_5_) );
NAND2_Z01 cordic_g442 ( .a(cordic_SumAngle_4_), .b(cordic_n_7), .o(cordic_n_65) );
BUF_X2 newInst_564 ( .a(newNet_563), .o(newNet_564) );
BUF_X2 newInst_141 ( .a(newNet_140), .o(newNet_141) );
BUF_X2 newInst_92 ( .a(newNet_91), .o(newNet_92) );
BUF_X2 newInst_57 ( .a(newNet_56), .o(newNet_57) );
INV_Z1 cordic_Add0_g46 ( .a(cordic_Add0_Btemp_15_), .o(cordic_Add0_n_16) );
NAND2_Z01 g15290 ( .a(n_219), .b(n_155), .o(n_365) );
INV_X2 newInst_422 ( .a(newNet_421), .o(newNet_422) );
fflopd cordic_X_reg_3_ ( .CK(newNet_133), .D(cordic_n_52), .Q(cordic_X_3_) );
NAND2_Z01 cordic_AddX_MUX_1_g293 ( .a(cordic_AddX_Y_1), .b(cordic_X_12_), .o(cordic_AddX_MUX_1_n_28) );
NAND2_Z01 cordic_Add0_Add_g697 ( .a(cordic_Add0_n_16), .b(cordic_Add0_Atemp_15_), .o(cordic_Add0_Add_n_10) );
AND2_X1 g14814 ( .a(n_701), .b(n_157), .o(n_705) );
NAND2_Z01 cordic_AddY_Add_g725 ( .a(cordic_AddY_Btemp1_0_), .b(cordic_AddY_Atemp_0_), .o(cordic_AddY_Add_n_9) );
BUF_X1 mybuffer0 ( .a(cordic_AngleCout), .o(PO_PAR64) );
NAND2_Z01 g15123 ( .a(n_445), .b(n_280), .o(n_486) );
BUF_X2 newInst_799 ( .a(newNet_798), .o(newNet_799) );
NAND2_Z01 cordic_AddY_Add_g722 ( .a(cordic_AddY_Btemp1_13_), .b(cordic_AddY_Atemp_13_), .o(cordic_AddY_Add_n_12) );
NAND2_Z01 cordic_AddX_MUX_1_g310 ( .a(cordic_BS1_12_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_11) );
INV_Z1 cordic_AddY_MUX_0_g321 ( .a(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_0) );
BUF_X2 newInst_304 ( .a(newNet_303), .o(newNet_304) );
NAND2_Z01 cordic_AddY_MUX_1_g280 ( .a(cordic_AddY_MUX_1_n_6), .b(cordic_AddY_MUX_1_n_23), .o(cordic_AddY_Btemp_11_) );
NAND2_Z01 cordic_Add0_Add_g633 ( .a(cordic_Add0_Add_n_72), .b(cordic_Add0_Add_n_9), .o(cordic_Add0_Add_n_74) );
NAND2_Z01 cordic_SH2_srl_35_26_g1179 ( .a(cordic_SH2_srl_35_26_n_42), .b(cordic_SH2_srl_35_26_n_39), .o(cordic_SH2_srl_35_26_n_73) );
BUF_X2 newInst_123 ( .a(newNet_122), .o(newNet_123) );
BUF_X2 newInst_99 ( .a(newNet_98), .o(newNet_99) );
BUF_X2 newInst_898 ( .a(newNet_897), .o(newNet_898) );
BUF_X2 newInst_534 ( .a(newNet_533), .o(newNet_534) );
fflopd cordic_Angle_reg_3_ ( .CK(newNet_237), .D(cordic_n_108), .Q(cordic_Angle_3_) );
fflopd cordic_Y_reg_10_ ( .CK(newNet_99), .D(cordic_n_38), .Q(cordic_Y_10_) );
INV_X1 g15505 ( .a(n_157), .o(n_156) );
NAND2_Z01 g14838 ( .a(n_681), .b(n_124), .o(n_685) );
BUF_X2 newInst_227 ( .a(newNet_226), .o(newNet_227) );
INV_Z1 cordic_Add0_g61 ( .a(cordic_Add0_Btemp_0_), .o(cordic_Add0_n_1) );
NAND2_Z01 cordic_SH2_srl_35_26_g1232 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_2_), .o(cordic_SH2_srl_35_26_n_17) );
AND2_X1 cordic_pla_g307 ( .a(cordic_iteration_1_), .b(cordic_iteration_0_), .o(cordic_pla_n_4) );
NAND2_Z01 cordic_SH2_srl_35_26_g1200 ( .a(cordic_SH2_srl_35_26_n_6), .b(cordic_SH2_srl_35_26_n_30), .o(cordic_SH2_srl_35_26_n_52) );
BUF_X2 newInst_977 ( .a(newNet_976), .o(newNet_977) );
fflopd CoreOutputReg_reg_0_ ( .CK(newNet_728), .D(n_414), .Q(CoreOutputReg_0_) );
BUF_X2 newInst_160 ( .a(newNet_159), .o(newNet_160) );
INV_X1 g15627 ( .a(n_31), .o(n_32) );
NAND3_Z1 g14829 ( .a(n_118), .b(n_687), .c(Check_Add_Parity), .o(n_691) );
AND2_X1 g56 ( .a(n_825), .b(n_856), .o(PO_AD_8) );
NAND3_Z1 cordic_SH1_srl_35_26_g1163 ( .a(cordic_SH1_srl_35_26_n_3), .b(cordic_SH1_srl_35_26_n_46), .c(cordic_iteration_2_), .o(cordic_SH1_srl_35_26_n_88) );
XNOR2_X1 cordic_Add0_Compl_g376 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_7_), .o(cordic_Add0_Compl_n_6) );
BUF_X2 newInst_1194 ( .a(newNet_1193), .o(newNet_1194) );
BUF_X2 newInst_740 ( .a(newNet_739), .o(newNet_740) );
BUF_X2 newInst_578 ( .a(newNet_577), .o(newNet_578) );
XOR2_X1 g15488 ( .a(n_81), .b(n_82), .o(n_175) );
NAND2_Z01 g14997 ( .a(n_572), .b(Config_Reg_15_), .o(n_580) );
BUF_X2 newInst_989 ( .a(newNet_988), .o(newNet_989) );
fflopd Config_Reg_reg_22_ ( .CK(newNet_963), .D(n_674), .Q(Config_Reg_22_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1110 ( .a(cordic_SH1_srl_35_26_n_131), .b(cordic_iteration_3_), .o(cordic_BS1_10_) );
NAND2_Z01 cordic_AddY_MUX_1_g315 ( .a(cordic_BS2_11_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_6) );
INV_X1 g13383 ( .a(PIO_PAR_Value_Hold), .o(n_896) );
AND2_X1 g33 ( .a(n_819), .b(n_856), .o(PO_AD_31) );
BUF_X2 newInst_1058 ( .a(newNet_644), .o(newNet_1058) );
BUF_X2 newInst_710 ( .a(newNet_683), .o(newNet_710) );
NAND2_Z01 cordic_Add0_MUX_1_g288 ( .a(cordic_tanangle_13_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_13) );
NAND2_Z01 g14984 ( .a(n_571), .b(CoreInput_3_), .o(n_593) );
AND2_X1 g13572 ( .a(PAR64_Int), .b(RESET), .o(n_715) );
XOR2_X1 cordic_AddX_Add_g659 ( .a(cordic_AddX_Add_n_73), .b(cordic_AddX_Add_n_22), .o(cordic_AddX_Stemp_14_) );
NOR2_Z1 g15631 ( .a(n_18), .b(Access_Type_1_2_), .o(n_36) );
NAND3_Z1 cordic_SH1_srl_35_26_g1117 ( .a(cordic_SH1_srl_35_26_n_110), .b(cordic_SH1_srl_35_26_n_111), .c(cordic_SH1_srl_35_26_n_109), .o(cordic_BS1_5_) );
XOR2_X1 cordic_AddX_Compl_g338 ( .a(cordic_AddX_Compl_n_41), .b(cordic_AddX_Compl_n_13), .o(CoreOutput_31_) );
NAND2_Z01 cordic_Add0_MUX_0_g289 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_0_), .o(cordic_Add0_MUX_0_n_14) );
NAND2_Z01 g15446 ( .a(n_144), .b(n_98), .o(n_208) );
BUF_X2 newInst_974 ( .a(newNet_973), .o(newNet_974) );
NAND2_Z01 cordic_Add0_MUX_0_g295 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_5_), .o(cordic_Add0_MUX_0_n_8) );
fflopd TAR_TRI_A_reg ( .CK(newNet_364), .D(n_573), .Q(TAR_TRI_A) );
BUF_X2 newInst_706 ( .a(newNet_705), .o(newNet_706) );
INV_X1 g15017 ( .a(n_564), .o(n_563) );
NAND2_Z01 cordic_AddY_MUX_0_g303 ( .a(cordic_BS2_4_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_18) );
XOR2_X1 g15607 ( .a(PI_AD_44), .b(PI_AD_38), .o(n_58) );
INV_X1 cordic_g483 ( .a(CoreOutput_19_), .o(cordic_n_24) );
BUF_X2 newInst_1102 ( .a(newNet_86), .o(newNet_1102) );
BUF_X2 newInst_723 ( .a(newNet_722), .o(newNet_723) );
BUF_X2 newInst_270 ( .a(newNet_269), .o(newNet_270) );
NAND2_Z01 g13484 ( .a(n_727), .b(n_766), .o(n_800) );
NAND2_Z01 g15293 ( .a(n_275), .b(Access_Type_1_0_), .o(n_362) );
NAND2_Z01 g13477 ( .a(n_733), .b(n_771), .o(n_807) );
NAND2_Z01 cordic_SH1_srl_35_26_g1168 ( .a(cordic_SH1_srl_35_26_n_51), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_84) );
BUF_X2 newInst_766 ( .a(newNet_765), .o(newNet_766) );
BUF_X2 newInst_550 ( .a(newNet_116), .o(newNet_550) );
NAND2_Z01 cordic_SH2_srl_35_26_g1174 ( .a(cordic_SH2_srl_35_26_n_43), .b(cordic_SH2_srl_35_26_n_45), .o(cordic_SH2_srl_35_26_n_78) );
INV_X2 cordic_SH2_srl_35_26_g1252 ( .a(cordic_iteration_0_), .o(cordic_SH2_srl_35_26_n_0) );
NAND2_Z01 cordic_Add0_MUX_0_g293 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_6_), .o(cordic_Add0_MUX_0_n_10) );
NAND2_Z01 cordic_AddX_MUX_0_g285 ( .a(cordic_AddX_MUX_0_n_19), .b(cordic_AddX_MUX_0_n_1), .o(cordic_AddX_Atemp_10_) );
BUF_X2 newInst_742 ( .a(newNet_741), .o(newNet_742) );
BUF_X2 newInst_196 ( .a(newNet_195), .o(newNet_196) );
NAND2_Z01 cordic_SH1_srl_35_26_g1228 ( .a(cordic_iteration_0_), .b(cordic_Y_15_), .o(cordic_SH1_srl_35_26_n_24) );
NAND3_Z1 cordic_SH1_srl_35_26_g1214 ( .a(cordic_SH1_srl_35_26_n_3), .b(cordic_SH1_srl_35_26_n_0), .c(cordic_Y_15_), .o(cordic_SH1_srl_35_26_n_41) );
NAND2_Z01 g15352 ( .a(n_214), .b(CoreOutputReg_14_), .o(n_309) );
BUF_X2 newInst_896 ( .a(newNet_895), .o(newNet_896) );
XOR2_X1 cordic_Add0_Add_g685 ( .a(cordic_Add0_n_15), .b(cordic_Add0_Atemp_14_), .o(cordic_Add0_Add_n_22) );
fflopd cordic_Y_reg_4_ ( .CK(newNet_57), .D(cordic_n_37), .Q(cordic_Y_4_) );
BUF_X2 newInst_1053 ( .a(newNet_1052), .o(newNet_1053) );
BUF_X2 newInst_501 ( .a(newNet_8), .o(newNet_501) );
NAND2_Z01 cordic_AddY_MUX_0_g285 ( .a(cordic_AddY_MUX_0_n_19), .b(cordic_AddY_MUX_0_n_1), .o(cordic_AddY_Atemp_10_) );
XOR2_X1 cordic_AddX_g202 ( .a(cordic_AddX_Btemp_7_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_7_) );
XOR2_X1 g15602 ( .a(PI_AD_23), .b(PI_AD_18), .o(n_63) );
XOR2_X1 g15315 ( .a(n_175), .b(n_176), .o(n_345) );
NOR3_Z1 g13505 ( .a(Idsel), .b(n_899), .c(PI_REQ64_L), .o(n_781) );
XOR2_X1 cordic_Add0_Add_g679 ( .a(cordic_Add0_n_14), .b(cordic_Add0_Atemp_13_), .o(cordic_Add0_Add_n_28) );
AND2_X1 g332 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_62) );
BUF_X2 newInst_758 ( .a(newNet_757), .o(newNet_758) );
NOR2_Z1 cordic_g428 ( .a(cordic_n_13), .b(Issue_Rst), .o(cordic_n_79) );
NAND2_Z01 cordic_SH1_srl_35_26_g1200 ( .a(cordic_SH1_srl_35_26_n_6), .b(cordic_SH1_srl_35_26_n_30), .o(cordic_SH1_srl_35_26_n_52) );
NAND2_Z01 cordic_AddX_MUX_0_g319 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_4_), .o(cordic_AddX_MUX_0_n_2) );
NAND2_Z01 g15364 ( .a(CoreOutput_19_), .b(n_2), .o(n_297) );
BUF_X2 newInst_421 ( .a(newNet_309), .o(newNet_421) );
NAND2_Z01 cordic_AddX_Add_g732 ( .a(cordic_AddX_Btemp1_1_), .b(cordic_AddX_Atemp_1_), .o(cordic_AddX_Add_n_2) );
NAND2_Z01 g15235 ( .a(n_274), .b(Access_Address_1_22_), .o(n_425) );
NAND2_Z01 g15067 ( .a(n_473), .b(PI_AD_2), .o(n_541) );
NAND2_Z01 g15511 ( .a(n_116), .b(CBE_par_1_), .o(n_150) );
NAND2_Z01 cordic_AddX_MUX_0_g320 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_10_), .o(cordic_AddX_MUX_0_n_1) );
XOR2_X1 cordic_Add0_Add_g687 ( .a(cordic_Add0_n_3), .b(cordic_Add0_Atemp_2_), .o(cordic_Add0_Add_n_20) );
NOR2_Z1 g13450 ( .a(n_794), .b(n_710), .o(n_832) );
fflopd CoreOutputReg_reg_21_ ( .CK(newNet_655), .D(n_400), .Q(CoreOutputReg_21_) );
NOR2_Z1 g13446 ( .a(n_795), .b(n_710), .o(n_836) );
NAND2_Z01 g15464 ( .a(n_128), .b(n_102), .o(n_213) );
XOR2_X1 g15316 ( .a(n_174), .b(n_170), .o(n_344) );
NAND2_Z01 g15239 ( .a(n_274), .b(Access_Address_1_25_), .o(n_421) );
BUF_X2 newInst_131 ( .a(newNet_130), .o(newNet_131) );
INV_Y1 cordic_SH1_srl_35_26_g1249 ( .a(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_3) );
NAND2_Z01 g15299 ( .a(n_272), .b(PI_CBE_L_3), .o(n_356) );
NAND2_Z01 cordic_Add0_MUX_1_g259 ( .a(cordic_Add0_MUX_1_n_12), .b(cordic_Add0_MUX_1_n_28), .o(cordic_Add0_Btemp_0_) );
fflopd Config_Reg_reg_11_ ( .CK(newNet_1046), .D(n_638), .Q(Config_Reg_11_) );
BUF_X2 newInst_755 ( .a(newNet_754), .o(newNet_755) );
BUF_X2 newInst_487 ( .a(newNet_486), .o(newNet_487) );
NAND3_Z1 g15304 ( .a(n_211), .b(n_198), .c(n_153), .o(n_351) );
fflopd CoreOutputReg_reg_19_ ( .CK(newNet_672), .D(n_403), .Q(CoreOutputReg_19_) );
NAND2_Z01 g13537 ( .a(Idsel), .b(Config_Reg_22_), .o(n_749) );
INV_X1 g14825 ( .a(n_694), .o(n_695) );
NAND2_Z01 cordic_AddY_MUX_0_g276 ( .a(cordic_AddY_MUX_0_n_29), .b(cordic_AddY_MUX_0_n_14), .o(cordic_AddY_Atemp_2_) );
NOR2_Z1 cordic_g468 ( .a(cordic_n_20), .b(Issue_Rst), .o(cordic_n_39) );
BUF_X2 newInst_1010 ( .a(newNet_1009), .o(newNet_1010) );
NAND3_Z1 g14820 ( .a(n_431), .b(n_692), .c(n_273), .o(n_699) );
fflopd Config_Reg_reg_14_ ( .CK(newNet_1019), .D(n_634), .Q(Config_Reg_14_) );
BUF_X2 newInst_384 ( .a(newNet_383), .o(newNet_384) );
NOR2_Z1 g13435 ( .a(n_813), .b(n_710), .o(n_847) );
NAND2_Z01 cordic_AddX_MUX_0_g279 ( .a(cordic_AddX_MUX_0_n_25), .b(cordic_AddX_MUX_0_n_12), .o(cordic_AddX_Atemp_0_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1170 ( .a(cordic_SH1_srl_35_26_n_48), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_82) );
BUF_X2 newInst_104 ( .a(newNet_103), .o(newNet_104) );
BUF_X2 newInst_177 ( .a(newNet_176), .o(newNet_177) );
fflopd cordic_Angle_reg_9_ ( .CK(newNet_212), .D(cordic_n_102), .Q(cordic_Angle_9_) );
fflopd CoreInput_reg_13_ ( .CK(newNet_797), .D(n_652), .Q(CoreInput_13_) );
fflopd Access_Address_1_reg_29_ ( .CK(newNet_1133), .D(n_472), .Q(Access_Address_1_29_) );
NAND2_Z01 g15390 ( .a(CoreOutput_28_), .b(n_2), .o(n_260) );
BUF_X2 newInst_1092 ( .a(newNet_47), .o(newNet_1092) );
BUF_X2 newInst_937 ( .a(newNet_507), .o(newNet_937) );
BUF_X2 newInst_565 ( .a(newNet_564), .o(newNet_565) );
fflopd PO_STOP_L_reg ( .CK(newNet_420), .D(n_568), .Q(PO_STOP_L) );
BUF_X2 newInst_934 ( .a(newNet_933), .o(newNet_934) );
BUF_X2 newInst_601 ( .a(newNet_600), .o(newNet_601) );
BUF_X2 newInst_981 ( .a(newNet_563), .o(newNet_981) );
NAND2_Z01 cordic_SH1_srl_35_26_g1140 ( .a(cordic_SH1_srl_35_26_n_93), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_112) );
BUF_X2 newInst_124 ( .a(newNet_123), .o(newNet_124) );
BUF_X2 newInst_719 ( .a(newNet_718), .o(newNet_719) );
NAND2_Z01 cordic_AddY_MUX_1_g297 ( .a(cordic_AddY_Y_1), .b(cordic_Y_7_), .o(cordic_AddY_MUX_1_n_24) );
NAND2_Z01 cordic_Add0_MUX_0_g273 ( .a(cordic_tanangle_1_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_30) );
NAND2_Z01 g15338 ( .a(n_184), .b(PI_AD_28), .o(n_323) );
BUF_X2 newInst_438 ( .a(newNet_437), .o(newNet_438) );
AND2_X1 cordic_Add0_Compl_g343 ( .a(cordic_Add0_Compl_n_37), .b(cordic_Add0_Compl_n_12), .o(cordic_Add0_Compl_n_39) );
NAND2_Z01 cordic_SH2_srl_35_26_g1107 ( .a(cordic_SH2_srl_35_26_n_130), .b(cordic_iteration_3_), .o(cordic_SH2_srl_35_26_n_145) );
XOR2_X1 cordic_Add0_Add_g680 ( .a(cordic_Add0_n_6), .b(cordic_Add0_Atemp_5_), .o(cordic_Add0_Add_n_27) );
BUF_X2 newInst_875 ( .a(newNet_571), .o(newNet_875) );
BUF_X2 newInst_110 ( .a(newNet_109), .o(newNet_110) );
NAND2_Z01 cordic_SH1_srl_35_26_g1177 ( .a(cordic_SH1_srl_35_26_n_51), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_75) );
BUF_X2 newInst_1064 ( .a(newNet_1063), .o(newNet_1064) );
BUF_X2 newInst_237 ( .a(newNet_236), .o(newNet_237) );
fflopd CoreInput_reg_15_ ( .CK(newNet_792), .D(n_649), .Q(CoreInput_15_) );
BUF_X2 newInst_685 ( .a(newNet_684), .o(newNet_685) );
BUF_X2 newInst_137 ( .a(newNet_136), .o(newNet_137) );
INV_X1 g15274 ( .a(n_382), .o(n_383) );
NOR2_Z6 cordic_AddY_g35 ( .a(cordic_AddY_n_5), .b(cordic_AngleCin), .o(cordic_AddY_Y_1) );
BUF_X2 newInst_956 ( .a(newNet_955), .o(newNet_956) );
BUF_X2 newInst_1204 ( .a(newNet_1203), .o(newNet_1204) );
BUF_X2 newInst_899 ( .a(newNet_898), .o(newNet_899) );
INV_X1 drc_bufs15659 ( .a(n_494), .o(n_7) );
NAND2_Z01 g14961 ( .a(n_572), .b(Config_Reg_27_), .o(n_616) );
BUF_X2 newInst_277 ( .a(newNet_276), .o(newNet_277) );
BUF_X2 newInst_86 ( .a(newNet_33), .o(newNet_86) );
XOR2_X1 cordic_Add0_Add_g670 ( .a(cordic_Add0_Add_n_35), .b(cordic_Add0_Add_n_20), .o(cordic_Add0_Stemp_2_) );
fflopd CoreOutputReg_reg_12_ ( .CK(newNet_709), .D(n_411), .Q(CoreOutputReg_12_) );
BUF_X2 newInst_117 ( .a(newNet_61), .o(newNet_117) );
NAND2_Z01 cordic_SH1_srl_35_26_g1141 ( .a(cordic_SH1_srl_35_26_n_101), .b(cordic_SH1_srl_35_26_n_20), .o(cordic_SH1_srl_35_26_n_111) );
NAND2_Z01 g15374 ( .a(n_214), .b(CoreOutputReg_23_), .o(n_287) );
NAND2_Z01 cordic_g421 ( .a(Issue_Rst), .b(CoreInput_6_), .o(cordic_n_86) );
BUF_X2 newInst_591 ( .a(newNet_590), .o(newNet_591) );
BUF_X2 newInst_866 ( .a(newNet_568), .o(newNet_866) );
XOR2_X1 cordic_Add0_Compl_g362 ( .a(cordic_Add0_Compl_n_17), .b(cordic_Add0_Compl_n_14), .o(cordic_SumAngle_2_) );
NAND2_Z01 g14998 ( .a(n_572), .b(Config_Reg_16_), .o(n_579) );
fflopd CoreOutputReg_reg_32_ ( .CK(newNet_597), .D(n_388), .Q(CoreOutputReg_32_) );
NAND2_Z01 g13559 ( .a(n_712), .b(CoreOutputReg_27_), .o(n_728) );
XOR2_X1 cordic_AddX_Compl_g356 ( .a(cordic_AddX_Compl_n_23), .b(cordic_AddX_Compl_n_5), .o(CoreOutput_22_) );
BUF_X2 newInst_1149 ( .a(newNet_1148), .o(newNet_1149) );
BUF_X2 newInst_739 ( .a(newNet_738), .o(newNet_739) );
BUF_X2 newInst_1039 ( .a(newNet_1038), .o(newNet_1039) );
NAND2_Z01 cordic_AddY_Add_g676 ( .a(cordic_AddY_Add_n_56), .b(cordic_AddY_Add_n_1), .o(cordic_AddY_Add_n_58) );
BUF_X2 newInst_555 ( .a(newNet_554), .o(newNet_555) );
BUF_X2 newInst_679 ( .a(newNet_678), .o(newNet_679) );
NOR2_Z1 cordic_g453 ( .a(cordic_n_23), .b(Issue_Rst), .o(cordic_n_54) );
BUF_X2 newInst_781 ( .a(newNet_780), .o(newNet_781) );
fflopd Config_Reg_reg_0_ ( .CK(newNet_1053), .D(n_639), .Q(Config_Reg_0_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1182 ( .a(cordic_SH1_srl_35_26_n_43), .b(cordic_SH1_srl_35_26_n_53), .o(cordic_SH1_srl_35_26_n_70) );
NAND2_Z01 g14981 ( .a(n_571), .b(CoreInput_16_), .o(n_596) );
BUF_X2 newInst_696 ( .a(newNet_695), .o(newNet_696) );
BUF_X2 newInst_344 ( .a(newNet_343), .o(newNet_344) );
NAND3_Z1 g15010 ( .a(n_514), .b(n_7), .c(n_10), .o(n_569) );
NOR2_Z1 cordic_g464 ( .a(cordic_n_8), .b(Issue_Rst), .o(cordic_n_43) );
XOR2_X1 g13404 ( .a(n_875), .b(PO_AD_21), .o(n_876) );
NAND2_Z01 cordic_Add0_Add_g645 ( .a(cordic_Add0_Add_n_60), .b(cordic_Add0_Add_n_7), .o(cordic_Add0_Add_n_62) );
fflopd Config_Reg_reg_31_ ( .CK(newNet_893), .D(n_662), .Q(Config_Reg_31_) );
BUF_X2 newInst_919 ( .a(newNet_918), .o(newNet_919) );
NAND2_Z01 cordic_AddX_MUX_1_g299 ( .a(cordic_AddX_Y_1), .b(cordic_X_6_), .o(cordic_AddX_MUX_1_n_22) );
NAND2_Z01 g15416 ( .a(n_3), .b(PI_AD_17), .o(n_234) );
NAND2_Z01 cordic_g394 ( .a(cordic_n_71), .b(cordic_n_93), .o(cordic_n_113) );
BUF_X2 newInst_1073 ( .a(newNet_1072), .o(newNet_1073) );
XOR2_X1 cordic_AddY_g202 ( .a(cordic_AddY_Btemp_7_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_7_) );
XOR2_X1 cordic_AddY_Compl_g360 ( .a(cordic_AddY_Compl_n_19), .b(cordic_AddY_Compl_n_16), .o(CoreOutput_3_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1159 ( .a(cordic_SH2_srl_35_26_n_83), .b(cordic_SH2_srl_35_26_n_65), .o(cordic_SH2_srl_35_26_n_93) );
NAND2_Z01 cordic_AddY_Add_g721 ( .a(cordic_AddY_Btemp1_10_), .b(cordic_AddY_Atemp_10_), .o(cordic_AddY_Add_n_13) );
NOR2_Z1 cordic_AddX_Compl_g381 ( .a(cordic_AddX_Compl_n_0), .b(cordic_AddX_Stemp_0_), .o(cordic_AddX_Compl_n_1) );
BUF_X2 newInst_597 ( .a(newNet_596), .o(newNet_597) );
NAND2_Z01 cordic_SH2_srl_35_26_g1198 ( .a(cordic_SH2_srl_35_26_n_13), .b(cordic_SH2_srl_35_26_n_26), .o(cordic_SH2_srl_35_26_n_54) );
NAND2_Z01 g14927 ( .a(n_594), .b(n_524), .o(n_647) );
BUF_X2 newInst_1035 ( .a(newNet_1034), .o(newNet_1035) );
BUF_X2 newInst_912 ( .a(newNet_911), .o(newNet_912) );
BUF_X2 newInst_84 ( .a(newNet_83), .o(newNet_84) );
BUF_X2 newInst_414 ( .a(newNet_413), .o(newNet_414) );
NAND2_Z01 g13523 ( .a(Idsel), .b(Config_Reg_12_), .o(n_763) );
NAND2_Z01 g13476 ( .a(n_738), .b(n_762), .o(n_808) );
fflopd Access_Address_1_reg_28_ ( .CK(newNet_1137), .D(n_475), .Q(Access_Address_1_28_) );
BUF_X2 newInst_651 ( .a(newNet_650), .o(newNet_651) );
XOR2_X1 cordic_AddY_g209 ( .a(cordic_AddY_Btemp_3_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_3_) );
NAND2_Z01 g15260 ( .a(n_291), .b(n_292), .o(n_400) );
BUF_X2 newInst_128 ( .a(newNet_62), .o(newNet_128) );
NAND2_Z01 cordic_SH1_srl_35_26_g1193 ( .a(cordic_SH1_srl_35_26_n_40), .b(cordic_SH1_srl_35_26_n_20), .o(cordic_SH1_srl_35_26_n_59) );
NAND2_Z01 cordic_AddX_MUX_0_g291 ( .a(cordic_BS1_9_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_30) );
NAND2_Z01 g15517 ( .a(n_95), .b(n_41), .o(n_145) );
INV_X2 newInst_610 ( .a(newNet_609), .o(newNet_610) );
NAND2_Z01 g15399 ( .a(n_214), .b(CoreOutputReg_33_), .o(n_251) );
BUF_X2 newInst_905 ( .a(newNet_330), .o(newNet_905) );
XOR2_X1 cordic_AddX_Add_g668 ( .a(cordic_AddX_Add_n_64), .b(cordic_AddX_Add_n_29), .o(cordic_AddX_Stemp_11_) );
NAND2_Z01 g13470 ( .a(n_742), .b(n_778), .o(n_814) );
BUF_X2 newInst_588 ( .a(newNet_587), .o(newNet_588) );
NAND2_Z01 cordic_AddX_Add_g672 ( .a(cordic_AddX_Add_n_61), .b(cordic_AddX_Add_n_27), .o(cordic_AddX_Add_n_62) );
BUF_X2 newInst_1142 ( .a(newNet_471), .o(newNet_1142) );
NAND2_Z01 cordic_AddX_MUX_1_g277 ( .a(cordic_AddX_MUX_1_n_10), .b(cordic_AddX_MUX_1_n_26), .o(cordic_AddX_Btemp_8_) );
NOR2_Z1 cordic_g461 ( .a(cordic_n_16), .b(Issue_Rst), .o(cordic_n_46) );
NAND2_Z01 g14977 ( .a(n_571), .b(CoreInput_12_), .o(n_600) );
BUF_X2 newInst_847 ( .a(newNet_846), .o(newNet_847) );
BUF_X2 newInst_1074 ( .a(newNet_1073), .o(newNet_1074) );
fflopd cordic_Xsign_reg ( .CK(newNet_116), .D(cordic_n_46), .Q(cordic_Xsign) );
NAND2_Z01 g15086 ( .a(n_4), .b(PI_AD_4), .o(n_522) );
INV_Y1 cordic_SH2_srl_35_26_g1249 ( .a(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_3) );
BUF_X2 newInst_638 ( .a(newNet_637), .o(newNet_638) );
NAND2_Z01 cordic_AddY_MUX_1_g309 ( .a(cordic_BS2_0_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_12) );
fflopd cordic_Ysign_reg ( .CK(newNet_198), .D(cordic_n_79), .Q(cordic_Ysign) );
BUF_X2 newInst_857 ( .a(newNet_751), .o(newNet_857) );
BUF_X2 newInst_0 ( .a(tau_clk), .o(newNet_0) );
fflopd CoreInput_reg_9_ ( .CK(newNet_734), .D(n_640), .Q(CoreInput_9_) );
XOR2_X1 g13397 ( .a(n_882), .b(PO_AD_16), .o(n_883) );
BUF_X2 newInst_852 ( .a(newNet_851), .o(newNet_852) );
AND2_X1 g350 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_44) );
BUF_X2 newInst_795 ( .a(newNet_366), .o(newNet_795) );
AND2_X1 cordic_AddY_Compl_g351 ( .a(cordic_AddY_Compl_n_29), .b(cordic_AddY_Compl_n_10), .o(cordic_AddY_Compl_n_31) );
fflopd CoreOutputReg_reg_2_ ( .CK(newNet_614), .D(n_391), .Q(CoreOutputReg_2_) );
NAND2_Z01 cordic_Add0_MUX_0_g288 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_13_), .o(cordic_Add0_MUX_0_n_15) );
BUF_X2 newInst_640 ( .a(newNet_639), .o(newNet_640) );
NAND2_Z01 g15015 ( .a(n_502), .b(PAR_Int), .o(n_567) );
XNOR2_X1 cordic_Add0_Compl_g367 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_9_), .o(cordic_Add0_Compl_n_15) );
NOR2_Z1 g15149 ( .a(n_445), .b(n_976), .o(n_463) );
XOR2_X1 cordic_Add0_Add_g658 ( .a(cordic_Add0_Add_n_47), .b(cordic_Add0_Add_n_30), .o(cordic_Add0_Stemp_6_) );
BUF_X2 newInst_615 ( .a(newNet_53), .o(newNet_615) );
NAND4_Z1 cordic_SH1_srl_35_26_g1105 ( .a(cordic_SH1_srl_35_26_n_68), .b(cordic_SH1_srl_35_26_n_117), .c(cordic_SH1_srl_35_26_n_144), .d(cordic_SH1_srl_35_26_n_73), .o(cordic_BS1_1_) );
BUF_X2 newInst_481 ( .a(newNet_480), .o(newNet_481) );
fflopd Access_Type_1_reg_2_ ( .CK(newNet_1101), .D(n_467), .Q(Access_Type_1_2_) );
BUF_X2 newInst_14 ( .a(newNet_13), .o(newNet_14) );
BUF_X2 newInst_265 ( .a(newNet_264), .o(newNet_265) );
AND2_X1 cordic_Add0_Compl_g357 ( .a(cordic_Add0_Compl_n_23), .b(cordic_Add0_Compl_n_5), .o(cordic_Add0_Compl_n_25) );
NAND2_Z01 cordic_AddY_Add_g664 ( .a(cordic_AddY_Add_n_68), .b(cordic_AddY_Add_n_4), .o(cordic_AddY_Add_n_70) );
XNOR2_X1 cordic_AddY_Compl_g369 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_14_), .o(cordic_AddY_Compl_n_13) );
XOR2_X1 g15611 ( .a(PI_AD_56), .b(PI_AD_49), .o(n_54) );
BUF_X2 newInst_215 ( .a(newNet_120), .o(newNet_215) );
NAND2_Z01 g15368 ( .a(CoreOutput_20_), .b(n_188), .o(n_293) );
XOR2_X1 cordic_AddY_Compl_g344 ( .a(cordic_AddY_Compl_n_35), .b(cordic_AddY_Compl_n_3), .o(CoreOutput_11_) );
BUF_X2 newInst_180 ( .a(newNet_179), .o(newNet_180) );
NAND2_Z01 cordic_SH1_srl_35_26_g1137 ( .a(cordic_SH1_srl_35_26_n_97), .b(cordic_SH1_srl_35_26_n_18), .o(cordic_SH1_srl_35_26_n_115) );
INV_X2 newInst_516 ( .a(newNet_515), .o(newNet_516) );
NAND2_Z01 g15251 ( .a(n_308), .b(n_309), .o(n_409) );
XOR2_X1 g15577 ( .a(PI_AD_26), .b(PI_AD_16), .o(n_88) );
NAND2_Z01 cordic_AddY_MUX_0_g296 ( .a(cordic_BS2_0_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_25) );
BUF_X2 newInst_460 ( .a(newNet_167), .o(newNet_460) );
BUF_X2 newInst_675 ( .a(newNet_674), .o(newNet_675) );
NAND2_Z01 cordic_SH2_srl_35_26_g1207 ( .a(cordic_SH2_srl_35_26_n_15), .b(cordic_SH2_srl_35_26_n_23), .o(cordic_SH2_srl_35_26_n_39) );
fflopd PO_TRDY_L_reg ( .CK(newNet_416), .D(n_478), .Q(PO_TRDY_L) );
BUF_X2 newInst_763 ( .a(newNet_762), .o(newNet_763) );
BUF_X2 newInst_380 ( .a(newNet_379), .o(newNet_380) );
BUF_X2 newInst_1005 ( .a(newNet_1004), .o(newNet_1005) );
BUF_X2 newInst_338 ( .a(newNet_337), .o(newNet_338) );
BUF_X2 newInst_746 ( .a(newNet_745), .o(newNet_746) );
BUF_X2 newInst_67 ( .a(newNet_66), .o(newNet_67) );
INV_X1 cordic_Add0_MUX_0_g302 ( .a(cordic_Angle_15_), .o(cordic_Add0_MUX_0_n_1) );
NAND2_Z01 cordic_pla_g304 ( .a(cordic_pla_n_2), .b(cordic_iteration_3_), .o(cordic_pla_n_8) );
NAND2_Z01 g14955 ( .a(n_572), .b(Config_Reg_21_), .o(n_622) );
XOR2_X1 cordic_AddX_Compl_g364 ( .a(cordic_AddX_Compl_n_11), .b(cordic_AddX_Compl_n_1), .o(CoreOutput_18_) );
NAND2_Z01 cordic_Add0_Add_g659 ( .a(cordic_Add0_Add_n_47), .b(cordic_Add0_Add_n_30), .o(cordic_Add0_Add_n_48) );
fflopd cordic_iteration_reg_0_ ( .CK(newNet_50), .D(cordic_n_35), .Q(cordic_iteration_0_) );
BUF_X2 newInst_77 ( .a(newNet_76), .o(newNet_77) );
BUF_X2 newInst_631 ( .a(newNet_630), .o(newNet_631) );
NAND2_Z01 cordic_g439 ( .a(cordic_SumAngle_1_), .b(cordic_n_7), .o(cordic_n_68) );
NAND2_Z01 cordic_SH1_srl_35_26_g1136 ( .a(cordic_SH1_srl_35_26_n_90), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_116) );
BUF_X2 newInst_824 ( .a(newNet_823), .o(newNet_824) );
fflopd CoreOutputReg_reg_6_ ( .CK(newNet_571), .D(n_376), .Q(CoreOutputReg_6_) );
fflopd CoreInput_reg_8_ ( .CK(newNet_737), .D(n_641), .Q(CoreInput_8_) );
BUF_X2 newInst_583 ( .a(newNet_582), .o(newNet_583) );
BUF_X2 newInst_419 ( .a(newNet_418), .o(newNet_419) );
XOR2_X1 cordic_Add0_Add_g661 ( .a(cordic_Add0_Add_n_44), .b(cordic_Add0_Add_n_27), .o(cordic_Add0_Stemp_5_) );
NAND2_Z01 cordic_pla_g275 ( .a(cordic_pla_n_23), .b(cordic_pla_n_2), .o(cordic_pla_n_36) );
AND2_X1 g359 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_35) );
BUF_X2 newInst_370 ( .a(newNet_369), .o(newNet_370) );
NAND2_Z01 cordic_SH2_srl_35_26_g1182 ( .a(cordic_SH2_srl_35_26_n_43), .b(cordic_SH2_srl_35_26_n_53), .o(cordic_SH2_srl_35_26_n_70) );
NAND3_Z1 g15144 ( .a(n_363), .b(n_357), .c(n_10), .o(n_467) );
NAND2_Z01 cordic_AddX_Add_g661 ( .a(cordic_AddX_Add_n_71), .b(cordic_AddX_Add_n_12), .o(cordic_AddX_Add_n_73) );
AND3_X1 g15571 ( .a(State_1_), .b(n_26), .c(State_2_), .o(n_106) );
NAND2_Z01 g13567 ( .a(n_712), .b(CoreOutputReg_6_), .o(n_720) );
BUF_X2 newInst_113 ( .a(newNet_112), .o(newNet_113) );
XOR2_X1 cordic_AddX_g207 ( .a(cordic_AddX_Btemp_10_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_10_) );
XOR2_X1 g15583 ( .a(PI_AD_30), .b(PI_AD_1), .o(n_82) );
NAND2_Z01 g14988 ( .a(n_571), .b(CoreInput_7_), .o(n_589) );
BUF_X2 newInst_1156 ( .a(newNet_1155), .o(newNet_1156) );
NAND2_Z01 g13468 ( .a(n_746), .b(n_779), .o(n_816) );
BUF_X2 newInst_1164 ( .a(newNet_1163), .o(newNet_1164) );
NAND2_Z01 cordic_AddX_Add_g685 ( .a(cordic_AddX_Add_n_47), .b(cordic_AddX_Add_n_11), .o(cordic_AddX_Add_n_49) );
BUF_X2 newInst_39 ( .a(newNet_38), .o(newNet_39) );
NAND2_Z01 cordic_AddY_MUX_0_g300 ( .a(cordic_BS2_5_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_21) );
AND2_X1 g15562 ( .a(n_32), .b(State_1_), .o(n_112) );
BUF_X2 newInst_548 ( .a(newNet_547), .o(newNet_548) );
BUF_X2 newInst_426 ( .a(newNet_425), .o(newNet_426) );
NAND2_Z01 cordic_AddY_MUX_1_g300 ( .a(cordic_AddY_Y_1), .b(cordic_Y_5_), .o(cordic_AddY_MUX_1_n_21) );
INV_X1 g15380 ( .a(n_280), .o(n_281) );
NAND2_Z01 g15536 ( .a(n_111), .b(n_10), .o(n_134) );
INV_X1 cordic_SH2_srl_35_26_g1152 ( .a(cordic_SH2_srl_35_26_n_95), .o(cordic_SH2_srl_35_26_n_94) );
BUF_X2 newInst_772 ( .a(newNet_771), .o(newNet_772) );
NAND2_Z01 cordic_SH1_srl_35_26_g1205 ( .a(cordic_SH1_srl_35_26_n_7), .b(cordic_SH1_srl_35_26_n_32), .o(cordic_SH1_srl_35_26_n_48) );
NAND2_Z01 cordic_AddX_Add_g675 ( .a(cordic_AddX_Add_n_58), .b(cordic_AddX_Add_n_21), .o(cordic_AddX_Add_n_59) );
NAND2_Z01 cordic_AddX_Add_g693 ( .a(cordic_AddX_Add_n_40), .b(cordic_AddX_Add_n_24), .o(cordic_AddX_Add_n_41) );
NAND2_Z01 g15403 ( .a(n_214), .b(CoreOutputReg_4_), .o(n_247) );
NAND2_Z01 g15334 ( .a(n_3), .b(PI_AD_27), .o(n_327) );
BUF_X2 newInst_205 ( .a(newNet_204), .o(newNet_205) );
NAND4_Z1 g14818 ( .a(n_46), .b(n_218), .c(n_687), .d(Check_Attr_Parity), .o(n_701) );
BUF_X2 newInst_560 ( .a(newNet_559), .o(newNet_560) );
NAND2_Z01 cordic_Add0_MUX_1_g292 ( .a(cordic_tanangle_3_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_9) );
INV_Z1 cordic_Add0_g49 ( .a(cordic_Add0_Btemp_12_), .o(cordic_Add0_n_13) );
BUF_X2 newInst_8 ( .a(newNet_7), .o(newNet_8) );
XOR2_X1 g13392 ( .a(n_887), .b(PO_AD_30), .o(n_888) );
AND2_X1 cordic_AddY_Compl_g349 ( .a(cordic_AddY_Compl_n_31), .b(cordic_AddY_Compl_n_15), .o(cordic_AddY_Compl_n_33) );
BUF_X2 newInst_151 ( .a(newNet_150), .o(newNet_151) );
BUF_X2 newInst_537 ( .a(newNet_536), .o(newNet_537) );
NAND2_Z01 g13566 ( .a(n_712), .b(CoreOutputReg_0_), .o(n_721) );
BUF_X2 newInst_163 ( .a(newNet_121), .o(newNet_163) );
NAND2_Z01 cordic_AddX_MUX_0_g278 ( .a(cordic_AddX_MUX_0_n_27), .b(cordic_AddX_MUX_0_n_13), .o(cordic_AddX_Atemp_1_) );
NAND2_Z01 cordic_AddY_MUX_0_g312 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_14_), .o(cordic_AddY_MUX_0_n_9) );
NAND2_Z01 cordic_AddY_Add_g728 ( .a(cordic_AddY_Btemp1_3_), .b(cordic_AddY_Atemp_3_), .o(cordic_AddY_Add_n_6) );
NAND2_Z01 g15413 ( .a(n_187), .b(Check_Data_Parity), .o(n_237) );
BUF_X2 newInst_810 ( .a(newNet_809), .o(newNet_810) );
BUF_X2 newInst_390 ( .a(newNet_389), .o(newNet_390) );
XOR2_X1 cordic_AddY_Add_g708 ( .a(cordic_AddY_Btemp1_4_), .b(cordic_AddY_Atemp_4_), .o(cordic_AddY_Add_n_26) );
NAND2_Z01 cordic_SH2_srl_35_26_g1124 ( .a(cordic_SH2_srl_35_26_n_124), .b(cordic_SH2_srl_35_26_n_106), .o(cordic_SH2_srl_35_26_n_128) );
BUF_X2 newInst_258 ( .a(newNet_257), .o(newNet_258) );
NAND2_Z01 cordic_SH1_srl_35_26_g1128 ( .a(cordic_SH1_srl_35_26_n_101), .b(cordic_iteration_2_), .o(cordic_SH1_srl_35_26_n_124) );
BUF_X2 newInst_448 ( .a(newNet_447), .o(newNet_448) );
NOR2_Z1 g15478 ( .a(n_119), .b(n_44), .o(n_181) );
BUF_X2 newInst_775 ( .a(newNet_128), .o(newNet_775) );
NAND2_Z01 cordic_SH1_srl_35_26_g1155 ( .a(cordic_SH1_srl_35_26_n_85), .b(cordic_SH1_srl_35_26_n_71), .o(cordic_SH1_srl_35_26_n_98) );
BUF_X2 newInst_406 ( .a(newNet_405), .o(newNet_406) );
BUF_X2 newInst_377 ( .a(newNet_316), .o(newNet_377) );
NOR4_Z1 g15479 ( .a(Access_Address_1_20_), .b(n_23), .c(n_27), .d(Access_Address_1_19_), .o(n_180) );
BUF_X2 newInst_75 ( .a(tau_clk), .o(newNet_75) );
fflopd Access_Type_1_reg_3_ ( .CK(newNet_1100), .D(n_466), .Q(Access_Type_1_3_) );
NAND2_Z01 cordic_AddX_MUX_1_g314 ( .a(cordic_BS1_15_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_7) );
NAND2_Z01 cordic_Add0_MUX_0_g262 ( .a(cordic_Add0_MUX_0_n_29), .b(cordic_Add0_MUX_0_n_12), .o(cordic_Add0_Atemp_7_) );
NOR2_Z1 cordic_Add0_MUX_1_g278 ( .a(cordic_Add0_MUX_1_n_2), .b(cordic_Add0_MUX_1_n_0), .o(cordic_Add0_Btemp_15_) );
NAND2_Z01 g15243 ( .a(n_336), .b(n_197), .o(n_417) );
BUF_X2 newInst_658 ( .a(newNet_657), .o(newNet_658) );
INV_X1 cordic_g501 ( .a(cordic_AddY_Stemp_0_), .o(cordic_n_6) );
BUF_X2 newInst_350 ( .a(newNet_349), .o(newNet_350) );
XOR2_X1 cordic_AddY_g198 ( .a(cordic_AddY_Btemp_14_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_14_) );
XOR2_X1 cordic_AddY_g205 ( .a(cordic_AddY_Btemp_5_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_5_) );
fflopd Config_Reg_reg_27_ ( .CK(newNet_919), .D(n_669), .Q(Config_Reg_27_) );
XOR2_X1 cordic_AddY_Add_g701 ( .a(cordic_AddY_Add_n_16), .b(cordic_AddY_Y_2), .o(cordic_AddY_Stemp_0_) );
BUF_X2 newInst_286 ( .a(newNet_285), .o(newNet_286) );
NAND2_Z01 cordic_SH2_srl_35_26_g1195 ( .a(cordic_SH2_srl_35_26_n_10), .b(cordic_SH2_srl_35_26_n_33), .o(cordic_SH2_srl_35_26_n_57) );
BUF_X2 newInst_161 ( .a(newNet_160), .o(newNet_161) );
NAND3_Z1 g15136 ( .a(n_323), .b(n_418), .c(n_10), .o(n_475) );
NAND2_Z01 g14934 ( .a(n_587), .b(n_517), .o(n_640) );
XNOR2_X1 cordic_Add0_Compl_g380 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_11_), .o(cordic_Add0_Compl_n_3) );
fflopd Config_Reg_reg_21_ ( .CK(newNet_972), .D(n_675), .Q(Config_Reg_21_) );
NAND2_Z01 g15620 ( .a(DevSel_Cnt_En), .b(n_10), .o(n_50) );
NAND2_Z01 g15057 ( .a(n_473), .b(PI_AD_21), .o(n_551) );
NAND2_Z01 g15350 ( .a(n_214), .b(CoreOutputReg_13_), .o(n_311) );
XOR2_X1 cordic_AddX_Add_g714 ( .a(cordic_AddX_Btemp1_2_), .b(cordic_AddX_Atemp_2_), .o(cordic_AddX_Add_n_20) );
XNOR2_X1 g13428 ( .a(Par64_Sgnl), .b(PAR64_Int_d), .o(n_854) );
BUF_X2 newInst_968 ( .a(newNet_967), .o(newNet_968) );
BUF_X2 newInst_602 ( .a(newNet_601), .o(newNet_602) );
XOR2_X1 cordic_AddY_Add_g689 ( .a(cordic_AddY_Add_n_43), .b(cordic_AddY_Add_n_26), .o(cordic_AddY_Stemp_4_) );
NAND2_Z01 cordic_AddY_MUX_1_g305 ( .a(cordic_BS2_3_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_16) );
NAND2_Z01 g15076 ( .a(n_4), .b(PI_AD_10), .o(n_532) );
BUF_X2 newInst_223 ( .a(newNet_222), .o(newNet_223) );
NAND2_Z01 g15508 ( .a(n_116), .b(CBE_par_2_), .o(n_153) );
NAND2_Z01 cordic_AddY_Add_g732 ( .a(cordic_AddY_Btemp1_1_), .b(cordic_AddY_Atemp_1_), .o(cordic_AddY_Add_n_2) );
NAND2_Z01 cordic_SH2_srl_35_26_g1165 ( .a(cordic_SH2_srl_35_26_n_54), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_87) );
BUF_X2 newInst_949 ( .a(newNet_948), .o(newNet_949) );
BUF_X2 newInst_95 ( .a(newNet_94), .o(newNet_95) );
BUF_X2 newInst_801 ( .a(newNet_800), .o(newNet_801) );
NAND2_Z01 g13507 ( .a(Idsel), .b(Config_Reg_3_), .o(n_779) );
XOR2_X1 cordic_AddY_g212 ( .a(cordic_AddY_Btemp_1_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_1_) );
BUF_X2 newInst_244 ( .a(newNet_243), .o(newNet_244) );
XOR2_X1 cordic_Add0_Compl_g348 ( .a(cordic_Add0_Compl_n_31), .b(cordic_Add0_Compl_n_15), .o(cordic_SumAngle_9_) );
NAND2_Z01 g15214 ( .a(n_346), .b(n_139), .o(n_438) );
NAND2_Z01 g13556 ( .a(n_712), .b(CoreOutputReg_13_), .o(n_731) );
NAND2_Z01 cordic_SH1_srl_35_26_g1132 ( .a(cordic_SH1_srl_35_26_n_96), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_120) );
NAND2_Z01 cordic_AddX_Add_g731 ( .a(cordic_AddX_Btemp1_2_), .b(cordic_AddX_Atemp_2_), .o(cordic_AddX_Add_n_3) );
NAND2_Z01 g15213 ( .a(n_385), .b(DevSel_Wait_Cnt_1_), .o(n_439) );
BUF_X2 newInst_1180 ( .a(newNet_1179), .o(newNet_1180) );
NAND2_Z01 cordic_Add0_MUX_1_g271 ( .a(cordic_AngleCin), .b(cordic_Angle_1_), .o(cordic_Add0_MUX_1_n_30) );
NAND2_Z01 cordic_AddX_MUX_1_g292 ( .a(cordic_AddX_Y_1), .b(cordic_X_2_), .o(cordic_AddX_MUX_1_n_29) );
NAND2_Z01 g15118 ( .a(n_446), .b(Par64_Sgnl), .o(n_491) );
XNOR2_X1 cordic_AddY_Compl_g378 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_15_), .o(cordic_AddY_Compl_n_2) );
XOR2_X1 g15503 ( .a(n_55), .b(n_56), .o(n_160) );
NAND2_Z01 g15465 ( .a(n_129), .b(Trdy_Wait_Cnt_0_), .o(n_194) );
BUF_X2 newInst_491 ( .a(newNet_490), .o(newNet_491) );
AND2_X1 g342 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_52) );
NAND2_Z01 g15408 ( .a(n_214), .b(CoreOutputReg_7_), .o(n_242) );
NAND2_Z01 g15359 ( .a(n_214), .b(CoreOutputReg_17_), .o(n_302) );
BUF_X2 newInst_829 ( .a(newNet_828), .o(newNet_829) );
INV_X2 newInst_469 ( .a(newNet_468), .o(newNet_469) );
NAND2_Z01 cordic_Add0_MUX_1_g268 ( .a(cordic_Add0_MUX_1_n_16), .b(cordic_Add0_MUX_1_n_17), .o(cordic_Add0_Btemp_2_) );
NAND2_Z01 g13430 ( .a(n_817), .b(Par_Sgnl), .o(n_852) );
BUF_X2 newInst_366 ( .a(newNet_365), .o(newNet_366) );
NOR2_Z1 cordic_SH1_srl_35_26_g1129 ( .a(cordic_SH1_srl_35_26_n_100), .b(cordic_SH1_srl_35_26_n_19), .o(cordic_BS1_13_) );
XOR2_X1 cordic_g353 ( .a(cordic_n_98), .b(cordic_iteration_2_), .o(cordic_n_119) );
NAND2_Z01 g15098 ( .a(n_473), .b(PI_AD_13), .o(n_510) );
NAND2_Z01 g14913 ( .a(n_608), .b(n_528), .o(n_661) );
NAND2_Z01 g15453 ( .a(n_132), .b(n_35), .o(n_217) );
BUF_X2 newInst_1130 ( .a(newNet_1129), .o(newNet_1130) );
BUF_X2 newInst_450 ( .a(newNet_449), .o(newNet_450) );
BUF_X2 newInst_815 ( .a(newNet_814), .o(newNet_815) );
XOR2_X1 cordic_Add0_Add_g637 ( .a(cordic_Add0_Add_n_68), .b(cordic_Add0_Add_n_28), .o(cordic_Add0_Stemp_13_) );
NAND2_Z01 cordic_g413 ( .a(Issue_Rst), .b(CoreInput_13_), .o(cordic_n_94) );
NAND2_Z01 cordic_Add0_MUX_1_g265 ( .a(cordic_Add0_MUX_1_n_5), .b(cordic_Add0_MUX_1_n_21), .o(cordic_Add0_Btemp_4_) );
NAND2_Z01 g14938 ( .a(n_583), .b(n_511), .o(n_636) );
AND2_X1 g48 ( .a(n_837), .b(n_856), .o(PO_AD_16) );
NAND2_Z01 cordic_SH2_srl_35_26_g1148 ( .a(cordic_SH2_srl_35_26_n_90), .b(cordic_SH2_srl_35_26_n_18), .o(cordic_SH2_srl_35_26_n_104) );
BUF_X2 newInst_1002 ( .a(newNet_1001), .o(newNet_1002) );
NAND2_Z01 cordic_AddX_MUX_0_g301 ( .a(cordic_BS1_13_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_20) );
NAND2_Z01 g13498 ( .a(n_719), .b(n_751), .o(n_786) );
BUF_X2 newInst_1178 ( .a(newNet_1177), .o(newNet_1178) );
NOR3_Z1 g15541 ( .a(n_24), .b(n_5), .c(DWord_Trans), .o(n_121) );
BUF_X2 newInst_467 ( .a(newNet_466), .o(newNet_467) );
NAND2_Z01 g13548 ( .a(n_712), .b(CoreOutputReg_17_), .o(n_738) );
BUF_X2 newInst_835 ( .a(newNet_834), .o(newNet_835) );
XOR2_X1 cordic_AddX_Add_g706 ( .a(cordic_AddX_Btemp1_6_), .b(cordic_AddX_Atemp_6_), .o(cordic_AddX_Add_n_28) );
BUF_X2 newInst_663 ( .a(newNet_662), .o(newNet_663) );
NAND3_Z1 g15000 ( .a(n_17), .b(n_564), .c(System_Busy), .o(n_577) );
NAND2_Z01 cordic_AddY_MUX_1_g275 ( .a(cordic_AddY_MUX_1_n_15), .b(cordic_AddY_MUX_1_n_30), .o(cordic_AddY_Btemp_9_) );
NAND2_Z01 g14970 ( .a(n_572), .b(Config_Reg_6_), .o(n_607) );
BUF_X2 newInst_147 ( .a(newNet_85), .o(newNet_147) );
INV_X1 cordic_g484 ( .a(CoreOutput_18_), .o(cordic_n_23) );
INV_X2 newInst_1127 ( .a(newNet_1126), .o(newNet_1127) );
XOR2_X1 g15496 ( .a(n_70), .b(n_69), .o(n_167) );
NAND3_Z1 g15128 ( .a(n_334), .b(n_427), .c(n_10), .o(n_482) );
NAND2_Z01 g13540 ( .a(n_712), .b(CoreOutputReg_3_), .o(n_746) );
BUF_X2 newInst_526 ( .a(newNet_525), .o(newNet_526) );
NAND2_Z01 cordic_Add0_Add_g638 ( .a(cordic_Add0_Add_n_68), .b(cordic_Add0_Add_n_28), .o(cordic_Add0_Add_n_69) );
AND2_X1 cordic_SH1_srl_35_26_g1149 ( .a(cordic_SH1_srl_35_26_n_89), .b(cordic_SH1_srl_35_26_n_1), .o(cordic_SH1_srl_35_26_n_103) );
INV_X1 cordic_g491 ( .a(CoreOutput_33_), .o(cordic_n_16) );
BUF_X2 newInst_1128 ( .a(newNet_1127), .o(newNet_1128) );
NAND2_Z01 cordic_SH2_srl_35_26_g1216 ( .a(cordic_iteration_0_), .b(cordic_X_13_), .o(cordic_SH2_srl_35_26_n_36) );
XOR2_X1 g15597 ( .a(PI_AD_43), .b(PI_AD_37), .o(n_68) );
NOR2_X6 g15455 ( .a(n_141), .b(RESET), .o(n_214) );
XOR2_X1 cordic_AddY_Add_g683 ( .a(cordic_AddY_Add_n_49), .b(cordic_AddY_Add_n_28), .o(cordic_AddY_Stemp_6_) );
INV_Z1 cordic_Add0_g54 ( .a(cordic_Add0_Btemp_7_), .o(cordic_Add0_n_8) );
NAND2_Z01 g14917 ( .a(n_604), .b(n_509), .o(n_657) );
BUF_X2 newInst_1021 ( .a(newNet_1020), .o(newNet_1021) );
BUF_X2 newInst_838 ( .a(newNet_837), .o(newNet_838) );
NAND2_Z01 g13530 ( .a(Idsel), .b(Config_Reg_9_), .o(n_756) );
NAND2_Z01 cordic_g400 ( .a(cordic_n_65), .b(cordic_n_87), .o(cordic_n_107) );
NAND2_Z01 cordic_SH2_srl_35_26_g1218 ( .a(cordic_iteration_0_), .b(cordic_X_1_), .o(cordic_SH2_srl_35_26_n_34) );
NAND2_Z01 cordic_AddY_MUX_0_g275 ( .a(cordic_AddY_MUX_0_n_30), .b(cordic_AddY_MUX_0_n_15), .o(cordic_AddY_Atemp_9_) );
INV_X1 cordic_AddX_Compl_g382 ( .a(cordic_AddX_Y_4), .o(cordic_AddX_Compl_n_0) );
fflopd Access_Address_1_reg_21_ ( .CK(newNet_1171), .D(n_484), .Q(Access_Address_1_21_) );
NAND2_Z01 g15551 ( .a(n_53), .b(Core_Cnt_2_), .o(n_105) );
BUF_X2 newInst_736 ( .a(newNet_735), .o(newNet_736) );
BUF_X2 newInst_608 ( .a(newNet_607), .o(newNet_608) );
NAND2_Z01 cordic_g446 ( .a(cordic_SumAngle_8_), .b(cordic_n_7), .o(cordic_n_61) );
NAND2_Z01 g14903 ( .a(n_618), .b(n_547), .o(n_671) );
NOR2_Z1 cordic_SH2_srl_35_26_g1112 ( .a(cordic_SH2_srl_35_26_n_129), .b(cordic_iteration_3_), .o(cordic_BS2_9_) );
BUF_X2 newInst_553 ( .a(newNet_552), .o(newNet_553) );
BUF_X2 newInst_220 ( .a(newNet_219), .o(newNet_220) );
NAND2_Z01 cordic_AddX_MUX_1_g306 ( .a(cordic_BS1_9_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_15) );
XNOR2_X1 cordic_AddY_Compl_g373 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_10_), .o(cordic_AddY_Compl_n_9) );
NAND2_Z01 g13512 ( .a(Idsel), .b(Config_Reg_19_), .o(n_774) );
BUF_X2 newInst_433 ( .a(newNet_432), .o(newNet_433) );
NAND2_Z01 g14993 ( .a(n_572), .b(Config_Reg_11_), .o(n_584) );
NAND2_Z01 g15068 ( .a(n_473), .b(PI_AD_30), .o(n_540) );
BUF_X2 newInst_964 ( .a(newNet_16), .o(newNet_964) );
NAND2_Z01 cordic_AddY_MUX_0_g289 ( .a(cordic_BS2_15_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_32) );
AND2_X1 g13502 ( .a(n_973), .b(Access_Type_1_0_), .o(n_799) );
NAND2_Z01 g15355 ( .a(CoreOutput_15_), .b(n_2), .o(n_306) );
XOR2_X1 g15002 ( .a(n_559), .b(n_164), .o(n_575) );
NAND2_Z01 g15297 ( .a(n_272), .b(PI_CBE_L_1), .o(n_358) );
BUF_X2 newInst_1111 ( .a(newNet_776), .o(newNet_1111) );
BUF_X2 newInst_616 ( .a(newNet_615), .o(newNet_616) );
INV_X2 cordic_g500 ( .a(Issue_Rst), .o(cordic_n_7) );
NAND2_Z01 g15220 ( .a(n_353), .b(n_209), .o(n_434) );
BUF_X2 newInst_945 ( .a(newNet_944), .o(newNet_945) );
NOR2_Z1 cordic_SH2_srl_35_26_g1247 ( .a(cordic_SH2_srl_35_26_n_1), .b(cordic_iteration_2_), .o(cordic_SH2_srl_35_26_n_20) );
NAND2_Z01 cordic_AddX_MUX_1_g318 ( .a(cordic_BS1_13_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_3) );
XOR2_X1 cordic_Add0_Add_g678 ( .a(cordic_Add0_n_8), .b(cordic_Add0_Atemp_7_), .o(cordic_Add0_Add_n_29) );
BUF_X2 newInst_924 ( .a(newNet_923), .o(newNet_924) );
BUF_X2 newInst_996 ( .a(newNet_540), .o(newNet_996) );
NOR2_Z1 cordic_pla_g284 ( .a(cordic_pla_n_5), .b(cordic_pla_n_13), .o(cordic_tanangle_10_) );
NAND2_Z01 g15052 ( .a(n_473), .b(PI_AD_17), .o(n_556) );
NAND2_Z01 g15448 ( .a(n_148), .b(n_10), .o(n_206) );
BUF_X2 newInst_359 ( .a(newNet_358), .o(newNet_359) );
BUF_X2 newInst_3 ( .a(newNet_2), .o(newNet_3) );
NAND2_Z01 cordic_SH2_srl_35_26_g1226 ( .a(cordic_iteration_0_), .b(cordic_X_11_), .o(cordic_SH2_srl_35_26_n_26) );
XOR2_X1 cordic_Add0_Compl_g337 ( .a(cordic_Add0_Compl_n_43), .b(cordic_Add0_Compl_n_2), .o(cordic_SumAngle_15_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1217 ( .a(cordic_iteration_0_), .b(cordic_Y_4_), .o(cordic_SH1_srl_35_26_n_35) );
NAND2_Z01 cordic_AddX_Add_g663 ( .a(cordic_AddX_Add_n_70), .b(cordic_AddX_Add_n_23), .o(cordic_AddX_Add_n_71) );
AND2_X1 g37 ( .a(n_832), .b(n_856), .o(PO_AD_27) );
NAND3_Z1 g15134 ( .a(n_330), .b(n_422), .c(n_10), .o(n_477) );
XOR2_X1 cordic_Add0_Add_g690 ( .a(cordic_Add0_n_9), .b(cordic_Add0_Atemp_8_), .o(cordic_Add0_Add_n_17) );
BUF_X2 newInst_991 ( .a(newNet_990), .o(newNet_991) );
BUF_X2 newInst_691 ( .a(newNet_690), .o(newNet_691) );
BUF_X2 newInst_403 ( .a(newNet_402), .o(newNet_403) );
NAND2_Z01 cordic_Add0_MUX_1_g285 ( .a(cordic_tanangle_2_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_16) );
INV_X1 cordic_g479 ( .a(CoreOutput_7_), .o(cordic_n_28) );
INV_X1 g15646 ( .a(Access_Type_1_0_), .o(n_19) );
BUF_X2 newInst_1112 ( .a(newNet_1111), .o(newNet_1112) );
NAND2_Z01 g13536 ( .a(Idsel), .b(Config_Reg_5_), .o(n_750) );
INV_Z1 cordic_g17 ( .a(cordic_AngleCin), .o(cordic_n_144) );
BUF_X2 newInst_1119 ( .a(newNet_1118), .o(newNet_1119) );
BUF_X2 newInst_204 ( .a(newNet_203), .o(newNet_204) );
BUF_X2 newInst_1018 ( .a(newNet_1017), .o(newNet_1018) );
BUF_X2 newInst_585 ( .a(newNet_584), .o(newNet_585) );
NAND2_Z01 cordic_SH1_srl_35_26_g1210 ( .a(cordic_SH1_srl_35_26_n_11), .b(cordic_SH1_srl_35_26_n_36), .o(cordic_SH1_srl_35_26_n_44) );
fflopd Config_Reg_reg_6_ ( .CK(newNet_865), .D(n_660), .Q(Config_Reg_6_) );
BUF_X2 newInst_374 ( .a(newNet_373), .o(newNet_374) );
AND2_X1 g32 ( .a(n_850), .b(n_856), .o(PO_AD_32) );
BUF_X2 newInst_1155 ( .a(newNet_1154), .o(newNet_1155) );
XNOR2_X1 cordic_AddX_Compl_g366 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_3_), .o(cordic_AddX_Compl_n_16) );
INV_Y1 cordic_Add0_MUX_0_g301 ( .a(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_2) );
NAND2_Z01 g13529 ( .a(Idsel), .b(Config_Reg_4_), .o(n_757) );
NAND4_Z1 g15020 ( .a(n_276), .b(n_367), .c(n_448), .d(n_117), .o(n_564) );
NAND2_Z01 g15271 ( .a(n_290), .b(n_253), .o(n_389) );
BUF_X2 newInst_788 ( .a(newNet_787), .o(newNet_788) );
BUF_X2 newInst_36 ( .a(newNet_35), .o(newNet_36) );
NAND2_Z01 cordic_AddX_MUX_1_g282 ( .a(cordic_AddX_MUX_1_n_5), .b(cordic_AddX_MUX_1_n_22), .o(cordic_AddX_Btemp_6_) );
BUF_X2 newInst_909 ( .a(newNet_908), .o(newNet_909) );
BUF_X2 newInst_856 ( .a(newNet_855), .o(newNet_856) );
XOR2_X1 cordic_AddX_Add_g718 ( .a(cordic_AddX_Btemp1_0_), .b(cordic_AddX_Atemp_0_), .o(cordic_AddX_Add_n_16) );
NAND2_Z01 g15063 ( .a(n_473), .b(PI_AD_26), .o(n_545) );
fflopd Burst_Trans_reg ( .CK(newNet_1095), .D(n_407), .Q(Burst_Trans) );
fflopd CoreOutputReg_reg_31_ ( .CK(newNet_598), .D(n_389), .Q(CoreOutputReg_31_) );
BUF_X2 newInst_574 ( .a(newNet_573), .o(newNet_574) );
BUF_X2 newInst_508 ( .a(newNet_436), .o(newNet_508) );
fflopd Config_Reg_reg_12_ ( .CK(newNet_1037), .D(n_636), .Q(Config_Reg_12_) );
NAND2_Z01 g15264 ( .a(n_282), .b(n_283), .o(n_396) );
AND2_X1 cordic_Add0_Compl_g359 ( .a(cordic_Add0_Compl_n_21), .b(cordic_Add0_Compl_n_7), .o(cordic_Add0_Compl_n_23) );
XOR2_X1 cordic_AddX_Add_g710 ( .a(cordic_AddX_Btemp1_3_), .b(cordic_AddX_Atemp_3_), .o(cordic_AddX_Add_n_24) );
BUF_X2 newInst_844 ( .a(newNet_843), .o(newNet_844) );
NAND2_Z01 g15632 ( .a(n_19), .b(Access_Type_1_2_), .o(n_29) );
BUF_X2 newInst_709 ( .a(newNet_708), .o(newNet_709) );
NAND2_Z01 g15628 ( .a(Trdy_Wait_Cnt_0_), .b(Trdy_Wait_Cnt_1_), .o(n_39) );
NOR2_Z1 cordic_g331 ( .a(cordic_n_121), .b(Issue_Rst), .o(cordic_n_123) );
NAND3_Z1 g15306 ( .a(n_211), .b(n_200), .c(n_151), .o(n_349) );
NOR2_Z1 g15560 ( .a(n_51), .b(RESET), .o(n_113) );
AND2_X1 cordic_AddY_Compl_g359 ( .a(cordic_AddY_Compl_n_21), .b(cordic_AddY_Compl_n_7), .o(cordic_AddY_Compl_n_23) );
NAND2_Z01 cordic_AddX_MUX_0_g312 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_14_), .o(cordic_AddX_MUX_0_n_9) );
NAND2_Z01 g14808 ( .a(n_703), .b(n_702), .o(n_708) );
BUF_X2 newInst_959 ( .a(newNet_958), .o(newNet_959) );
NAND2_Z01 g15121 ( .a(n_444), .b(n_132), .o(n_488) );
BUF_X2 newInst_1086 ( .a(newNet_1085), .o(newNet_1086) );
NAND2_Z01 cordic_AddY_MUX_0_g301 ( .a(cordic_BS2_13_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_20) );
NAND2_Z01 cordic_AddY_Add_g696 ( .a(cordic_AddY_Add_n_37), .b(cordic_AddY_Add_n_20), .o(cordic_AddY_Add_n_38) );
NAND2_Z01 cordic_AddX_MUX_0_g308 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_1_), .o(cordic_AddX_MUX_0_n_13) );
BUF_X2 newInst_65 ( .a(newNet_64), .o(newNet_65) );
XOR2_X1 g15603 ( .a(PI_AD_46), .b(PI_AD_45), .o(n_62) );
NOR2_Z1 g15481 ( .a(n_135), .b(n_157), .o(n_187) );
BUF_X2 newInst_345 ( .a(newNet_344), .o(newNet_345) );
NAND2_Z01 cordic_AddY_Add_g673 ( .a(cordic_AddY_Add_n_59), .b(cordic_AddY_Add_n_5), .o(cordic_AddY_Add_n_61) );
XOR2_X1 cordic_AddX_Add_g662 ( .a(cordic_AddX_Add_n_70), .b(cordic_AddX_Add_n_23), .o(cordic_AddX_Stemp_13_) );
fflopd CoreOutputReg_reg_7_ ( .CK(newNet_562), .D(n_375), .Q(CoreOutputReg_7_) );
NAND2_Z01 cordic_Add0_MUX_0_g278 ( .a(cordic_tanangle_5_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_25) );
NAND2_Z01 cordic_Add0_MUX_1_g256 ( .a(cordic_Add0_MUX_1_n_4), .b(cordic_Add0_MUX_1_n_22), .o(cordic_Add0_Btemp_12_) );
NAND2_Z01 g13543 ( .a(n_712), .b(CoreOutputReg_2_), .o(n_743) );
NAND2_Z01 g14989 ( .a(n_571), .b(CoreInput_8_), .o(n_588) );
BUF_X2 newInst_715 ( .a(newNet_714), .o(newNet_715) );
BUF_X2 newInst_226 ( .a(newNet_225), .o(newNet_226) );
AND2_X1 g47 ( .a(n_840), .b(n_856), .o(PO_AD_17) );
BUF_X2 newInst_1167 ( .a(newNet_1166), .o(newNet_1167) );
NAND2_Z01 cordic_SH1_srl_35_26_g1120 ( .a(cordic_SH1_srl_35_26_n_125), .b(cordic_SH1_srl_35_26_n_121), .o(cordic_SH1_srl_35_26_n_132) );
BUF_X2 newInst_504 ( .a(newNet_503), .o(newNet_504) );
NAND2_Z01 cordic_Add0_MUX_1_g298 ( .a(cordic_tanangle_9_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_3) );
NAND2_Z01 g15388 ( .a(CoreOutput_27_), .b(n_188), .o(n_262) );
BUF_X2 newInst_698 ( .a(newNet_697), .o(newNet_698) );
BUF_X2 newInst_232 ( .a(newNet_231), .o(newNet_232) );
BUF_X2 newInst_558 ( .a(newNet_557), .o(newNet_558) );
BUF_X2 newInst_1025 ( .a(newNet_1024), .o(newNet_1025) );
fflopd CoreOutputReg_reg_10_ ( .CK(newNet_723), .D(n_413), .Q(CoreOutputReg_10_) );
NAND2_Z01 cordic_AddX_MUX_0_g292 ( .a(cordic_BS1_2_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_29) );
BUF_X2 newInst_1196 ( .a(newNet_1195), .o(newNet_1196) );
XOR2_X1 cordic_Add0_Add_g673 ( .a(cordic_Add0_Add_n_32), .b(cordic_Add0_Add_n_18), .o(cordic_Add0_Stemp_1_) );
NAND2_Z01 g14940 ( .a(n_581), .b(n_508), .o(n_634) );
BUF_X2 newInst_830 ( .a(newNet_829), .o(newNet_830) );
AND2_X1 cordic_pla_g268 ( .a(cordic_tanangle_2_), .b(cordic_pla_n_28), .o(cordic_tanangle_1_) );
NAND2_Z01 g15211 ( .a(n_385), .b(DevSel_Wait_Cnt_2_), .o(n_441) );
BUF_X2 newInst_1101 ( .a(newNet_758), .o(newNet_1101) );
BUF_X2 newInst_913 ( .a(newNet_912), .o(newNet_913) );
NAND2_Z01 cordic_SH2_srl_35_26_g1224 ( .a(cordic_iteration_0_), .b(cordic_X_9_), .o(cordic_SH2_srl_35_26_n_28) );
NAND2_Z01 g15460 ( .a(n_138), .b(PI_CBE_L_2), .o(n_198) );
XOR2_X1 cordic_AddY_Add_g674 ( .a(cordic_AddY_Add_n_58), .b(cordic_AddY_Add_n_21), .o(cordic_AddY_Stemp_9_) );
BUF_X2 newInst_411 ( .a(newNet_410), .o(newNet_411) );
BUF_X2 newInst_29 ( .a(newNet_28), .o(newNet_29) );
XOR2_X1 cordic_AddY_Compl_g354 ( .a(cordic_AddY_Compl_n_25), .b(cordic_AddY_Compl_n_4), .o(CoreOutput_6_) );
NAND2_Z01 g15417 ( .a(n_3), .b(PI_AD_18), .o(n_233) );
AND2_X1 cordic_AddY_Compl_g363 ( .a(cordic_AddY_Compl_n_17), .b(cordic_AddY_Compl_n_14), .o(cordic_AddY_Compl_n_19) );
NAND2_Z01 cordic_AddX_MUX_0_g282 ( .a(cordic_AddX_MUX_0_n_22), .b(cordic_AddX_MUX_0_n_5), .o(cordic_AddX_Atemp_6_) );
XOR2_X1 g13400 ( .a(n_879), .b(PO_AD_12), .o(n_880) );
NAND2_Z01 g14902 ( .a(n_619), .b(n_548), .o(n_672) );
NAND3_Z1 g15125 ( .a(n_333), .b(n_426), .c(n_10), .o(n_484) );
NAND2_Z01 g15250 ( .a(n_310), .b(n_311), .o(n_410) );
BUF_X2 newInst_735 ( .a(newNet_175), .o(newNet_735) );
NAND2_Z01 cordic_AddY_MUX_1_g316 ( .a(cordic_BS2_6_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_5) );
BUF_X2 newInst_1160 ( .a(newNet_1159), .o(newNet_1160) );
fflopd CoreCnt_En_reg ( .CK(newNet_844), .D(n_326), .Q(CoreCnt_En) );
NAND2_Z01 g14956 ( .a(n_572), .b(Config_Reg_22_), .o(n_621) );
NAND2_Z01 g14994 ( .a(n_572), .b(Config_Reg_12_), .o(n_583) );
INV_X1 g15640 ( .a(DevSel_Wait_Cnt_1_), .o(n_25) );
BUF_X2 newInst_1169 ( .a(newNet_153), .o(newNet_1169) );
XOR2_X1 cordic_AddY_Add_g706 ( .a(cordic_AddY_Btemp1_6_), .b(cordic_AddY_Atemp_6_), .o(cordic_AddY_Add_n_28) );
NOR2_Z1 g13432 ( .a(n_781), .b(n_710), .o(n_850) );
XOR2_X1 g15160 ( .a(n_344), .b(n_345), .o(n_452) );
fflopd Config_Reg_reg_28_ ( .CK(newNet_916), .D(n_668), .Q(Config_Reg_28_) );
NAND2_Z01 g15301 ( .a(n_267), .b(n_50), .o(n_354) );
NAND2_Z01 g14969 ( .a(n_572), .b(Config_Reg_5_), .o(n_608) );
BUF_X2 newInst_1069 ( .a(newNet_1068), .o(newNet_1069) );
BUF_X2 newInst_387 ( .a(newNet_386), .o(newNet_387) );
XNOR2_X1 cordic_AddX_Compl_g376 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_7_), .o(cordic_AddX_Compl_n_6) );
NAND2_Z01 cordic_Add0_MUX_0_g257 ( .a(cordic_Add0_MUX_0_n_24), .b(cordic_Add0_MUX_0_n_15), .o(cordic_Add0_Atemp_13_) );
NAND2_Z01 g15152 ( .a(n_444), .b(n_278), .o(n_460) );
INV_X1 cordic_g493 ( .a(CoreOutput_6_), .o(cordic_n_14) );
XOR2_X1 cordic_AddY_g203 ( .a(cordic_AddY_Btemp_11_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_11_) );
BUF_X2 newInst_263 ( .a(newNet_94), .o(newNet_263) );
XOR2_X1 cordic_Add0_Compl_g364 ( .a(cordic_Add0_Compl_n_11), .b(cordic_Add0_Compl_n_1), .o(cordic_SumAngle_1_) );
NOR4_Z1 g15442 ( .a(DevSel_Cnt_En), .b(n_110), .c(n_157), .d(PI_FRAME_L), .o(n_266) );
INV_X1 g15111 ( .a(n_495), .o(n_496) );
BUF_X2 newInst_482 ( .a(newNet_481), .o(newNet_482) );
NAND2_Z01 cordic_SH1_srl_35_26_g1223 ( .a(cordic_iteration_0_), .b(cordic_Y_3_), .o(cordic_SH1_srl_35_26_n_29) );
INV_X1 cordic_SH1_srl_35_26_g1119 ( .a(cordic_SH1_srl_35_26_n_132), .o(cordic_SH1_srl_35_26_n_133) );
BUF_X2 newInst_630 ( .a(newNet_385), .o(newNet_630) );
BUF_X2 newInst_1106 ( .a(newNet_1105), .o(newNet_1106) );
NOR2_Z1 g13459 ( .a(n_787), .b(n_710), .o(n_823) );
NAND2_Z01 g13520 ( .a(Idsel), .b(Config_Reg_14_), .o(n_766) );
NAND2_Z01 cordic_g415 ( .a(Issue_Rst), .b(CoreInput_15_), .o(cordic_n_92) );
BUF_X2 newInst_1077 ( .a(newNet_1076), .o(newNet_1077) );
NAND2_Z01 cordic_SH1_srl_35_26_g1209 ( .a(cordic_SH1_srl_35_26_n_14), .b(cordic_SH1_srl_35_26_n_25), .o(cordic_SH1_srl_35_26_n_45) );
BUF_X2 newInst_1118 ( .a(newNet_1117), .o(newNet_1118) );
INV_X3 g13577 ( .a(TAR_TRI_A), .o(n_710) );
BUF_X2 newInst_727 ( .a(newNet_726), .o(newNet_727) );
BUF_X2 newInst_432 ( .a(newNet_431), .o(newNet_432) );
BUF_X2 newInst_157 ( .a(newNet_156), .o(newNet_157) );
NAND2_Z01 cordic_AddY_MUX_0_g280 ( .a(cordic_AddY_MUX_0_n_23), .b(cordic_AddY_MUX_0_n_6), .o(cordic_AddY_Atemp_11_) );
NAND2_Z01 cordic_AddX_MUX_1_g280 ( .a(cordic_AddX_MUX_1_n_6), .b(cordic_AddX_MUX_1_n_23), .o(cordic_AddX_Btemp_11_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1160 ( .a(cordic_SH2_srl_35_26_n_82), .b(cordic_SH2_srl_35_26_n_63), .o(cordic_SH2_srl_35_26_n_92) );
NAND2_Z01 cordic_AddY_Add_g693 ( .a(cordic_AddY_Add_n_40), .b(cordic_AddY_Add_n_24), .o(cordic_AddY_Add_n_41) );
BUF_X2 newInst_1016 ( .a(newNet_1015), .o(newNet_1016) );
BUF_X2 newInst_122 ( .a(newNet_121), .o(newNet_122) );
fflopd Idsel_reg ( .CK(newNet_467), .D(n_492), .Q(Idsel) );
NAND2_Z01 g15116 ( .a(n_441), .b(n_195), .o(n_493) );
NAND2_Z01 g15427 ( .a(n_215), .b(State_1_), .o(n_227) );
NAND2_Z01 g15266 ( .a(n_262), .b(n_263), .o(n_394) );
XOR2_X1 g15581 ( .a(PI_AD_31), .b(PI_AD_0), .o(n_84) );
XOR2_X1 g13417 ( .a(n_862), .b(PO_AD_3), .o(n_863) );
BUF_X2 newInst_753 ( .a(newNet_752), .o(newNet_753) );
BUF_X2 newInst_109 ( .a(newNet_108), .o(newNet_109) );
NAND3_X1 g2 ( .a(n_1062), .b(Set_Data_Parity), .c(n_10), .o(n_1063) );
NAND2_Z01 g14908 ( .a(n_613), .b(n_541), .o(n_666) );
BUF_X2 newInst_761 ( .a(newNet_760), .o(newNet_761) );
BUF_X2 newInst_336 ( .a(newNet_335), .o(newNet_336) );
BUF_X2 newInst_518 ( .a(newNet_284), .o(newNet_518) );
NAND2_Z01 cordic_Add0_Add_g635 ( .a(cordic_Add0_Add_n_71), .b(cordic_Add0_Add_n_22), .o(cordic_Add0_Add_n_72) );
NAND2_Z01 cordic_g436 ( .a(cordic_SumAngle_13_), .b(cordic_n_7), .o(cordic_n_71) );
BUF_X2 newInst_1097 ( .a(newNet_1096), .o(newNet_1097) );
INV_X1 cordic_pla_g298 ( .a(cordic_pla_n_12), .o(cordic_pla_n_13) );
BUF_X2 newInst_408 ( .a(newNet_407), .o(newNet_408) );
XOR2_X1 g13412 ( .a(n_867), .b(PO_AD_24), .o(n_868) );
AND2_X1 cordic_AddY_Compl_g347 ( .a(cordic_AddY_Compl_n_33), .b(cordic_AddY_Compl_n_9), .o(cordic_AddY_Compl_n_35) );
fflopd Access_Address_1_reg_24_ ( .CK(newNet_1153), .D(n_479), .Q(Access_Address_1_24_) );
NAND2_Z01 g14964 ( .a(n_572), .b(Config_Reg_2_), .o(n_613) );
BUF_X2 newInst_243 ( .a(newNet_242), .o(newNet_243) );
NAND2_Z01 cordic_SH2_srl_35_26_g1136 ( .a(cordic_SH2_srl_35_26_n_90), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_116) );
fflopd Trdy_Wait_Cnt_reg_0_ ( .CK(newNet_321), .D(n_228), .Q(Trdy_Wait_Cnt_0_) );
NAND2_Z01 g14919 ( .a(n_602), .b(n_532), .o(n_655) );
NAND2_Z01 g15073 ( .a(n_473), .b(PI_AD_6), .o(n_535) );
BUF_X2 newInst_902 ( .a(newNet_901), .o(newNet_902) );
BUF_X2 newInst_701 ( .a(newNet_700), .o(newNet_701) );
NAND2_Z01 cordic_SH2_srl_35_26_g1132 ( .a(cordic_SH2_srl_35_26_n_96), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_120) );
NAND3_Z1 g15569 ( .a(DevSel_Wait_Cnt_0_), .b(n_13), .c(DevSel_Wait_Cnt_1_), .o(n_95) );
NAND2_Z01 cordic_AddX_MUX_0_g283 ( .a(cordic_AddX_MUX_0_n_31), .b(cordic_AddX_MUX_0_n_9), .o(cordic_AddX_Atemp_14_) );
NAND2_Z01 g15327 ( .a(n_3), .b(PI_AD_20), .o(n_334) );
NOR2_Z1 cordic_g448 ( .a(cordic_n_18), .b(Issue_Rst), .o(cordic_n_59) );
NAND2_Z01 g13509 ( .a(Idsel), .b(Config_Reg_1_), .o(n_777) );
AND2_X1 g55 ( .a(n_827), .b(n_856), .o(PO_AD_9) );
NAND2_Z01 cordic_AddX_MUX_1_g273 ( .a(cordic_AddX_MUX_1_n_7), .b(cordic_AddX_MUX_1_n_32), .o(cordic_AddX_Btemp_15_) );
NAND2_Z01 g14933 ( .a(n_588), .b(n_518), .o(n_641) );
NAND2_Z01 g15324 ( .a(n_204), .b(n_40), .o(n_337) );
fflopd cordic_Y_reg_13_ ( .CK(newNet_85), .D(cordic_n_43), .Q(cordic_Y_13_) );
BUF_X2 newInst_485 ( .a(newNet_234), .o(newNet_485) );
NAND2_Z01 g15105 ( .a(n_473), .b(PI_AD_16), .o(n_503) );
BUF_X2 newInst_490 ( .a(newNet_489), .o(newNet_490) );
NAND2_Z01 cordic_Add0_Add_g706 ( .a(cordic_Add0_n_9), .b(cordic_Add0_Atemp_8_), .o(cordic_Add0_Add_n_1) );
BUF_X2 newInst_668 ( .a(newNet_667), .o(newNet_668) );
INV_X1 cordic_g487 ( .a(CoreOutput_2_), .o(cordic_n_20) );
BUF_X2 newInst_1203 ( .a(newNet_1202), .o(newNet_1203) );
NAND2_Z01 g15531 ( .a(n_5), .b(n_10), .o(n_139) );
BUF_X2 newInst_323 ( .a(newNet_322), .o(newNet_323) );
INV_Z1 cordic_Add0_g59 ( .a(cordic_Add0_Btemp_2_), .o(cordic_Add0_n_3) );
INV_X1 g15475 ( .a(n_183), .o(n_182) );
NAND2_Z01 cordic_SH2_srl_35_26_g1178 ( .a(cordic_SH2_srl_35_26_n_42), .b(cordic_SH2_srl_35_26_n_53), .o(cordic_SH2_srl_35_26_n_74) );
NAND2_Z01 cordic_SH2_srl_35_26_g1108 ( .a(cordic_SH2_srl_35_26_n_128), .b(cordic_iteration_3_), .o(cordic_SH2_srl_35_26_n_144) );
fflopd PIO_PAR_Value_Hold_reg ( .CK(newNet_1201), .D(n_1063), .Q(PIO_PAR_Value_Hold) );
XOR2_X1 cordic_AddX_g211 ( .a(cordic_AddX_Btemp_2_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_2_) );
AND2_X1 g52 ( .a(n_833), .b(n_856), .o(PO_AD_12) );
XOR2_X1 g15504 ( .a(n_54), .b(n_68), .o(n_159) );
NAND2_Z01 g15218 ( .a(n_347), .b(n_271), .o(n_435) );
BUF_X2 newInst_303 ( .a(newNet_290), .o(newNet_303) );
BUF_X2 newInst_397 ( .a(newNet_396), .o(newNet_397) );
BUF_X2 newInst_1140 ( .a(newNet_1139), .o(newNet_1140) );
NAND2_Z01 g14923 ( .a(n_598), .b(n_527), .o(n_651) );
fflopd Check_Attr_Parity_reg ( .CK(newNet_1065), .D(n_707), .Q(Check_Attr_Parity) );
NOR2_Z1 g13461 ( .a(n_815), .b(n_710), .o(n_821) );
NAND2_Z01 cordic_g402 ( .a(cordic_n_63), .b(cordic_n_85), .o(cordic_n_105) );
BUF_X2 newInst_891 ( .a(newNet_890), .o(newNet_891) );
BUF_X2 newInst_339 ( .a(newNet_338), .o(newNet_339) );
NAND2_Z01 cordic_SH1_srl_35_26_g1161 ( .a(cordic_SH1_srl_35_26_n_79), .b(cordic_SH1_srl_35_26_n_61), .o(cordic_SH1_srl_35_26_n_91) );
AND2_X1 cordic_AddX_Compl_g359 ( .a(cordic_AddX_Compl_n_21), .b(cordic_AddX_Compl_n_7), .o(cordic_AddX_Compl_n_23) );
BUF_X2 newInst_676 ( .a(newNet_675), .o(newNet_676) );
BUF_X2 newInst_307 ( .a(newNet_306), .o(newNet_307) );
NAND2_Z01 g15255 ( .a(n_301), .b(n_302), .o(n_405) );
NAND2_Z01 cordic_SH2_srl_35_26_g1128 ( .a(cordic_SH2_srl_35_26_n_101), .b(cordic_iteration_2_), .o(cordic_SH2_srl_35_26_n_124) );
fflopd cordic_Y_reg_5_ ( .CK(newNet_55), .D(cordic_n_57), .Q(cordic_Y_5_) );
fflopd cordic_iteration_reg_2_ ( .CK(newNet_293), .D(cordic_n_122), .Q(cordic_iteration_2_) );
XOR2_X1 cordic_AddY_Add_g713 ( .a(cordic_AddY_Btemp1_9_), .b(cordic_AddY_Atemp_9_), .o(cordic_AddY_Add_n_21) );
NAND2_Z01 cordic_SH1_srl_35_26_g1180 ( .a(cordic_SH1_srl_35_26_n_42), .b(cordic_SH1_srl_35_26_n_49), .o(cordic_SH1_srl_35_26_n_72) );
NAND2_Z01 cordic_SH1_srl_35_26_g1109 ( .a(cordic_SH1_srl_35_26_n_132), .b(cordic_iteration_3_), .o(cordic_SH1_srl_35_26_n_143) );
XOR2_X1 g15590 ( .a(PI_AD_28), .b(PI_AD_7), .o(n_75) );
BUF_X2 newInst_363 ( .a(newNet_222), .o(newNet_363) );
NAND2_Z01 g13518 ( .a(Idsel), .b(Config_Reg_28_), .o(n_768) );
BUF_X2 newInst_254 ( .a(newNet_253), .o(newNet_254) );
BUF_X2 newInst_1001 ( .a(newNet_1000), .o(newNet_1001) );
NAND2_Z01 cordic_Add0_MUX_0_g291 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_7_), .o(cordic_Add0_MUX_0_n_12) );
NAND2_Z01 cordic_pla_g300 ( .a(cordic_pla_n_1), .b(cordic_iteration_0_), .o(cordic_pla_n_11) );
NAND2_Z01 cordic_AddY_MUX_0_g305 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_3_), .o(cordic_AddY_MUX_0_n_16) );
NAND2_Z01 cordic_AddX_Add_g657 ( .a(cordic_AddX_Add_n_76), .b(cordic_AddX_Add_n_25), .o(cordic_AddX_Add_n_77) );
BUF_X2 newInst_950 ( .a(newNet_949), .o(newNet_950) );
NAND2_Z01 g15246 ( .a(n_319), .b(n_320), .o(n_414) );
NAND2_Z01 g15432 ( .a(n_186), .b(n_192), .o(n_225) );
BUF_X2 newInst_800 ( .a(newNet_799), .o(newNet_800) );
INV_X2 cordic_Add0_g45 ( .a(cordic_Add0_Y_3), .o(cordic_AngleCout) );
NAND2_Z01 g15240 ( .a(n_274), .b(Access_Address_1_27_), .o(n_420) );
BUF_X2 newInst_861 ( .a(newNet_860), .o(newNet_861) );
NAND2_Z01 cordic_AddX_MUX_1_g289 ( .a(cordic_AddX_Y_1), .b(cordic_X_15_), .o(cordic_AddX_MUX_1_n_32) );
NAND2_Z01 g15410 ( .a(n_214), .b(CoreOutputReg_8_), .o(n_240) );
BUF_X2 newInst_803 ( .a(newNet_802), .o(newNet_803) );
BUF_X2 newInst_354 ( .a(newNet_353), .o(newNet_354) );
NAND2_Z01 cordic_Add0_Add_g698 ( .a(cordic_Add0_n_15), .b(cordic_Add0_Atemp_14_), .o(cordic_Add0_Add_n_9) );
BUF_X2 newInst_533 ( .a(newNet_532), .o(newNet_533) );
NAND2_Z01 cordic_AddX_MUX_1_g294 ( .a(cordic_AddX_Y_1), .b(cordic_X_1_), .o(cordic_AddX_MUX_1_n_27) );
NAND2_Z01 g15347 ( .a(n_214), .b(CoreOutputReg_12_), .o(n_314) );
XOR2_X1 cordic_Add0_Compl_g344 ( .a(cordic_Add0_Compl_n_35), .b(cordic_Add0_Compl_n_3), .o(cordic_SumAngle_11_) );
NAND2_Z01 g15450 ( .a(n_135), .b(PO_SERR_L), .o(n_218) );
NAND2_Z01 cordic_g425 ( .a(Issue_Rst), .b(CoreInput_0_), .o(cordic_n_82) );
BUF_X2 newInst_620 ( .a(newNet_552), .o(newNet_620) );
BUF_X2 newInst_946 ( .a(newNet_945), .o(newNet_946) );
fflopd PAR_Int_d_reg ( .CK(newNet_1204), .D(n_716), .Q(PAR_Int_d) );
BUF_X2 newInst_1175 ( .a(newNet_1174), .o(newNet_1175) );
NAND2_Z01 cordic_SH2_srl_35_26_g1156 ( .a(cordic_SH2_srl_35_26_n_86), .b(cordic_SH2_srl_35_26_n_69), .o(cordic_SH2_srl_35_26_n_97) );
fflopd cordic_Angle_reg_4_ ( .CK(newNet_234), .D(cordic_n_107), .Q(cordic_Angle_4_) );
NAND3_Z1 g15140 ( .a(n_322), .b(n_415), .c(n_10), .o(n_471) );
NOR2_Z1 g15009 ( .a(n_564), .b(n_463), .o(n_570) );
BUF_X2 newInst_1047 ( .a(newNet_29), .o(newNet_1047) );
INV_X2 newInst_140 ( .a(newNet_139), .o(newNet_140) );
XNOR2_X1 cordic_AddY_Compl_g377 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_5_), .o(cordic_AddY_Compl_n_5) );
BUF_X2 newInst_89 ( .a(newNet_88), .o(newNet_89) );
XNOR2_X1 cordic_Add0_Compl_g378 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_15_), .o(cordic_Add0_Compl_n_2) );
INV_X1 cordic_g507 ( .a(CoreOutput_14_), .o(cordic_n_0) );
NAND2_Z01 cordic_AddY_MUX_1_g281 ( .a(cordic_AddY_MUX_1_n_8), .b(cordic_AddY_MUX_1_n_24), .o(cordic_AddY_Btemp_7_) );
NAND2_Z01 cordic_AddY_MUX_0_g278 ( .a(cordic_AddY_MUX_0_n_27), .b(cordic_AddY_MUX_0_n_13), .o(cordic_AddY_Atemp_1_) );
NAND2_Z01 g15282 ( .a(n_235), .b(n_325), .o(n_373) );
NAND2_Z01 g15124 ( .a(n_445), .b(n_157), .o(n_485) );
BUF_X2 newInst_840 ( .a(newNet_839), .o(newNet_840) );
NAND2_Z01 cordic_SH2_srl_35_26_g1186 ( .a(cordic_SH2_srl_35_26_n_47), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_66) );
BUF_X2 newInst_386 ( .a(newNet_385), .o(newNet_386) );
NAND2_Z01 cordic_SH2_srl_35_26_g1205 ( .a(cordic_SH2_srl_35_26_n_7), .b(cordic_SH2_srl_35_26_n_32), .o(cordic_SH2_srl_35_26_n_48) );
BUF_X2 newInst_525 ( .a(newNet_524), .o(newNet_525) );
NAND3_Z1 g15313 ( .a(n_185), .b(n_183), .c(n_49), .o(n_346) );
BUF_X2 newInst_266 ( .a(newNet_265), .o(newNet_266) );
NAND2_Z01 g14905 ( .a(n_616), .b(n_544), .o(n_669) );
NAND2_Z01 cordic_AddY_MUX_1_g287 ( .a(cordic_AddY_MUX_1_n_2), .b(cordic_AddY_MUX_1_n_18), .o(cordic_AddY_Btemp_4_) );
BUF_X2 newInst_515 ( .a(newNet_514), .o(newNet_515) );
NAND2_Z01 cordic_g443 ( .a(cordic_SumAngle_5_), .b(cordic_n_7), .o(cordic_n_64) );
BUF_X2 newInst_916 ( .a(newNet_915), .o(newNet_916) );
BUF_X2 newInst_773 ( .a(newNet_772), .o(newNet_773) );
fflopd cordic_Y_reg_8_ ( .CK(newNet_205), .D(cordic_n_80), .Q(cordic_Y_8_) );
NAND2_Z01 cordic_AddX_Add_g681 ( .a(cordic_AddX_Add_n_52), .b(cordic_AddX_Add_n_30), .o(cordic_AddX_Add_n_53) );
XOR2_X1 cordic_AddY_Add_g703 ( .a(cordic_AddY_Btemp1_5_), .b(cordic_AddY_Atemp_5_), .o(cordic_AddY_Add_n_31) );
BUF_X2 newInst_112 ( .a(newNet_111), .o(newNet_112) );
BUF_X2 newInst_561 ( .a(newNet_560), .o(newNet_561) );
NAND2_Z01 cordic_AddY_MUX_1_g312 ( .a(cordic_BS2_14_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_9) );
BUF_X2 newInst_884 ( .a(newNet_883), .o(newNet_884) );
BUF_X2 newInst_730 ( .a(newNet_729), .o(newNet_730) );
BUF_X2 newInst_236 ( .a(newNet_235), .o(newNet_236) );
NAND2_Z01 cordic_g432 ( .a(cordic_AngleCout), .b(cordic_n_7), .o(cordic_n_75) );
AND2_X1 g334 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_60) );
NAND2_Z01 cordic_AddY_Add_g690 ( .a(cordic_AddY_Add_n_43), .b(cordic_AddY_Add_n_26), .o(cordic_AddY_Add_n_44) );
NAND3_Z1 g15223 ( .a(n_6), .b(n_281), .c(TAR_TRI_D), .o(n_431) );
NAND2_Z01 cordic_Add0_MUX_1_g293 ( .a(cordic_tanangle_6_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_8) );
AND2_X1 g355 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_39) );
NAND2_Z01 g15288 ( .a(n_270), .b(PI_IRDY_L), .o(n_367) );
NAND2_Z01 g14941 ( .a(n_580), .b(n_507), .o(n_633) );
BUF_X2 newInst_240 ( .a(newNet_239), .o(newNet_240) );
XOR2_X1 g15579 ( .a(PI_AD_53), .b(PI_AD_41), .o(n_86) );
BUF_X2 newInst_897 ( .a(newNet_896), .o(newNet_897) );
NAND2_Z01 cordic_AddY_MUX_1_g307 ( .a(cordic_BS2_2_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_14) );
NAND3_Z1 cordic_SH1_srl_35_26_g1116 ( .a(cordic_SH1_srl_35_26_n_114), .b(cordic_SH1_srl_35_26_n_103), .c(cordic_SH1_srl_35_26_n_112), .o(cordic_BS1_6_) );
BUF_X2 newInst_1098 ( .a(newNet_1097), .o(newNet_1098) );
BUF_X2 newInst_819 ( .a(newNet_818), .o(newNet_819) );
NAND2_Z01 cordic_AddX_MUX_1_g287 ( .a(cordic_AddX_MUX_1_n_2), .b(cordic_AddX_MUX_1_n_18), .o(cordic_AddX_Btemp_4_) );
INV_X1 cordic_SH1_srl_35_26_g1152 ( .a(cordic_SH1_srl_35_26_n_95), .o(cordic_SH1_srl_35_26_n_94) );
BUF_X2 newInst_416 ( .a(newNet_415), .o(newNet_416) );
BUF_X2 newInst_22 ( .a(newNet_21), .o(newNet_22) );
NAND2_Z01 cordic_AddY_MUX_1_g308 ( .a(cordic_BS2_1_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_13) );
NAND2_Z01 cordic_Add0_MUX_0_g263 ( .a(cordic_Add0_MUX_0_n_26), .b(cordic_Add0_MUX_0_n_7), .o(cordic_Add0_Atemp_10_) );
BUF_X2 newInst_1151 ( .a(newNet_1150), .o(newNet_1151) );
NAND2_Z01 cordic_AddX_MUX_1_g296 ( .a(cordic_AddX_Y_1), .b(cordic_X_0_), .o(cordic_AddX_MUX_1_n_25) );
NAND2_Z01 cordic_Add0_MUX_0_g271 ( .a(cordic_tanangle_11_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_32) );
NAND2_Z01 g15108 ( .a(n_462), .b(n_461), .o(n_500) );
BUF_X2 newInst_495 ( .a(newNet_494), .o(newNet_495) );
BUF_X2 newInst_455 ( .a(newNet_121), .o(newNet_455) );
NAND2_Z01 cordic_AddX_Add_g697 ( .a(cordic_AddX_Add_n_35), .b(cordic_AddX_Add_n_2), .o(cordic_AddX_Add_n_37) );
NOR2_Z2 cordic_AddX_g66 ( .a(cordic_AddX_Y_3), .b(cordic_AddX_n_0), .o(cordic_AddX_Y_4) );
BUF_X2 newInst_689 ( .a(newNet_688), .o(newNet_689) );
BUF_X2 newInst_542 ( .a(newNet_541), .o(newNet_542) );
NAND2_Z01 cordic_AddY_MUX_0_g293 ( .a(cordic_BS2_12_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_28) );
XOR2_X1 cordic_Add0_Add_g681 ( .a(cordic_Add0_n_11), .b(cordic_Add0_Atemp_10_), .o(cordic_Add0_Add_n_26) );
NAND2_Z01 g15078 ( .a(n_494), .b(PI_AD_12), .o(n_530) );
NAND2_Z01 cordic_SH1_srl_35_26_g1175 ( .a(cordic_SH1_srl_35_26_n_42), .b(cordic_SH1_srl_35_26_n_55), .o(cordic_SH1_srl_35_26_n_77) );
NAND2_Z01 cordic_SH1_srl_35_26_g1159 ( .a(cordic_SH1_srl_35_26_n_83), .b(cordic_SH1_srl_35_26_n_65), .o(cordic_SH1_srl_35_26_n_93) );
NAND2_Z01 cordic_SH2_srl_35_26_g1141 ( .a(cordic_SH2_srl_35_26_n_101), .b(cordic_SH2_srl_35_26_n_20), .o(cordic_SH2_srl_35_26_n_111) );
NAND2_Z01 cordic_pla_g278 ( .a(cordic_pla_n_22), .b(cordic_pla_n_9), .o(cordic_tanangle_6_) );
XOR2_X1 g13394 ( .a(n_885), .b(PO_AD_19), .o(n_886) );
NAND2_Z01 g15091 ( .a(n_4), .b(PI_AD_9), .o(n_517) );
BUF_X2 newInst_119 ( .a(newNet_118), .o(newNet_119) );
BUF_X2 newInst_672 ( .a(newNet_671), .o(newNet_672) );
NAND2_Z01 cordic_SH2_srl_35_26_g1145 ( .a(cordic_SH2_srl_35_26_n_95), .b(cordic_SH2_srl_35_26_n_20), .o(cordic_SH2_srl_35_26_n_107) );
BUF_X2 newInst_793 ( .a(newNet_252), .o(newNet_793) );
BUF_X2 newInst_446 ( .a(newNet_445), .o(newNet_446) );
fflopd Access_Address_1_reg_30_ ( .CK(newNet_1131), .D(n_470), .Q(Access_Address_1_30_) );
BUF_X2 newInst_349 ( .a(newNet_348), .o(newNet_349) );
INV_X1 cordic_SH1_srl_35_26_g1123 ( .a(cordic_SH1_srl_35_26_n_128), .o(cordic_SH1_srl_35_26_n_129) );
INV_X1 cordic_g505 ( .a(CoreOutput_11_), .o(cordic_n_2) );
INV_X2 newInst_46 ( .a(newNet_15), .o(newNet_46) );
INV_X1 cordic_SH1_srl_35_26_g1251 ( .a(cordic_iteration_3_), .o(cordic_SH1_srl_35_26_n_1) );
NAND2_Z01 cordic_SH1_srl_35_26_g1226 ( .a(cordic_iteration_0_), .b(cordic_Y_11_), .o(cordic_SH1_srl_35_26_n_26) );
NAND2_Z01 g13561 ( .a(n_712), .b(CoreOutputReg_15_), .o(n_726) );
BUF_X2 newInst_219 ( .a(newNet_218), .o(newNet_219) );
BUF_X2 newInst_154 ( .a(newNet_6), .o(newNet_154) );
NAND2_Z01 g15405 ( .a(n_214), .b(CoreOutputReg_5_), .o(n_245) );
AND2_X1 cordic_Add0_Compl_g361 ( .a(cordic_Add0_Compl_n_19), .b(cordic_Add0_Compl_n_16), .o(cordic_Add0_Compl_n_21) );
NAND2_Z01 g13534 ( .a(Idsel), .b(Config_Reg_7_), .o(n_752) );
NAND3_Z1 g13424 ( .a(n_853), .b(n_857), .c(n_852), .o(n_1047) );
BUF_X2 newInst_292 ( .a(newNet_291), .o(newNet_292) );
INV_X1 g15194 ( .a(n_446), .o(n_447) );
NAND2_Z01 g15082 ( .a(n_4), .b(PI_AD_15), .o(n_526) );
BUF_X2 newInst_72 ( .a(newNet_71), .o(newNet_72) );
BUF_X2 newInst_126 ( .a(newNet_125), .o(newNet_126) );
NAND2_Z01 cordic_AddX_g65 ( .a(cordic_n_144), .b(cordic_Xsign), .o(cordic_AddX_n_2) );
NAND3_Z1 g15019 ( .a(n_30), .b(n_497), .c(Access_Type_1_1_), .o(n_565) );
NAND2_Z01 g15394 ( .a(n_214), .b(CoreOutputReg_2_), .o(n_256) );
BUF_X2 newInst_820 ( .a(newNet_819), .o(newNet_820) );
XOR2_X1 g15494 ( .a(n_62), .b(n_73), .o(n_169) );
BUF_X2 newInst_315 ( .a(newNet_314), .o(newNet_315) );
INV_X1 g15614 ( .a(n_48), .o(n_47) );
AND2_X1 cordic_SH2_srl_35_26_g1192 ( .a(cordic_SH2_srl_35_26_n_41), .b(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_60) );
NAND2_Z01 cordic_pla_g293 ( .a(cordic_pla_n_15), .b(cordic_pla_n_6), .o(cordic_pla_n_17) );
NAND2_Z01 g15397 ( .a(n_214), .b(CoreOutputReg_31_), .o(n_253) );
BUF_X2 newInst_1042 ( .a(newNet_1041), .o(newNet_1042) );
BUF_X2 newInst_130 ( .a(newNet_129), .o(newNet_130) );
XOR2_X1 g15499 ( .a(n_64), .b(n_65), .o(n_164) );
NAND2_Z01 g15557 ( .a(n_38), .b(State_1_), .o(n_115) );
BUF_X2 newInst_1158 ( .a(newNet_1157), .o(newNet_1158) );
NAND2_Z01 cordic_AddY_MUX_0_g309 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_0_), .o(cordic_AddY_MUX_0_n_12) );
NAND2_Z01 g15463 ( .a(n_145), .b(n_49), .o(n_195) );
AND2_X1 g357 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_37) );
NOR2_Z2 cordic_AddY_g66 ( .a(cordic_AddY_Y_3), .b(cordic_AddY_n_0), .o(cordic_AddY_Y_4) );
BUF_X2 newInst_1062 ( .a(newNet_1061), .o(newNet_1062) );
BUF_X2 newInst_174 ( .a(newNet_173), .o(newNet_174) );
XOR2_X1 cordic_AddY_Compl_g358 ( .a(cordic_AddY_Compl_n_21), .b(cordic_AddY_Compl_n_7), .o(CoreOutput_4_) );
INV_X1 cordic_g408 ( .a(cordic_n_98), .o(cordic_n_99) );
NAND2_Z01 g15515 ( .a(n_103), .b(n_8), .o(n_158) );
NAND2_Z01 cordic_Add0_Add_g668 ( .a(cordic_Add0_Add_n_38), .b(cordic_Add0_Add_n_23), .o(cordic_Add0_Add_n_39) );
XOR2_X1 cordic_Add0_Compl_g350 ( .a(cordic_Add0_Compl_n_29), .b(cordic_Add0_Compl_n_10), .o(cordic_SumAngle_8_) );
NAND2_Z01 cordic_AddX_Add_g726 ( .a(cordic_AddX_Btemp1_15_), .b(cordic_AddX_Atemp_15_), .o(cordic_AddX_Add_n_8) );
INV_X1 cordic_pla_g309 ( .a(cordic_iteration_2_), .o(cordic_pla_n_2) );
INV_X1 cordic_g494 ( .a(CoreOutput_16_), .o(cordic_n_13) );
NAND2_Z01 g15529 ( .a(n_106), .b(n_112), .o(n_125) );
BUF_X2 newInst_271 ( .a(newNet_270), .o(newNet_271) );
NAND2_Z01 cordic_Add0_MUX_0_g297 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_4_), .o(cordic_Add0_MUX_0_n_6) );
BUF_X2 newInst_1188 ( .a(newNet_473), .o(newNet_1188) );
BUF_X2 newInst_82 ( .a(newNet_81), .o(newNet_82) );
NAND2_Z01 cordic_Add0_Add_g654 ( .a(cordic_Add0_Add_n_51), .b(cordic_Add0_Add_n_15), .o(cordic_Add0_Add_n_53) );
INV_X1 cordic_AddY_g36 ( .a(cordic_Ysign), .o(cordic_AddY_n_5) );
BUF_X2 newInst_284 ( .a(newNet_283), .o(newNet_284) );
BUF_X2 newInst_91 ( .a(newNet_90), .o(newNet_91) );
BUF_X2 newInst_15 ( .a(newNet_14), .o(newNet_15) );
BUF_X2 newInst_882 ( .a(newNet_881), .o(newNet_882) );
XOR2_X1 cordic_AddX_Add_g703 ( .a(cordic_AddX_Btemp1_5_), .b(cordic_AddX_Atemp_5_), .o(cordic_AddX_Add_n_31) );
fflopd CoreInput_reg_6_ ( .CK(newNet_749), .D(n_643), .Q(CoreInput_6_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1139 ( .a(cordic_SH1_srl_35_26_n_93), .b(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_113) );
fflopd cordic_Angle_reg_14_ ( .CK(newNet_251), .D(cordic_n_112), .Q(cordic_Angle_14_) );
NAND2_Z01 cordic_Add0_MUX_1_g275 ( .a(cordic_AngleCin), .b(cordic_Angle_6_), .o(cordic_Add0_MUX_1_n_26) );
NOR2_Z1 g13464 ( .a(n_783), .b(n_710), .o(n_818) );
AND2_X1 g340 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_54) );
XOR2_X1 g15584 ( .a(PI_AD_10), .b(PI_AD_2), .o(n_81) );
NAND3_Z1 g15155 ( .a(n_233), .b(n_369), .c(n_10), .o(n_457) );
INV_X1 cordic_g504 ( .a(CoreOutput_22_), .o(cordic_n_3) );
NAND2_Z01 g15056 ( .a(n_473), .b(PI_AD_20), .o(n_552) );
NAND2_Z01 cordic_SH1_srl_35_26_g1237 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_9_), .o(cordic_SH1_srl_35_26_n_12) );
BUF_X2 newInst_407 ( .a(newNet_247), .o(newNet_407) );
NAND2_Z01 cordic_SH2_srl_35_26_g1242 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_7_), .o(cordic_SH2_srl_35_26_n_7) );
NAND2_Z01 cordic_SH1_srl_35_26_g1142 ( .a(cordic_SH1_srl_35_26_n_91), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_110) );
NAND2_Z01 g13478 ( .a(n_729), .b(n_772), .o(n_806) );
BUF_X2 newInst_628 ( .a(newNet_627), .o(newNet_628) );
NAND2_Z01 g15339 ( .a(n_3), .b(PI_AD_31), .o(n_322) );
NAND2_Z01 g14928 ( .a(n_593), .b(n_523), .o(n_646) );
XNOR2_X1 cordic_Add0_Compl_g373 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_10_), .o(cordic_Add0_Compl_n_9) );
BUF_X2 newInst_967 ( .a(newNet_966), .o(newNet_967) );
BUF_X2 newInst_906 ( .a(newNet_905), .o(newNet_906) );
fflopd Access_Address_1_reg_16_ ( .CK(newNet_1190), .D(n_459), .Q(Access_Address_1_16_) );
NAND3_Z1 g14841 ( .a(n_629), .b(n_566), .c(n_10), .o(n_682) );
INV_X2 newInst_187 ( .a(newNet_186), .o(newNet_187) );
NAND3_Z1 g15224 ( .a(n_6), .b(n_281), .c(Idsel), .o(n_430) );
BUF_X2 newInst_876 ( .a(newNet_875), .o(newNet_876) );
BUF_X2 newInst_536 ( .a(newNet_535), .o(newNet_536) );
BUF_X2 newInst_85 ( .a(newNet_84), .o(newNet_85) );
fflopd cordic_Angle_reg_10_ ( .CK(newNet_286), .D(cordic_n_118), .Q(cordic_Angle_10_) );
fflopd cordic_X_reg_4_ ( .CK(newNet_127), .D(cordic_n_51), .Q(cordic_X_4_) );
BUF_X2 newInst_1038 ( .a(newNet_519), .o(newNet_1038) );
AND2_X1 cordic_AddX_Compl_g355 ( .a(cordic_AddX_Compl_n_25), .b(cordic_AddX_Compl_n_4), .o(cordic_AddX_Compl_n_27) );
BUF_X2 newInst_116 ( .a(newNet_115), .o(newNet_116) );
AND2_X1 g349 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_45) );
fflopd cordic_Y_reg_15_ ( .CK(newNet_74), .D(cordic_n_41), .Q(cordic_Y_15_) );
BUF_X2 newInst_1181 ( .a(newNet_77), .o(newNet_1181) );
BUF_X2 newInst_186 ( .a(newNet_185), .o(newNet_186) );
XOR2_X1 g15576 ( .a(PI_CBE_L_3), .b(PI_CBE_L_0), .o(n_89) );
fflopd cordic_X_reg_9_ ( .CK(newNet_572), .D(cordic_n_29), .Q(cordic_X_9_) );
BUF_X2 newInst_718 ( .a(newNet_717), .o(newNet_718) );
NAND2_Z01 cordic_AddY_MUX_1_g282 ( .a(cordic_AddY_MUX_1_n_5), .b(cordic_AddY_MUX_1_n_22), .o(cordic_AddY_Btemp_6_) );
fflopd CoreOutputReg_reg_23_ ( .CK(newNet_640), .D(n_398), .Q(CoreOutputReg_23_) );
NAND2_Z01 g15109 ( .a(n_460), .b(n_384), .o(n_499) );
NAND2_Z01 cordic_pla_g280 ( .a(cordic_pla_n_7), .b(cordic_pla_n_14), .o(cordic_pla_n_30) );
BUF_X2 newInst_1115 ( .a(newNet_1114), .o(newNet_1115) );
XOR2_X1 cordic_Add0_Add_g646 ( .a(cordic_Add0_Add_n_59), .b(cordic_Add0_Add_n_26), .o(cordic_Add0_Stemp_10_) );
BUF_X2 newInst_472 ( .a(newNet_471), .o(newNet_472) );
XNOR2_X1 cordic_AddX_Compl_g372 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_8_), .o(cordic_AddX_Compl_n_10) );
NOR2_Z1 cordic_Add0_MUX_0_g292 ( .a(cordic_Add0_MUX_0_n_0), .b(cordic_AngleCin), .o(cordic_Add0_Atemp_14_) );
BUF_X2 newInst_320 ( .a(newNet_319), .o(newNet_320) );
AND2_X1 cordic_SH2_srl_35_26_g1149 ( .a(cordic_SH2_srl_35_26_n_89), .b(cordic_SH2_srl_35_26_n_1), .o(cordic_SH2_srl_35_26_n_103) );
NOR2_Z1 cordic_SH2_srl_35_26_g1213 ( .a(cordic_SH2_srl_35_26_n_19), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_42) );
XOR2_X1 cordic_AddX_Add_g715 ( .a(cordic_AddX_Btemp1_12_), .b(cordic_AddX_Atemp_12_), .o(cordic_AddX_Add_n_19) );
XOR2_X1 g13416 ( .a(n_863), .b(PO_AD_29), .o(n_864) );
XOR2_X1 cordic_AddX_g206 ( .a(cordic_AddX_Btemp_13_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_13_) );
BUF_X2 newInst_1072 ( .a(newNet_854), .o(newNet_1072) );
NAND2_Z01 g15414 ( .a(n_184), .b(PI_IDSEL), .o(n_236) );
BUF_X2 newInst_1150 ( .a(newNet_1149), .o(newNet_1150) );
fflopd Config_Reg_reg_24_ ( .CK(newNet_943), .D(n_672), .Q(Config_Reg_24_) );
BUF_X2 newInst_592 ( .a(newNet_591), .o(newNet_592) );
BUF_X2 newInst_278 ( .a(newNet_148), .o(newNet_278) );
NAND2_Z01 g13490 ( .a(n_728), .b(n_767), .o(n_794) );
BUF_X2 newInst_1122 ( .a(newNet_0), .o(newNet_1122) );
BUF_X2 newInst_682 ( .a(newNet_681), .o(newNet_682) );
BUF_X2 newInst_910 ( .a(newNet_151), .o(newNet_910) );
BUF_X2 newInst_146 ( .a(newNet_145), .o(newNet_146) );
NAND3_Z1 g15129 ( .a(n_331), .b(n_425), .c(n_10), .o(n_481) );
NAND2_Z01 cordic_SH1_srl_35_26_g1220 ( .a(cordic_iteration_0_), .b(cordic_Y_8_), .o(cordic_SH1_srl_35_26_n_32) );
NAND2_Z01 cordic_AddX_Add_g690 ( .a(cordic_AddX_Add_n_43), .b(cordic_AddX_Add_n_26), .o(cordic_AddX_Add_n_44) );
INV_X1 g15275 ( .a(n_381), .o(n_380) );
BUF_X2 newInst_784 ( .a(newNet_783), .o(newNet_784) );
BUF_X2 newInst_437 ( .a(newNet_436), .o(newNet_437) );
NAND2_Z01 g15272 ( .a(n_312), .b(n_252), .o(n_388) );
NAND2_Z01 cordic_SH1_srl_35_26_g1147 ( .a(cordic_SH1_srl_35_26_n_99), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_105) );
NAND2_Z01 g15016 ( .a(n_500), .b(PAR64_Int), .o(n_566) );
BUF_X2 newInst_451 ( .a(newNet_450), .o(newNet_451) );
XOR2_X1 cordic_AddX_Compl_g350 ( .a(cordic_AddX_Compl_n_29), .b(cordic_AddX_Compl_n_10), .o(CoreOutput_25_) );
BUF_X2 newInst_870 ( .a(newNet_869), .o(newNet_870) );
NAND2_Z01 g15102 ( .a(n_489), .b(n_269), .o(n_506) );
NAND2_Z01 g15516 ( .a(n_94), .b(n_42), .o(n_146) );
BUF_X2 newInst_848 ( .a(newNet_847), .o(newNet_848) );
NAND2_Z01 cordic_g422 ( .a(Issue_Rst), .b(CoreInput_7_), .o(cordic_n_85) );
NAND2_Z01 g15521 ( .a(n_91), .b(n_47), .o(n_142) );
BUF_X2 newInst_995 ( .a(newNet_994), .o(newNet_995) );
NAND2_Z01 g15287 ( .a(n_281), .b(TAR_TRI_T), .o(n_368) );
BUF_X2 newInst_83 ( .a(newNet_82), .o(newNet_83) );
BUF_X2 newInst_1179 ( .a(newNet_1178), .o(newNet_1179) );
NAND3_Z1 g15156 ( .a(n_335), .b(n_428), .c(n_10), .o(n_456) );
fflopd State_reg_2_ ( .CK(newNet_376), .D(n_697), .Q(State_2_) );
NAND2_Z01 cordic_pla_g294 ( .a(cordic_pla_n_13), .b(cordic_pla_n_1), .o(cordic_pla_n_22) );
NOR2_Z1 cordic_g463 ( .a(cordic_n_10), .b(Issue_Rst), .o(cordic_n_44) );
BUF_X2 newInst_752 ( .a(newNet_751), .o(newNet_752) );
XOR2_X1 cordic_AddY_Compl_g350 ( .a(cordic_AddY_Compl_n_29), .b(cordic_AddY_Compl_n_10), .o(CoreOutput_8_) );
NAND2_Z01 g13471 ( .a(n_743), .b(n_769), .o(n_813) );
NAND2_Z01 g15422 ( .a(n_217), .b(n_11), .o(n_277) );
BUF_X2 newInst_259 ( .a(newNet_258), .o(newNet_259) );
XNOR2_X1 cordic_Add0_Compl_g375 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_4_), .o(cordic_Add0_Compl_n_7) );
NAND2_Z01 cordic_AddY_Add_g699 ( .a(cordic_AddY_Add_n_34), .b(cordic_AddY_Add_n_18), .o(cordic_AddY_Add_n_35) );
XOR2_X1 g15487 ( .a(n_83), .b(n_84), .o(n_176) );
XOR2_X1 cordic_Add0_Add_g686 ( .a(cordic_Add0_n_10), .b(cordic_Add0_Atemp_9_), .o(cordic_Add0_Add_n_21) );
BUF_X2 newInst_568 ( .a(newNet_567), .o(newNet_568) );
NAND2_Z01 g14990 ( .a(n_0), .b(CoreInput_9_), .o(n_587) );
BUF_X2 newInst_757 ( .a(newNet_327), .o(newNet_757) );
BUF_X2 newInst_1093 ( .a(newNet_1092), .o(newNet_1093) );
NOR2_Z1 cordic_SH1_srl_35_26_g1213 ( .a(cordic_SH1_srl_35_26_n_19), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_42) );
AND2_X1 cordic_AddX_Compl_g363 ( .a(cordic_AddX_Compl_n_17), .b(cordic_AddX_Compl_n_14), .o(cordic_AddX_Compl_n_19) );
NAND2_Z01 g13482 ( .a(n_726), .b(n_761), .o(n_802) );
fflopd PAR64_Int_d_reg ( .CK(newNet_1205), .D(n_715), .Q(PAR64_Int_d) );
BUF_X2 newInst_324 ( .a(newNet_323), .o(newNet_324) );
AND2_X1 g51 ( .a(n_829), .b(n_856), .o(PO_AD_13) );
NAND3_Z1 g15018 ( .a(n_490), .b(n_491), .c(n_10), .o(n_562) );
NOR2_Z1 g13436 ( .a(n_812), .b(n_710), .o(n_846) );
BUF_X2 newInst_1059 ( .a(newNet_1058), .o(newNet_1059) );
NAND2_Z01 cordic_AddX_Add_g733 ( .a(cordic_AddX_Btemp1_8_), .b(cordic_AddX_Atemp_8_), .o(cordic_AddX_Add_n_1) );
NAND2_Z01 g15351 ( .a(CoreOutput_13_), .b(n_188), .o(n_310) );
BUF_X2 newInst_634 ( .a(newNet_633), .o(newNet_634) );
NAND2_Z01 g13469 ( .a(n_720), .b(n_773), .o(n_815) );
BUF_X2 newInst_598 ( .a(newNet_310), .o(newNet_598) );
NAND2_Z01 g13547 ( .a(n_712), .b(CoreOutputReg_20_), .o(n_739) );
BUF_X2 newInst_975 ( .a(newNet_974), .o(newNet_975) );
NAND3_Z1 cordic_SH1_srl_35_26_g1164 ( .a(cordic_SH1_srl_35_26_n_3), .b(cordic_SH1_srl_35_26_n_46), .c(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_89) );
BUF_X2 newInst_484 ( .a(newNet_483), .o(newNet_484) );
NAND2_Z01 cordic_AddY_MUX_1_g290 ( .a(cordic_AddY_Y_1), .b(cordic_Y_14_), .o(cordic_AddY_MUX_1_n_31) );
NAND3_Z1 g15143 ( .a(n_364), .b(n_358), .c(n_10), .o(n_468) );
fflopd CoreOutputReg_reg_22_ ( .CK(newNet_644), .D(n_399), .Q(CoreOutputReg_22_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1194 ( .a(cordic_SH1_srl_35_26_n_41), .b(cordic_SH1_srl_35_26_n_19), .o(cordic_BS1_15_) );
INV_X1 cordic_g482 ( .a(CoreOutput_8_), .o(cordic_n_25) );
NAND2_Z01 g15630 ( .a(n_26), .b(State_2_), .o(n_37) );
NAND2_Z01 g15510 ( .a(n_116), .b(CBE_par_3_), .o(n_151) );
BUF_X2 newInst_825 ( .a(newNet_824), .o(newNet_825) );
INV_Y3 g15655 ( .a(RESET), .o(n_10) );
NAND2_Z01 g13483 ( .a(n_736), .b(n_774), .o(n_801) );
NAND2_Z01 g15459 ( .a(n_138), .b(PI_CBE_L_0), .o(n_199) );
BUF_X2 newInst_1079 ( .a(newNet_342), .o(newNet_1079) );
BUF_X2 newInst_963 ( .a(newNet_962), .o(newNet_963) );
fflopd cordic_Angle_reg_11_ ( .CK(newNet_277), .D(cordic_n_117), .Q(cordic_Angle_11_) );
INV_X1 g15656 ( .a(PI_CBE_L_1), .o(n_9) );
BUF_X2 newInst_170 ( .a(newNet_169), .o(newNet_170) );
NAND2_Z01 cordic_AddY_MUX_0_g302 ( .a(cordic_BS2_10_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_19) );
NAND2_Z01 cordic_AddY_MUX_0_g299 ( .a(cordic_BS2_6_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_22) );
XOR2_X1 cordic_AddX_Compl_g360 ( .a(cordic_AddX_Compl_n_19), .b(cordic_AddX_Compl_n_16), .o(CoreOutput_20_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1246 ( .a(cordic_SH1_srl_35_26_n_2), .b(cordic_iteration_3_), .o(cordic_SH1_srl_35_26_n_21) );
NAND2_Z01 cordic_AddX_MUX_0_g286 ( .a(cordic_AddX_MUX_0_n_21), .b(cordic_AddX_MUX_0_n_4), .o(cordic_AddX_Atemp_5_) );
NAND2_Z01 g15254 ( .a(n_304), .b(n_305), .o(n_406) );
BUF_X2 newInst_162 ( .a(newNet_161), .o(newNet_162) );
BUF_X2 newInst_705 ( .a(newNet_90), .o(newNet_705) );
XOR2_X1 cordic_AddX_g210 ( .a(cordic_AddX_Btemp_9_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_9_) );
NAND2_Z01 g13506 ( .a(Idsel), .b(Config_Reg_31_), .o(n_780) );
BUF_X2 newInst_879 ( .a(newNet_878), .o(newNet_879) );
NAND2_Z01 cordic_SH1_srl_35_26_g1227 ( .a(cordic_iteration_0_), .b(cordic_Y_6_), .o(cordic_SH1_srl_35_26_n_25) );
BUF_X2 newInst_936 ( .a(newNet_935), .o(newNet_936) );
BUF_X2 newInst_836 ( .a(newNet_835), .o(newNet_836) );
XOR2_X1 cordic_AddY_Add_g709 ( .a(cordic_AddY_Btemp1_15_), .b(cordic_AddY_Atemp_15_), .o(cordic_AddY_Add_n_25) );
BUF_X2 newInst_765 ( .a(newNet_764), .o(newNet_765) );
BUF_X2 newInst_332 ( .a(newNet_331), .o(newNet_332) );
XOR2_X1 g15317 ( .a(n_173), .b(n_167), .o(n_343) );
NAND3_Z1 g15563 ( .a(Access_Type_1_1_), .b(Access_Type_1_0_), .c(Access_Type_1_2_), .o(n_98) );
fflopd CoreInput_reg_16_ ( .CK(newNet_782), .D(n_650), .Q(CoreInput_16_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1156 ( .a(cordic_SH1_srl_35_26_n_86), .b(cordic_SH1_srl_35_26_n_69), .o(cordic_SH1_srl_35_26_n_97) );
AND2_X1 cordic_g475 ( .a(CoreOutput_32_), .b(Issue_Rst), .o(cordic_n_32) );
INV_X1 cordic_SH2_srl_35_26_g1251 ( .a(cordic_iteration_3_), .o(cordic_SH2_srl_35_26_n_1) );
NAND2_Z01 cordic_AddX_MUX_1_g305 ( .a(cordic_BS1_3_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_16) );
BUF_X2 newInst_1067 ( .a(newNet_1066), .o(newNet_1067) );
BUF_X2 newInst_743 ( .a(newNet_742), .o(newNet_743) );
NOR2_Z1 g13445 ( .a(n_803), .b(n_710), .o(n_837) );
NAND2_Z01 g15292 ( .a(n_275), .b(Access_Type_1_2_), .o(n_363) );
NAND2_Z01 g15234 ( .a(n_274), .b(Access_Address_1_21_), .o(n_426) );
BUF_X2 newInst_289 ( .a(newNet_288), .o(newNet_289) );
BUF_X2 newInst_580 ( .a(newNet_219), .o(newNet_580) );
NOR2_Z1 cordic_g452 ( .a(cordic_n_22), .b(Issue_Rst), .o(cordic_n_55) );
BUF_X2 newInst_1046 ( .a(newNet_1045), .o(newNet_1046) );
NAND2_Z01 cordic_AddX_MUX_0_g316 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_6_), .o(cordic_AddX_MUX_0_n_5) );
BUF_X2 newInst_694 ( .a(newNet_607), .o(newNet_694) );
NAND2_Z01 g15298 ( .a(n_272), .b(PI_CBE_L_2), .o(n_357) );
NOR2_Z1 g13455 ( .a(n_790), .b(n_710), .o(n_827) );
NAND2_Z01 g13551 ( .a(n_712), .b(CoreOutputReg_24_), .o(n_735) );
BUF_X2 newInst_697 ( .a(newNet_696), .o(newNet_697) );
BUF_X2 newInst_659 ( .a(newNet_658), .o(newNet_659) );
BUF_X2 newInst_420 ( .a(newNet_419), .o(newNet_420) );
BUF_X2 newInst_208 ( .a(newNet_207), .o(newNet_208) );
BUF_X2 newInst_52 ( .a(newNet_38), .o(newNet_52) );
BUF_X2 newInst_954 ( .a(newNet_953), .o(newNet_954) );
NAND2_Z01 cordic_SH2_srl_35_26_g1175 ( .a(cordic_SH2_srl_35_26_n_42), .b(cordic_SH2_srl_35_26_n_55), .o(cordic_SH2_srl_35_26_n_77) );
BUF_X2 newInst_895 ( .a(newNet_881), .o(newNet_895) );
BUF_X2 newInst_575 ( .a(newNet_574), .o(newNet_575) );
NAND2_Z01 cordic_Add0_MUX_1_g280 ( .a(cordic_AngleCin), .b(cordic_Angle_4_), .o(cordic_Add0_MUX_1_n_21) );
XOR2_X1 cordic_Add0_Compl_g342 ( .a(cordic_Add0_Compl_n_37), .b(cordic_Add0_Compl_n_12), .o(cordic_SumAngle_12_) );
XOR2_X1 cordic_AddX_g203 ( .a(cordic_AddX_Btemp_11_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_11_) );
NAND2_Z01 g13429 ( .a(n_711), .b(PAR_Int_d), .o(n_853) );
BUF_X2 newInst_105 ( .a(newNet_104), .o(newNet_105) );
NOR2_Z1 g15564 ( .a(n_44), .b(Core_Cnt_0_), .o(n_97) );
NAND2_Z01 cordic_SH2_srl_35_26_g1199 ( .a(cordic_SH2_srl_35_26_n_17), .b(cordic_SH2_srl_35_26_n_29), .o(cordic_SH2_srl_35_26_n_53) );
NAND2_Z01 cordic_AddX_MUX_0_g318 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_13_), .o(cordic_AddX_MUX_0_n_3) );
NAND2_Z01 cordic_AddX_Add_g658 ( .a(cordic_AddX_Add_n_74), .b(cordic_AddX_Add_n_10), .o(cordic_AddX_Add_n_76) );
fflopd Check_Add_Parity_reg ( .CK(newNet_1070), .D(n_700), .Q(Check_Add_Parity) );
BUF_X2 newInst_1105 ( .a(newNet_919), .o(newNet_1105) );
NAND3_Z1 g15305 ( .a(n_211), .b(n_196), .c(n_150), .o(n_350) );
BUF_X2 newInst_927 ( .a(newNet_926), .o(newNet_927) );
BUF_X2 newInst_804 ( .a(newNet_803), .o(newNet_804) );
BUF_X2 newInst_367 ( .a(newNet_366), .o(newNet_367) );
NOR2_Z1 g15309 ( .a(n_271), .b(PI_IRDY_L), .o(n_348) );
INV_X1 cordic_Add0_MUX_1_g300 ( .a(cordic_Angle_14_), .o(cordic_Add0_MUX_1_n_1) );
NAND2_Z01 cordic_AddY_MUX_0_g315 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_11_), .o(cordic_AddY_MUX_0_n_6) );
NAND2_Z01 g14960 ( .a(n_572), .b(Config_Reg_26_), .o(n_617) );
INV_X1 cordic_SH2_srl_35_26_g1125 ( .a(cordic_SH2_srl_35_26_n_126), .o(cordic_SH2_srl_35_26_n_127) );
NAND2_Z01 g14985 ( .a(n_571), .b(CoreInput_4_), .o(n_592) );
NAND2_Z01 g15619 ( .a(State_0_), .b(State_2_), .o(n_51) );
NAND3_Z1 cordic_SH2_srl_35_26_g1164 ( .a(cordic_SH2_srl_35_26_n_3), .b(cordic_SH2_srl_35_26_n_46), .c(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_89) );
fflopd CoreOutputReg_reg_18_ ( .CK(newNet_683), .D(n_404), .Q(CoreOutputReg_18_) );
NAND2_Z01 cordic_AddY_Add_g730 ( .a(cordic_AddY_Btemp1_12_), .b(cordic_AddY_Atemp_12_), .o(cordic_AddY_Add_n_4) );
fflopd cordic_Y_reg_3_ ( .CK(newNet_61), .D(cordic_n_50), .Q(cordic_Y_3_) );
NAND2_Z01 cordic_AddY_Add_g684 ( .a(cordic_AddY_Add_n_49), .b(cordic_AddY_Add_n_28), .o(cordic_AddY_Add_n_50) );
AND2_X1 g42 ( .a(n_818), .b(n_856), .o(PO_AD_22) );
XOR2_X1 g15490 ( .a(n_76), .b(n_77), .o(n_173) );
BUF_X2 newInst_76 ( .a(newNet_75), .o(newNet_76) );
BUF_X2 newInst_394 ( .a(newNet_393), .o(newNet_394) );
XOR2_X1 cordic_AddY_g199 ( .a(cordic_AddY_Btemp_12_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_12_) );
BUF_X2 newInst_222 ( .a(newNet_221), .o(newNet_222) );
NOR2_Z2 g15137 ( .a(n_445), .b(n_35), .o(n_494) );
BUF_X2 newInst_777 ( .a(newNet_776), .o(newNet_777) );
BUF_X2 newInst_45 ( .a(newNet_44), .o(newNet_45) );
NAND2_Z01 g13508 ( .a(Idsel), .b(Config_Reg_21_), .o(n_778) );
BUF_X2 newInst_646 ( .a(newNet_645), .o(newNet_646) );
NAND2_Z01 cordic_AddY_MUX_0_g274 ( .a(cordic_AddY_MUX_0_n_28), .b(cordic_AddY_MUX_0_n_11), .o(cordic_AddY_Atemp_12_) );
AND2_X1 g351 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_43) );
NAND2_Z01 cordic_AddX_MUX_0_g303 ( .a(cordic_BS1_4_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_18) );
NAND2_Z01 g15621 ( .a(Trdy_Cnt_En), .b(n_10), .o(n_48) );
BUF_X2 newInst_178 ( .a(newNet_177), .o(newNet_178) );
XNOR2_X1 cordic_Add0_Compl_g368 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_2_), .o(cordic_Add0_Compl_n_14) );
NAND2_Z01 cordic_SH1_srl_35_26_g1241 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_3_), .o(cordic_SH1_srl_35_26_n_8) );
NAND2_Z01 cordic_AddY_MUX_0_g284 ( .a(cordic_AddY_MUX_0_n_20), .b(cordic_AddY_MUX_0_n_3), .o(cordic_AddY_Atemp_13_) );
XOR2_X1 cordic_AddY_g206 ( .a(cordic_AddY_Btemp_13_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_13_) );
BUF_X2 newInst_164 ( .a(newNet_163), .o(newNet_164) );
NAND2_Z01 cordic_SH1_srl_35_26_g1131 ( .a(cordic_SH1_srl_35_26_n_99), .b(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_121) );
NAND2_Z01 cordic_g390 ( .a(cordic_n_73), .b(cordic_n_95), .o(cordic_n_117) );
NOR2_Z1 g13441 ( .a(n_805), .b(n_710), .o(n_841) );
NAND2_Z01 g14918 ( .a(n_603), .b(n_533), .o(n_656) );
NAND2_Z01 cordic_AddY_Add_g655 ( .a(cordic_AddY_Add_n_77), .b(cordic_AddY_Add_n_8), .o(cordic_AddY_Y_3) );
BUF_X2 newInst_335 ( .a(newNet_334), .o(newNet_335) );
XOR2_X1 g15495 ( .a(n_72), .b(n_66), .o(n_168) );
NAND2_Z01 cordic_Add0_Add_g692 ( .a(cordic_Add0_n_8), .b(cordic_Add0_Atemp_7_), .o(cordic_Add0_Add_n_15) );
BUF_X2 newInst_920 ( .a(newNet_460), .o(newNet_920) );
BUF_X2 newInst_521 ( .a(newNet_520), .o(newNet_521) );
NAND2_Z01 g14974 ( .a(n_571), .b(CoreInput_0_), .o(n_603) );
NAND2_Z01 g15341 ( .a(n_214), .b(CoreOutputReg_0_), .o(n_320) );
BUF_X2 newInst_262 ( .a(newNet_261), .o(newNet_262) );
NOR2_Z6 cordic_AddX_g35 ( .a(cordic_n_144), .b(cordic_AddX_n_5), .o(cordic_AddX_Y_1) );
NAND2_Z01 g15328 ( .a(n_3), .b(PI_AD_21), .o(n_333) );
XOR2_X1 g15502 ( .a(n_57), .b(n_71), .o(n_161) );
NAND2_Z01 cordic_AddX_Add_g688 ( .a(cordic_AddX_Add_n_44), .b(cordic_AddX_Add_n_7), .o(cordic_AddX_Add_n_46) );
NAND3_Z1 cordic_pla_g271 ( .a(cordic_pla_n_30), .b(cordic_pla_n_21), .c(cordic_pla_n_9), .o(cordic_tanangle_3_) );
NAND2_Z01 cordic_AddX_Add_g725 ( .a(cordic_AddX_Btemp1_0_), .b(cordic_AddX_Atemp_0_), .o(cordic_AddX_Add_n_9) );
NAND2_Z01 g13557 ( .a(n_712), .b(CoreOutputReg_28_), .o(n_730) );
NOR2_Z1 g15215 ( .a(n_382), .b(n_215), .o(n_448) );
BUF_X2 newInst_978 ( .a(newNet_977), .o(newNet_978) );
fflopd cordic_X_reg_2_ ( .CK(newNet_135), .D(cordic_n_53), .Q(cordic_X_2_) );
NAND3_Z1 g15159 ( .a(n_273), .b(n_368), .c(n_185), .o(n_453) );
fflopd cordic_X_reg_0_ ( .CK(newNet_178), .D(cordic_n_60), .Q(cordic_X_0_) );
NAND2_Z01 cordic_AddY_Add_g726 ( .a(cordic_AddY_Btemp1_15_), .b(cordic_AddY_Atemp_15_), .o(cordic_AddY_Add_n_8) );
AND2_X1 g59 ( .a(n_820), .b(n_856), .o(PO_AD_5) );
NAND2_Z01 cordic_SH1_srl_35_26_g1230 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_13_), .o(cordic_SH1_srl_35_26_n_22) );
fflopd cordic_Y_reg_2_ ( .CK(newNet_62), .D(cordic_n_39), .Q(cordic_Y_2_) );
BUF_X2 newInst_285 ( .a(newNet_284), .o(newNet_285) );
XOR2_X1 cordic_AddY_g211 ( .a(cordic_AddY_Btemp_2_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_2_) );
BUF_X2 newInst_476 ( .a(newNet_475), .o(newNet_476) );
BUF_X2 newInst_302 ( .a(newNet_301), .o(newNet_302) );
BUF_X2 newInst_98 ( .a(newNet_97), .o(newNet_98) );
NAND2_Z01 cordic_AddY_MUX_1_g304 ( .a(cordic_AddY_Y_1), .b(cordic_Y_3_), .o(cordic_AddY_MUX_1_n_17) );
AND2_X1 cordic_g478 ( .a(CoreOutput_26_), .b(Issue_Rst), .o(cordic_n_29) );
NOR2_Z1 g14999 ( .a(n_570), .b(n_202), .o(n_578) );
BUF_X2 newInst_865 ( .a(newNet_864), .o(newNet_865) );
BUF_X2 newInst_27 ( .a(newNet_26), .o(newNet_27) );
NAND2_Z01 g14830 ( .a(n_686), .b(n_138), .o(n_690) );
NOR2_Z1 g14828 ( .a(n_688), .b(n_186), .o(n_692) );
NAND2_Z01 g15209 ( .a(n_381), .b(Par_Sgnl), .o(n_443) );
AND2_X1 g15436 ( .a(n_186), .b(TAR_TRI_S), .o(n_222) );
INV_X1 cordic_SH2_srl_35_26_g1121 ( .a(cordic_SH2_srl_35_26_n_130), .o(cordic_SH2_srl_35_26_n_131) );
NAND2_Z01 g14896 ( .a(n_625), .b(n_554), .o(n_678) );
XOR2_X1 cordic_AddY_Add_g677 ( .a(cordic_AddY_Add_n_55), .b(cordic_AddY_Add_n_17), .o(cordic_AddY_Stemp_8_) );
NAND2_Z01 cordic_g399 ( .a(cordic_n_66), .b(cordic_n_88), .o(cordic_n_108) );
fflopd Access_Type_1_reg_0_ ( .CK(newNet_1110), .D(n_469), .Q(Access_Type_1_0_) );
BUF_X2 newInst_603 ( .a(newNet_602), .o(newNet_603) );
BUF_X2 newInst_56 ( .a(newNet_11), .o(newNet_56) );
BUF_X2 newInst_136 ( .a(newNet_86), .o(newNet_136) );
NAND2_Z01 g14952 ( .a(n_572), .b(Config_Reg_19_), .o(n_625) );
NAND2_Z01 g13497 ( .a(n_741), .b(n_752), .o(n_787) );
BUF_X2 newInst_1136 ( .a(newNet_1135), .o(newNet_1136) );
XOR2_X1 g15580 ( .a(PI_AD_55), .b(PI_AD_50), .o(n_85) );
NAND2_Z01 cordic_AddY_MUX_1_g311 ( .a(cordic_BS2_8_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_10) );
NAND2_Z01 cordic_AddX_MUX_0_g277 ( .a(cordic_AddX_MUX_0_n_26), .b(cordic_AddX_MUX_0_n_10), .o(cordic_AddX_Atemp_8_) );
XOR2_X1 cordic_AddX_Add_g656 ( .a(cordic_AddX_Add_n_76), .b(cordic_AddX_Add_n_25), .o(cordic_AddX_Stemp_15_) );
fflopd cordic_AngleCin_reg ( .CK(newNet_268), .D(cordic_n_116), .Q(cordic_AngleCin) );
XOR2_X1 g13398 ( .a(n_881), .b(PO_AD_22), .o(n_882) );
BUF_X2 newInst_609 ( .a(newNet_608), .o(newNet_609) );
BUF_X2 newInst_327 ( .a(newNet_326), .o(newNet_327) );
XOR2_X1 cordic_AddX_Add_g707 ( .a(cordic_AddX_Btemp1_10_), .b(cordic_AddX_Atemp_10_), .o(cordic_AddX_Add_n_27) );
NAND2_Z01 cordic_Add0_MUX_1_g267 ( .a(cordic_Add0_MUX_1_n_9), .b(cordic_Add0_MUX_1_n_19), .o(cordic_Add0_Btemp_3_) );
NAND2_Z01 g15519 ( .a(n_115), .b(n_10), .o(n_157) );
BUF_X2 newInst_814 ( .a(newNet_813), .o(newNet_814) );
NAND2_Z01 cordic_SH1_srl_35_26_g1165 ( .a(cordic_SH1_srl_35_26_n_54), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_87) );
NOR2_Z1 g15456 ( .a(n_141), .b(OutputAvail), .o(n_202) );
NAND2_Z01 cordic_g410 ( .a(cordic_iteration_0_), .b(cordic_iteration_1_), .o(cordic_n_98) );
NAND2_Z01 g15120 ( .a(n_444), .b(n_217), .o(n_489) );
NAND2_Z01 g15371 ( .a(CoreOutput_31_), .b(n_2), .o(n_290) );
BUF_X2 newInst_664 ( .a(newNet_663), .o(newNet_664) );
NAND2_Z01 cordic_SH2_srl_35_26_g1217 ( .a(cordic_iteration_0_), .b(cordic_X_4_), .o(cordic_SH2_srl_35_26_n_35) );
BUF_X2 newInst_796 ( .a(newNet_795), .o(newNet_796) );
NAND2_Z01 cordic_SH2_srl_35_26_g1113 ( .a(cordic_SH2_srl_35_26_n_126), .b(cordic_iteration_3_), .o(cordic_SH2_srl_35_26_n_139) );
fflopd cordic_X_reg_11_ ( .CK(newNet_39), .D(cordic_n_34), .Q(cordic_X_11_) );
BUF_X2 newInst_639 ( .a(newNet_638), .o(newNet_639) );
NAND2_Z01 g14937 ( .a(n_585), .b(n_513), .o(n_637) );
INV_X1 g15546 ( .a(n_118), .o(n_117) );
BUF_X2 newInst_807 ( .a(newNet_806), .o(newNet_807) );
NAND2_Z01 cordic_SH2_srl_35_26_g1219 ( .a(cordic_iteration_0_), .b(cordic_X_12_), .o(cordic_SH2_srl_35_26_n_33) );
AND2_X1 g63 ( .a(n_846), .b(n_856), .o(PO_AD_1) );
NAND2_Z01 g15454 ( .a(n_45), .b(n_158), .o(n_216) );
INV_X1 cordic_SH2_srl_35_26_g1231 ( .a(cordic_SH2_srl_35_26_n_19), .o(cordic_SH2_srl_35_26_n_18) );
NAND2_Z01 cordic_Add0_MUX_1_g260 ( .a(cordic_Add0_MUX_1_n_10), .b(cordic_Add0_MUX_1_n_29), .o(cordic_Add0_Btemp_7_) );
NAND2_Z01 cordic_Add0_Add_g639 ( .a(cordic_Add0_Add_n_66), .b(cordic_Add0_Add_n_4), .o(cordic_Add0_Add_n_68) );
NOR3_Z1 g15540 ( .a(n_19), .b(n_34), .c(Access_Type_1_3_), .o(n_131) );
BUF_X2 newInst_1054 ( .a(newNet_670), .o(newNet_1054) );
NAND2_Z01 cordic_g414 ( .a(Issue_Rst), .b(CoreInput_14_), .o(cordic_n_93) );
BUF_X2 newInst_1171 ( .a(newNet_1170), .o(newNet_1171) );
NAND2_Z01 cordic_g404 ( .a(cordic_n_61), .b(cordic_n_83), .o(cordic_n_103) );
XOR2_X1 g15610 ( .a(PI_AD_59), .b(PI_AD_47), .o(n_55) );
NAND2_Z01 cordic_AddY_MUX_1_g273 ( .a(cordic_AddY_MUX_1_n_7), .b(cordic_AddY_MUX_1_n_32), .o(cordic_AddY_Btemp_15_) );
BUF_X2 newInst_436 ( .a(newNet_435), .o(newNet_436) );
NAND2_Z01 cordic_Add0_MUX_0_g279 ( .a(cordic_tanangle_13_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_24) );
XNOR2_X1 cordic_AddY_Compl_g372 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_8_), .o(cordic_AddY_Compl_n_10) );
BUF_X2 newInst_887 ( .a(newNet_886), .o(newNet_887) );
INV_X1 g14831 ( .a(n_689), .o(n_688) );
BUF_X2 newInst_250 ( .a(newNet_249), .o(newNet_250) );
NAND2_Z01 cordic_SH2_srl_35_26_g1109 ( .a(cordic_SH2_srl_35_26_n_132), .b(cordic_iteration_3_), .o(cordic_SH2_srl_35_26_n_143) );
XOR2_X1 cordic_AddX_Compl_g337 ( .a(cordic_AddX_Compl_n_43), .b(cordic_AddX_Compl_n_2), .o(CoreOutput_32_) );
NAND2_Z01 cordic_AddX_MUX_0_g302 ( .a(cordic_BS1_10_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_19) );
NAND4_Z1 cordic_SH2_srl_35_26_g1104 ( .a(cordic_SH2_srl_35_26_n_76), .b(cordic_SH2_srl_35_26_n_120), .c(cordic_SH2_srl_35_26_n_145), .d(cordic_SH2_srl_35_26_n_74), .o(cordic_BS2_2_) );
fflopd Dual_Cycle_reg ( .CK(newNet_484), .D(n_365), .Q(Dual_Cycle) );
NAND2_Z01 cordic_AddY_Add_g681 ( .a(cordic_AddY_Add_n_52), .b(cordic_AddY_Add_n_30), .o(cordic_AddY_Add_n_53) );
BUF_X2 newInst_1157 ( .a(newNet_1156), .o(newNet_1157) );
BUF_X2 newInst_280 ( .a(newNet_279), .o(newNet_280) );
NAND2_Z01 g15367 ( .a(n_214), .b(CoreOutputReg_20_), .o(n_294) );
NOR2_Z1 cordic_g429 ( .a(cordic_n_17), .b(Issue_Rst), .o(cordic_n_78) );
NOR2_Z1 g15471 ( .a(n_112), .b(n_133), .o(n_191) );
NAND2_Z01 cordic_AddY_Add_g667 ( .a(cordic_AddY_Add_n_65), .b(cordic_AddY_Add_n_14), .o(cordic_AddY_Add_n_67) );
NAND2_Z01 cordic_SH2_srl_35_26_g1210 ( .a(cordic_SH2_srl_35_26_n_11), .b(cordic_SH2_srl_35_26_n_36), .o(cordic_SH2_srl_35_26_n_44) );
AND2_X1 g36 ( .a(n_838), .b(n_856), .o(PO_AD_28) );
NAND2_Z01 cordic_AddX_MUX_1_g309 ( .a(cordic_BS1_0_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_12) );
NAND2_Z01 cordic_Add0_MUX_1_g297 ( .a(cordic_tanangle_12_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_4) );
NAND2_Z01 g14817 ( .a(n_695), .b(Trdy_Cnt_En), .o(n_702) );
BUF_X2 newInst_319 ( .a(newNet_318), .o(newNet_319) );
BUF_X2 newInst_61 ( .a(newNet_60), .o(newNet_61) );
BUF_X2 newInst_461 ( .a(newNet_9), .o(newNet_461) );
fflopd cordic_Y_reg_0_ ( .CK(newNet_110), .D(cordic_n_47), .Q(cordic_Y_0_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1229 ( .a(cordic_iteration_0_), .b(cordic_X_2_), .o(cordic_SH2_srl_35_26_n_23) );
AND2_X1 cordic_AddY_Compl_g343 ( .a(cordic_AddY_Compl_n_37), .b(cordic_AddY_Compl_n_12), .o(cordic_AddY_Compl_n_39) );
AND2_X1 g15470 ( .a(n_127), .b(System_Busy), .o(n_192) );
NAND2_Z01 cordic_SH2_srl_35_26_g1206 ( .a(cordic_SH2_srl_35_26_n_5), .b(cordic_SH2_srl_35_26_n_27), .o(cordic_SH2_srl_35_26_n_47) );
NOR2_Z1 cordic_g470 ( .a(cordic_n_5), .b(Issue_Rst), .o(cordic_n_37) );
INV_Z1 cordic_Add0_g55 ( .a(cordic_Add0_Btemp_6_), .o(cordic_Add0_n_7) );
XOR2_X1 g15594 ( .a(PI_AD_58), .b(PI_AD_48), .o(n_71) );
NAND2_Z01 g15096 ( .a(n_473), .b(PI_AD_11), .o(n_512) );
NAND2_Z01 cordic_SH1_srl_35_26_g1135 ( .a(cordic_SH1_srl_35_26_n_92), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_117) );
XNOR2_X1 cordic_AddY_Compl_g368 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_2_), .o(cordic_AddY_Compl_n_14) );
BUF_X2 newInst_127 ( .a(newNet_86), .o(newNet_127) );
NAND2_Z01 cordic_AddX_Add_g666 ( .a(cordic_AddX_Add_n_67), .b(cordic_AddX_Add_n_19), .o(cordic_AddX_Add_n_68) );
BUF_X2 newInst_1094 ( .a(newNet_1093), .o(newNet_1094) );
NAND2_Z01 cordic_SH2_srl_35_26_g1236 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_10_), .o(cordic_SH2_srl_35_26_n_13) );
BUF_X2 newInst_41 ( .a(newNet_40), .o(newNet_41) );
NAND2_Z01 cordic_AddY_MUX_1_g303 ( .a(cordic_AddY_Y_1), .b(cordic_Y_4_), .o(cordic_AddY_MUX_1_n_18) );
BUF_X2 newInst_1013 ( .a(newNet_1012), .o(newNet_1013) );
XOR2_X1 g13409 ( .a(n_870), .b(PO_AD_8), .o(n_871) );
NAND2_Z01 g13501 ( .a(n_748), .b(n_749), .o(n_783) );
fflopd Access_Address_1_reg_22_ ( .CK(newNet_1168), .D(n_481), .Q(Access_Address_1_22_) );
fflopd cordic_Y_reg_14_ ( .CK(newNet_80), .D(cordic_n_42), .Q(cordic_Y_14_) );
AND2_X1 g338 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_56) );
NAND2_Z01 cordic_AddY_Add_g733 ( .a(cordic_AddY_Btemp1_8_), .b(cordic_AddY_Atemp_8_), .o(cordic_AddY_Add_n_1) );
NAND2_Z01 cordic_Add0_Add_g663 ( .a(cordic_Add0_Add_n_42), .b(cordic_Add0_Add_n_8), .o(cordic_Add0_Add_n_44) );
NAND2_Z01 g15398 ( .a(n_214), .b(CoreOutputReg_32_), .o(n_252) );
NAND2_Z01 cordic_Add0_Add_g662 ( .a(cordic_Add0_Add_n_44), .b(cordic_Add0_Add_n_27), .o(cordic_Add0_Add_n_45) );
INV_X1 cordic_Add0_MUX_0_g303 ( .a(cordic_Angle_14_), .o(cordic_Add0_MUX_0_n_0) );
NAND2_Z01 cordic_Add0_Add_g703 ( .a(cordic_Add0_n_13), .b(cordic_Add0_Atemp_12_), .o(cordic_Add0_Add_n_4) );
AND2_X1 g15637 ( .a(Access_Address_1_16_), .b(Access_Address_1_17_), .o(n_27) );
BUF_X2 newInst_358 ( .a(newNet_357), .o(newNet_358) );
NAND4_Z1 cordic_SH1_srl_35_26_g1104 ( .a(cordic_SH1_srl_35_26_n_76), .b(cordic_SH1_srl_35_26_n_120), .c(cordic_SH1_srl_35_26_n_145), .d(cordic_SH1_srl_35_26_n_74), .o(cordic_BS1_2_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1183 ( .a(cordic_SH2_srl_35_26_n_48), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_69) );
BUF_X2 newInst_982 ( .a(newNet_981), .o(newNet_982) );
BUF_X2 newInst_547 ( .a(newNet_546), .o(newNet_547) );
NAND2_Z01 g13544 ( .a(n_712), .b(CoreOutputReg_21_), .o(n_742) );
BUF_X2 newInst_31 ( .a(newNet_30), .o(newNet_31) );
NAND2_Z01 g15335 ( .a(n_218), .b(n_178), .o(n_326) );
NAND2_Z01 g15363 ( .a(n_214), .b(CoreOutputReg_19_), .o(n_298) );
XOR2_X1 cordic_Add0_Add_g688 ( .a(cordic_Add0_n_13), .b(cordic_Add0_Atemp_12_), .o(cordic_Add0_Add_n_19) );
NAND2_Z01 cordic_Add0_MUX_0_g267 ( .a(cordic_Add0_MUX_0_n_22), .b(cordic_Add0_MUX_0_n_6), .o(cordic_Add0_Atemp_4_) );
BUF_X2 newInst_442 ( .a(newNet_441), .o(newNet_442) );
NAND2_Z01 cordic_Add0_Add_g641 ( .a(cordic_Add0_Add_n_65), .b(cordic_Add0_Add_n_19), .o(cordic_Add0_Add_n_66) );
fflopd cordic_Angle_reg_7_ ( .CK(newNet_217), .D(cordic_n_104), .Q(cordic_Angle_7_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1153 ( .a(cordic_SH2_srl_35_26_n_67), .b(cordic_SH2_srl_35_26_n_38), .o(cordic_SH2_srl_35_26_n_101) );
NAND2_Z01 cordic_AddY_Add_g669 ( .a(cordic_AddY_Add_n_64), .b(cordic_AddY_Add_n_29), .o(cordic_AddY_Add_n_65) );
BUF_X2 newInst_447 ( .a(newNet_15), .o(newNet_447) );
NAND2_Z01 cordic_AddX_MUX_1_g283 ( .a(cordic_AddX_MUX_1_n_9), .b(cordic_AddX_MUX_1_n_31), .o(cordic_AddX_Btemp_14_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1127 ( .a(cordic_SH1_srl_35_26_n_95), .b(cordic_iteration_2_), .o(cordic_SH1_srl_35_26_n_125) );
NAND2_Z01 cordic_Add0_MUX_1_g279 ( .a(cordic_AngleCin), .b(cordic_Angle_12_), .o(cordic_Add0_MUX_1_n_22) );
BUF_X2 newInst_917 ( .a(newNet_355), .o(newNet_917) );
BUF_X2 newInst_489 ( .a(newNet_488), .o(newNet_489) );
BUF_X2 newInst_458 ( .a(newNet_457), .o(newNet_458) );
NAND2_Z01 cordic_SH1_srl_35_26_g1242 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_7_), .o(cordic_SH1_srl_35_26_n_7) );
NAND2_Z01 cordic_AddX_MUX_0_g311 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_8_), .o(cordic_AddX_MUX_0_n_10) );
XOR2_X1 cordic_AddY_Add_g718 ( .a(cordic_AddY_Btemp1_0_), .b(cordic_AddY_Atemp_0_), .o(cordic_AddY_Add_n_16) );
AND2_X1 g61 ( .a(n_849), .b(n_856), .o(PO_AD_3) );
AND3_X1 g15570 ( .a(n_12), .b(n_39), .c(Trdy_Wait_Cnt_3_), .o(n_94) );
BUF_X2 newInst_425 ( .a(newNet_424), .o(newNet_425) );
BUF_X2 newInst_1133 ( .a(newNet_1132), .o(newNet_1133) );
BUF_X2 newInst_1144 ( .a(newNet_191), .o(newNet_1144) );
NAND2_Z01 g15092 ( .a(n_455), .b(n_433), .o(n_516) );
BUF_X2 newInst_66 ( .a(newNet_65), .o(newNet_66) );
BUF_X2 newInst_1165 ( .a(newNet_1164), .o(newNet_1165) );
BUF_X2 newInst_614 ( .a(newNet_613), .o(newNet_614) );
NAND2_Z01 g13565 ( .a(n_712), .b(CoreOutputReg_9_), .o(n_722) );
BUF_X2 newInst_776 ( .a(newNet_156), .o(newNet_776) );
NAND2_Z01 cordic_AddX_Add_g676 ( .a(cordic_AddX_Add_n_56), .b(cordic_AddX_Add_n_1), .o(cordic_AddX_Add_n_58) );
BUF_X2 newInst_724 ( .a(newNet_696), .o(newNet_724) );
NOR2_Z1 g15537 ( .a(n_114), .b(PI_FRAME_L), .o(n_122) );
BUF_X2 newInst_152 ( .a(newNet_151), .o(newNet_152) );
BUF_X2 newInst_78 ( .a(newNet_77), .o(newNet_78) );
fflopd CoreInput_reg_3_ ( .CK(newNet_767), .D(n_646), .Q(CoreInput_3_) );
INV_X1 cordic_SH1_srl_35_26_g1204 ( .a(cordic_SH1_srl_35_26_n_41), .o(cordic_SH1_srl_35_26_n_40) );
fflopd CoreInput_reg_14_ ( .CK(newNet_794), .D(n_651), .Q(CoreInput_14_) );
BUF_X2 newInst_9 ( .a(newNet_8), .o(newNet_9) );
NAND2_Z01 cordic_AddY_Add_g729 ( .a(cordic_AddY_Btemp1_9_), .b(cordic_AddY_Atemp_9_), .o(cordic_AddY_Add_n_5) );
NAND2_Z01 cordic_Add0_Add_g630 ( .a(cordic_Add0_Add_n_75), .b(cordic_Add0_Add_n_10), .o(cordic_Add0_Y_3) );
BUF_X2 newInst_1081 ( .a(newNet_1080), .o(newNet_1081) );
NAND2_Z01 g15064 ( .a(n_473), .b(PI_AD_27), .o(n_544) );
NAND2_Z01 g15244 ( .a(n_274), .b(Access_Address_1_30_), .o(n_416) );
NAND2_Z01 cordic_pla_g288 ( .a(cordic_pla_n_4), .b(cordic_pla_n_1), .o(cordic_pla_n_21) );
INV_X1 drc_bufs15665 ( .a(n_6), .o(n_3) );
INV_X1 g15383 ( .a(n_268), .o(n_269) );
BUF_X2 newInst_539 ( .a(newNet_538), .o(newNet_539) );
NAND2_Z01 cordic_AddY_MUX_0_g319 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_4_), .o(cordic_AddY_MUX_0_n_2) );
AND2_X1 g337 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_57) );
BUF_X2 newInst_417 ( .a(newNet_30), .o(newNet_417) );
NAND2_Z01 cordic_AddY_g63 ( .a(cordic_AddY_n_3), .b(cordic_AddY_n_2), .o(CoreOutput_16_) );
BUF_X2 newInst_1061 ( .a(newNet_1060), .o(newNet_1061) );
AND2_X1 cordic_AddX_Compl_g343 ( .a(cordic_AddX_Compl_n_37), .b(cordic_AddX_Compl_n_12), .o(cordic_AddX_Compl_n_39) );
NOR2_Z1 cordic_pla_g290 ( .a(cordic_pla_n_4), .b(cordic_pla_n_8), .o(cordic_pla_n_19) );
NAND2_Z01 cordic_SH2_srl_35_26_g1209 ( .a(cordic_SH2_srl_35_26_n_14), .b(cordic_SH2_srl_35_26_n_25), .o(cordic_SH2_srl_35_26_n_45) );
BUF_X2 newInst_54 ( .a(newNet_53), .o(newNet_54) );
BUF_X2 newInst_707 ( .a(newNet_706), .o(newNet_707) );
BUF_X2 newInst_445 ( .a(newNet_444), .o(newNet_445) );
NAND2_Z01 cordic_AddY_MUX_1_g306 ( .a(cordic_BS2_9_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_15) );
BUF_X2 newInst_456 ( .a(newNet_455), .o(newNet_456) );
NAND2_Z01 cordic_Add0_Add_g651 ( .a(cordic_Add0_Add_n_54), .b(cordic_Add0_Add_n_1), .o(cordic_Add0_Add_n_56) );
BUF_X2 newInst_1131 ( .a(newNet_1130), .o(newNet_1131) );
NAND2_Z01 g15418 ( .a(n_213), .b(Trdy_Wait_Cnt_2_), .o(n_232) );
BUF_X2 newInst_440 ( .a(newNet_439), .o(newNet_440) );
BUF_X2 newInst_885 ( .a(newNet_884), .o(newNet_885) );
NAND2_Z01 cordic_AddX_MUX_1_g288 ( .a(cordic_AddX_MUX_1_n_16), .b(cordic_AddX_MUX_1_n_17), .o(cordic_AddX_Btemp_3_) );
BUF_X2 newInst_914 ( .a(newNet_913), .o(newNet_914) );
INV_X1 drc_bufs15696 ( .a(n_116), .o(n_5) );
BUF_X2 newInst_951 ( .a(newNet_950), .o(newNet_951) );
BUF_X2 newInst_382 ( .a(newNet_381), .o(newNet_382) );
BUF_X2 newInst_373 ( .a(newNet_372), .o(newNet_373) );
AND2_X1 g352 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_42) );
BUF_X2 newInst_546 ( .a(newNet_545), .o(newNet_546) );
INV_X2 newInst_1033 ( .a(newNet_1032), .o(newNet_1033) );
BUF_X2 newInst_1076 ( .a(newNet_1075), .o(newNet_1076) );
NOR2_Z1 cordic_SH2_srl_35_26_g1211 ( .a(cordic_SH2_srl_35_26_n_19), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_43) );
NAND2_Z01 cordic_g406 ( .a(cordic_n_99), .b(cordic_iteration_2_), .o(cordic_n_101) );
BUF_X2 newInst_930 ( .a(newNet_880), .o(newNet_930) );
BUF_X2 newInst_388 ( .a(newNet_120), .o(newNet_388) );
NAND2_Z01 g15212 ( .a(n_360), .b(n_186), .o(n_440) );
INV_X2 cordic_AddY_drc_bufs ( .a(cordic_AddY_n_0), .o(cordic_AddY_Y_2) );
XNOR2_X1 cordic_g407 ( .a(cordic_iteration_0_), .b(cordic_iteration_1_), .o(cordic_n_100) );
BUF_X2 newInst_593 ( .a(newNet_592), .o(newNet_593) );
XOR2_X1 g13391 ( .a(n_888), .b(PO_AD_2), .o(n_889) );
BUF_X2 newInst_806 ( .a(newNet_805), .o(newNet_806) );
XOR2_X1 g15598 ( .a(PI_AD_22), .b(PI_AD_4), .o(n_67) );
BUF_X2 newInst_1199 ( .a(newNet_627), .o(newNet_1199) );
BUF_X2 newInst_760 ( .a(newNet_759), .o(newNet_760) );
XOR2_X1 cordic_g334 ( .a(cordic_n_101), .b(cordic_iteration_3_), .o(cordic_n_121) );
NAND2_Z01 g15379 ( .a(CoreOutput_25_), .b(n_188), .o(n_282) );
NOR2_Z1 cordic_pla_g273 ( .a(cordic_pla_n_23), .b(cordic_iteration_2_), .o(cordic_tanangle_13_) );
NAND2_Z01 g15554 ( .a(n_47), .b(n_39), .o(n_102) );
NAND2_Z01 cordic_SH1_srl_35_26_g1225 ( .a(cordic_iteration_0_), .b(cordic_Y_7_), .o(cordic_SH1_srl_35_26_n_27) );
INV_X2 newInst_845 ( .a(newNet_390), .o(newNet_845) );
BUF_X2 newInst_813 ( .a(newNet_812), .o(newNet_813) );
NAND2_Z01 cordic_AddX_MUX_0_g294 ( .a(cordic_BS1_1_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_27) );
BUF_X2 newInst_562 ( .a(newNet_561), .o(newNet_562) );
BUF_X2 newInst_333 ( .a(newNet_332), .o(newNet_333) );
AND2_X1 cordic_AddY_Compl_g353 ( .a(cordic_AddY_Compl_n_27), .b(cordic_AddY_Compl_n_6), .o(cordic_AddY_Compl_n_29) );
NAND2_Z01 cordic_AddY_MUX_1_g313 ( .a(cordic_BS2_7_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_8) );
NAND2_Z01 g13513 ( .a(Idsel), .b(Config_Reg_6_), .o(n_773) );
NAND2_Z01 cordic_AddX_Add_g694 ( .a(cordic_AddX_Add_n_38), .b(cordic_AddX_Add_n_3), .o(cordic_AddX_Add_n_40) );
NAND2_Z01 g15117 ( .a(n_430), .b(n_236), .o(n_492) );
NAND2_Z01 cordic_Add0_Add_g636 ( .a(cordic_Add0_Add_n_69), .b(cordic_Add0_Add_n_12), .o(cordic_Add0_Add_n_71) );
NAND4_Z1 cordic_SH2_srl_35_26_g1105 ( .a(cordic_SH2_srl_35_26_n_68), .b(cordic_SH2_srl_35_26_n_117), .c(cordic_SH2_srl_35_26_n_144), .d(cordic_SH2_srl_35_26_n_73), .o(cordic_BS2_1_) );
fflopd cordic_Angle_reg_5_ ( .CK(newNet_233), .D(cordic_n_106), .Q(cordic_Angle_5_) );
AND2_X1 g15534 ( .a(n_115), .b(RESET), .o(n_137) );
NAND2_Z01 g15409 ( .a(CoreOutput_7_), .b(n_188), .o(n_241) );
NAND2_Z01 g15079 ( .a(n_4), .b(PI_AD_13), .o(n_529) );
BUF_X2 newInst_1141 ( .a(newNet_1140), .o(newNet_1141) );
BUF_X2 newInst_73 ( .a(newNet_29), .o(newNet_73) );
NAND4_Z1 cordic_SH1_srl_35_26_g1103 ( .a(cordic_SH1_srl_35_26_n_78), .b(cordic_SH1_srl_35_26_n_122), .c(cordic_SH1_srl_35_26_n_139), .d(cordic_SH1_srl_35_26_n_77), .o(cordic_BS1_3_) );
NAND2_Z01 cordic_Add0_MUX_1_g272 ( .a(cordic_AngleCin), .b(cordic_Angle_7_), .o(cordic_Add0_MUX_1_n_29) );
BUF_X2 newInst_903 ( .a(newNet_902), .o(newNet_903) );
NOR2_Z1 g15476 ( .a(n_136), .b(n_113), .o(n_189) );
AND2_X1 cordic_AddX_Compl_g339 ( .a(cordic_AddX_Compl_n_41), .b(cordic_AddX_Compl_n_13), .o(cordic_AddX_Compl_n_43) );
XOR2_X1 cordic_AddX_Compl_g340 ( .a(cordic_AddX_Compl_n_39), .b(cordic_AddX_Compl_n_8), .o(CoreOutput_30_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1138 ( .a(cordic_SH1_srl_35_26_n_96), .b(cordic_SH1_srl_35_26_n_18), .o(cordic_SH1_srl_35_26_n_114) );
AND2_X1 g13425 ( .a(n_854), .b(PI_REQ64_L), .o(n_857) );
NOR2_Z1 g13451 ( .a(n_792), .b(n_710), .o(n_831) );
AND2_X1 g54 ( .a(n_841), .b(n_856), .o(PO_AD_10) );
NAND2_Z01 cordic_g401 ( .a(cordic_n_64), .b(cordic_n_86), .o(cordic_n_106) );
BUF_X2 newInst_1201 ( .a(newNet_1200), .o(newNet_1201) );
NAND2_Z01 cordic_AddX_Add_g719 ( .a(cordic_AddX_Btemp1_7_), .b(cordic_AddX_Atemp_7_), .o(cordic_AddX_Add_n_15) );
XOR2_X1 g15591 ( .a(PI_AD_25), .b(PI_AD_8), .o(n_74) );
NAND2_Z01 cordic_Add0_Add_g642 ( .a(cordic_Add0_Add_n_63), .b(cordic_Add0_Add_n_14), .o(cordic_Add0_Add_n_65) );
BUF_X2 newInst_1189 ( .a(newNet_1188), .o(newNet_1189) );
NAND2_Z01 g14924 ( .a(n_596), .b(n_504), .o(n_650) );
AND2_X1 g345 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_49) );
BUF_X2 newInst_673 ( .a(newNet_262), .o(newNet_673) );
BUF_X2 newInst_494 ( .a(newNet_493), .o(newNet_494) );
BUF_X2 newInst_431 ( .a(newNet_172), .o(newNet_431) );
NAND2_Z01 cordic_g437 ( .a(cordic_SumAngle_14_), .b(cordic_n_7), .o(cordic_n_70) );
NAND2_Z01 g14929 ( .a(n_592), .b(n_522), .o(n_645) );
BUF_X2 newInst_1202 ( .a(newNet_1135), .o(newNet_1202) );
INV_Z1 g8018 ( .a(State_2_), .o(n_898) );
NOR2_Z1 g15468 ( .a(n_139), .b(Dual_Cycle), .o(n_193) );
BUF_X2 newInst_12 ( .a(newNet_11), .o(newNet_12) );
BUF_X2 newInst_1193 ( .a(newNet_1192), .o(newNet_1193) );
BUF_X2 newInst_1126 ( .a(newNet_1125), .o(newNet_1126) );
BUF_X2 newInst_316 ( .a(newNet_315), .o(newNet_316) );
BUF_X2 newInst_88 ( .a(newNet_87), .o(newNet_88) );
NAND2_Z01 cordic_SH1_srl_35_26_g1174 ( .a(cordic_SH1_srl_35_26_n_43), .b(cordic_SH1_srl_35_26_n_45), .o(cordic_SH1_srl_35_26_n_78) );
NAND2_Z01 g15402 ( .a(CoreOutput_3_), .b(n_2), .o(n_248) );
BUF_X2 newInst_17 ( .a(newNet_2), .o(newNet_17) );
BUF_X2 newInst_1099 ( .a(newNet_1098), .o(newNet_1099) );
BUF_X2 newInst_317 ( .a(newNet_316), .o(newNet_317) );
BUF_X2 newInst_21 ( .a(newNet_20), .o(newNet_21) );
INV_X1 g15652 ( .a(DevSel_Wait_Cnt_2_), .o(n_13) );
BUF_X2 newInst_1004 ( .a(newNet_496), .o(newNet_1004) );
BUF_X2 newInst_260 ( .a(newNet_259), .o(newNet_260) );
BUF_X2 newInst_111 ( .a(newNet_96), .o(newNet_111) );
BUF_X2 newInst_49 ( .a(newNet_48), .o(newNet_49) );
BUF_X2 newInst_1182 ( .a(newNet_1181), .o(newNet_1182) );
INV_X1 cordic_g480 ( .a(cordic_AddX_Stemp_0_), .o(cordic_n_27) );
BUF_X2 newInst_242 ( .a(newNet_241), .o(newNet_242) );
NAND2_Z01 g15462 ( .a(n_138), .b(PI_CBE_L_1), .o(n_196) );
NAND2_Z01 cordic_AddX_MUX_0_g287 ( .a(cordic_AddX_MUX_0_n_18), .b(cordic_AddX_MUX_0_n_2), .o(cordic_AddX_Atemp_4_) );
NAND2_Z01 g15393 ( .a(CoreOutput_2_), .b(n_2), .o(n_257) );
NAND2_Z01 cordic_AddX_Add_g729 ( .a(cordic_AddX_Btemp1_9_), .b(cordic_AddX_Atemp_9_), .o(cordic_AddX_Add_n_5) );
BUF_X2 newInst_214 ( .a(newNet_213), .o(newNet_214) );
NAND2_Z01 g14895 ( .a(n_627), .b(n_555), .o(n_679) );
NAND2_Z01 g15069 ( .a(n_473), .b(PI_AD_31), .o(n_539) );
NAND2_Z01 cordic_Add0_Add_g699 ( .a(cordic_Add0_n_5), .b(cordic_Add0_Atemp_4_), .o(cordic_Add0_Add_n_8) );
NAND2_Z01 cordic_AddX_MUX_1_g290 ( .a(cordic_AddX_Y_1), .b(cordic_X_14_), .o(cordic_AddX_MUX_1_n_31) );
BUF_X2 newInst_385 ( .a(newNet_384), .o(newNet_385) );
BUF_X2 newInst_97 ( .a(newNet_96), .o(newNet_97) );
NAND2_Z01 g14911 ( .a(n_609), .b(n_536), .o(n_663) );
NAND2_Z01 cordic_SH1_srl_35_26_g1190 ( .a(cordic_SH1_srl_35_26_n_52), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_62) );
NAND2_Z01 cordic_SH1_srl_35_26_g1172 ( .a(cordic_SH1_srl_35_26_n_47), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_80) );
BUF_X2 newInst_306 ( .a(newNet_305), .o(newNet_306) );
BUF_X2 newInst_165 ( .a(newNet_164), .o(newNet_165) );
INV_X1 cordic_Add0_Compl_g382 ( .a(cordic_AngleCout), .o(cordic_Add0_Compl_n_0) );
NAND2_Z01 cordic_AddX_MUX_0_g304 ( .a(cordic_BS1_3_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_17) );
NAND2_Z01 cordic_AddY_Add_g727 ( .a(cordic_AddY_Btemp1_4_), .b(cordic_AddY_Atemp_4_), .o(cordic_AddY_Add_n_7) );
AND2_X1 g41 ( .a(n_822), .b(n_856), .o(PO_AD_23) );
NAND2_Z01 cordic_SH1_srl_35_26_g1203 ( .a(cordic_SH1_srl_35_26_n_22), .b(cordic_SH1_srl_35_26_n_31), .o(cordic_SH1_srl_35_26_n_50) );
NAND3_Z1 g15532 ( .a(Access_Type_1_3_), .b(n_36), .c(Idsel), .o(n_124) );
BUF_X2 newInst_524 ( .a(newNet_523), .o(newNet_524) );
NAND2_Z01 g15089 ( .a(n_494), .b(PI_AD_7), .o(n_519) );
AND2_X1 g15219 ( .a(n_381), .b(n_193), .o(n_446) );
BUF_X2 newInst_787 ( .a(newNet_786), .o(newNet_787) );
BUF_X2 newInst_210 ( .a(newNet_209), .o(newNet_210) );
NAND2_Z01 cordic_g426 ( .a(Issue_Rst), .b(CoreInput_10_), .o(cordic_n_81) );
BUF_X2 newInst_821 ( .a(newNet_820), .o(newNet_821) );
INV_X1 cordic_pla_g305 ( .a(cordic_pla_n_6), .o(cordic_pla_n_5) );
NAND3_Z1 cordic_SH2_srl_35_26_g1118 ( .a(cordic_SH2_srl_35_26_n_105), .b(cordic_SH2_srl_35_26_n_107), .c(cordic_SH2_srl_35_26_n_104), .o(cordic_BS2_4_) );
BUF_X2 newInst_59 ( .a(newNet_58), .o(newNet_59) );
BUF_X2 newInst_69 ( .a(newNet_68), .o(newNet_69) );
BUF_X2 newInst_255 ( .a(newNet_111), .o(newNet_255) );
XOR2_X1 g15501 ( .a(n_58), .b(n_59), .o(n_162) );
XOR2_X1 cordic_Add0_Add_g691 ( .a(cordic_Add0_Add_n_0), .b(cordic_Add0_Atemp_0_), .o(cordic_Add0_Stemp_0_) );
BUF_X2 newInst_424 ( .a(newNet_423), .o(newNet_424) );
XOR2_X1 g13405 ( .a(n_874), .b(PO_AD_9), .o(n_875) );
NAND2_Z01 cordic_AddX_Add_g687 ( .a(cordic_AddX_Add_n_46), .b(cordic_AddX_Add_n_31), .o(cordic_AddX_Add_n_47) );
XOR2_X1 g15545 ( .a(n_52), .b(Core_Cnt_2_), .o(n_119) );
BUF_X2 newInst_860 ( .a(newNet_362), .o(newNet_860) );
NOR2_Z1 g13460 ( .a(n_786), .b(n_710), .o(n_822) );
XOR2_X1 cordic_AddY_Compl_g371 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_1_), .o(cordic_AddY_Compl_n_11) );
BUF_X2 newInst_360 ( .a(newNet_359), .o(newNet_360) );
BUF_X2 newInst_33 ( .a(newNet_32), .o(newNet_33) );
NAND2_Z01 g14827 ( .a(n_689), .b(n_147), .o(n_693) );
BUF_X2 newInst_778 ( .a(newNet_777), .o(newNet_778) );
NOR2_Z1 cordic_pla_g301 ( .a(cordic_pla_n_2), .b(cordic_iteration_1_), .o(cordic_pla_n_10) );
BUF_X2 newInst_984 ( .a(newNet_238), .o(newNet_984) );
fflopd CoreOutputReg_reg_27_ ( .CK(newNet_622), .D(n_394), .Q(CoreOutputReg_27_) );
fflopd DevSel_Wait_Cnt_reg_0_ ( .CK(newNet_507), .D(n_454), .Q(DevSel_Wait_Cnt_0_) );
BUF_X2 newInst_771 ( .a(newNet_770), .o(newNet_771) );
NAND2_Z02 g15008 ( .a(n_563), .b(n_474), .o(n_571) );
BUF_X2 newInst_841 ( .a(newNet_840), .o(newNet_841) );
NAND2_Z01 cordic_Add0_Add_g660 ( .a(cordic_Add0_Add_n_45), .b(cordic_Add0_Add_n_13), .o(cordic_Add0_Add_n_47) );
BUF_X2 newInst_686 ( .a(newNet_685), .o(newNet_686) );
INV_X1 g13486 ( .a(n_798), .o(n_967) );
NAND2_Z01 g15426 ( .a(n_194), .b(n_96), .o(n_228) );
BUF_X2 newInst_1187 ( .a(newNet_231), .o(newNet_1187) );
NAND2_Z01 cordic_AddX_Add_g691 ( .a(cordic_AddX_Add_n_41), .b(cordic_AddX_Add_n_6), .o(cordic_AddX_Add_n_43) );
NAND2_Z01 g15070 ( .a(n_473), .b(PI_AD_3), .o(n_538) );
INV_Z1 cordic_Add0_g48 ( .a(cordic_Add0_Btemp_13_), .o(cordic_Add0_n_14) );
NAND2_Z01 cordic_Add0_MUX_0_g290 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_11_), .o(cordic_Add0_MUX_0_n_13) );
BUF_X2 newInst_747 ( .a(newNet_746), .o(newNet_747) );
NAND2_Z01 g15354 ( .a(n_214), .b(CoreOutputReg_15_), .o(n_307) );
BUF_X2 newInst_1088 ( .a(newNet_1087), .o(newNet_1088) );
INV_X2 newInst_986 ( .a(newNet_879), .o(newNet_986) );
NAND4_Z1 g14822 ( .a(n_279), .b(n_273), .c(n_690), .d(n_225), .o(n_697) );
AND2_X1 cordic_pla_g269 ( .a(cordic_tanangle_2_), .b(cordic_pla_n_10), .o(cordic_tanangle_0_) );
BUF_X2 newInst_780 ( .a(newNet_779), .o(newNet_780) );
NAND2_Z01 cordic_AddY_MUX_0_g318 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_13_), .o(cordic_AddY_MUX_0_n_3) );
BUF_X2 newInst_947 ( .a(newNet_946), .o(newNet_947) );
BUF_X2 newInst_867 ( .a(newNet_866), .o(newNet_867) );
BUF_X2 newInst_532 ( .a(newNet_403), .o(newNet_532) );
NAND2_Z01 cordic_SH2_srl_35_26_g1230 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_13_), .o(cordic_SH2_srl_35_26_n_22) );
XOR2_X1 cordic_Add0_Add_g682 ( .a(cordic_Add0_n_5), .b(cordic_Add0_Atemp_4_), .o(cordic_Add0_Add_n_25) );
NAND2_Z01 cordic_AddY_MUX_0_g273 ( .a(cordic_AddY_MUX_0_n_32), .b(cordic_AddY_MUX_0_n_7), .o(cordic_AddY_Atemp_15_) );
NAND2_Z01 cordic_AddY_Add_g682 ( .a(cordic_AddY_Add_n_50), .b(cordic_AddY_Add_n_0), .o(cordic_AddY_Add_n_52) );
NAND2_Z01 g15285 ( .a(n_274), .b(Access_Address_1_17_), .o(n_370) );
BUF_X2 newInst_125 ( .a(newNet_124), .o(newNet_125) );
XNOR2_X1 cordic_AddY_Compl_g376 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_7_), .o(cordic_AddY_Compl_n_6) );
AND2_X1 g46 ( .a(n_842), .b(n_856), .o(PO_AD_18) );
AND2_X1 g15635 ( .a(DevSel_Wait_Cnt_0_), .b(DevSel_Wait_Cnt_1_), .o(n_28) );
BUF_X2 newInst_135 ( .a(newNet_134), .o(newNet_135) );
NAND2_Z01 cordic_AddY_MUX_0_g320 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_10_), .o(cordic_AddY_MUX_0_n_1) );
NAND2_Z01 cordic_AddX_MUX_0_g309 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_0_), .o(cordic_AddX_MUX_0_n_12) );
NAND2_Z01 cordic_AddY_MUX_1_g294 ( .a(cordic_AddY_Y_1), .b(cordic_Y_1_), .o(cordic_AddY_MUX_1_n_27) );
NAND2_Z01 cordic_AddX_MUX_0_g293 ( .a(cordic_BS1_12_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_28) );
BUF_X2 newInst_64 ( .a(newNet_63), .o(newNet_64) );
NAND2_Z01 g13546 ( .a(n_712), .b(CoreOutputReg_1_), .o(n_740) );
XOR2_X1 g15161 ( .a(n_342), .b(n_343), .o(n_451) );
NAND2_Z01 cordic_Add0_MUX_1_g295 ( .a(cordic_tanangle_10_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_6) );
BUF_X2 newInst_1026 ( .a(newNet_1025), .o(newNet_1026) );
NAND2_Z01 cordic_g391 ( .a(cordic_n_75), .b(cordic_n_82), .o(cordic_n_116) );
NAND2_Z01 cordic_Add0_Add_g705 ( .a(cordic_Add0_n_2), .b(cordic_Add0_Atemp_1_), .o(cordic_Add0_Add_n_2) );
BUF_X2 newInst_353 ( .a(newNet_352), .o(newNet_353) );
NAND2_Z01 cordic_AddX_Add_g655 ( .a(cordic_AddX_Add_n_77), .b(cordic_AddX_Add_n_8), .o(cordic_AddX_Y_3) );
BUF_X2 newInst_604 ( .a(newNet_603), .o(newNet_604) );
INV_X2 newInst_328 ( .a(newNet_327), .o(newNet_328) );
INV_Z1 cordic_Add0_g56 ( .a(cordic_Add0_Btemp_5_), .o(cordic_Add0_n_6) );
BUF_X2 newInst_738 ( .a(newNet_591), .o(newNet_738) );
BUF_X2 newInst_288 ( .a(newNet_287), .o(newNet_288) );
NAND2_Z01 g15365 ( .a(n_214), .b(CoreOutputReg_1_), .o(n_296) );
BUF_X2 newInst_1087 ( .a(newNet_1086), .o(newNet_1087) );
NAND2_Z01 cordic_AddY_Add_g675 ( .a(cordic_AddY_Add_n_58), .b(cordic_AddY_Add_n_21), .o(cordic_AddY_Add_n_59) );
XOR2_X1 cordic_AddX_g200 ( .a(cordic_AddX_Btemp_8_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_8_) );
BUF_X2 newInst_979 ( .a(newNet_978), .o(newNet_979) );
NAND2_Z01 cordic_Add0_MUX_0_g269 ( .a(cordic_Add0_MUX_0_n_20), .b(cordic_Add0_MUX_0_n_9), .o(cordic_Add0_Atemp_3_) );
XOR2_X1 g15321 ( .a(n_159), .b(n_160), .o(n_339) );
BUF_X2 newInst_81 ( .a(newNet_34), .o(newNet_81) );
NAND2_Z01 cordic_Add0_MUX_0_g274 ( .a(cordic_tanangle_7_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_29) );
INV_X1 g15643 ( .a(PO_TRDY_L), .o(n_22) );
NAND2_Z01 g13489 ( .a(n_717), .b(n_760), .o(n_795) );
NAND2_Z01 cordic_AddX_Add_g684 ( .a(cordic_AddX_Add_n_49), .b(cordic_AddX_Add_n_28), .o(cordic_AddX_Add_n_50) );
BUF_X2 newInst_1100 ( .a(newNet_1099), .o(newNet_1100) );
BUF_X2 newInst_567 ( .a(newNet_566), .o(newNet_567) );
NAND4_Z1 g15222 ( .a(n_33), .b(n_1047), .c(n_203), .d(n_10), .o(n_432) );
BUF_X2 newInst_768 ( .a(newNet_91), .o(newNet_768) );
BUF_X2 newInst_670 ( .a(newNet_669), .o(newNet_670) );
BUF_X2 newInst_405 ( .a(newNet_404), .o(newNet_405) );
fflopd cordic_Y_reg_1_ ( .CK(newNet_72), .D(cordic_n_40), .Q(cordic_Y_1_) );
NAND2_Z01 g13472 ( .a(n_740), .b(n_777), .o(n_812) );
NAND2_Z01 g14900 ( .a(n_621), .b(n_550), .o(n_674) );
NAND2_Z01 cordic_SH2_srl_35_26_g1220 ( .a(cordic_iteration_0_), .b(cordic_X_8_), .o(cordic_SH2_srl_35_26_n_32) );
NAND2_Z01 cordic_AddY_Add_g734 ( .a(cordic_AddY_Btemp1_6_), .b(cordic_AddY_Atemp_6_), .o(cordic_AddY_Add_n_0) );
BUF_X2 newInst_50 ( .a(newNet_49), .o(newNet_50) );
NAND2_Z01 cordic_Add0_Compl_g365 ( .a(cordic_Add0_Compl_n_11), .b(cordic_Add0_Compl_n_1), .o(cordic_Add0_Compl_n_17) );
NAND2_Z01 cordic_g433 ( .a(cordic_SumAngle_10_), .b(cordic_n_7), .o(cordic_n_74) );
XOR2_X1 cordic_Add0_Add_g677 ( .a(cordic_Add0_n_7), .b(cordic_Add0_Atemp_6_), .o(cordic_Add0_Add_n_30) );
NAND2_Z01 g14899 ( .a(n_622), .b(n_551), .o(n_675) );
NAND2_Z01 g13524 ( .a(Idsel), .b(Config_Reg_17_), .o(n_762) );
BUF_X2 newInst_552 ( .a(newNet_551), .o(newNet_552) );
NAND3_Z1 g15153 ( .a(n_229), .b(n_371), .c(n_10), .o(n_459) );
AND2_X1 cordic_AddX_Compl_g351 ( .a(cordic_AddX_Compl_n_29), .b(cordic_AddX_Compl_n_10), .o(cordic_AddX_Compl_n_31) );
NAND3_Z1 cordic_SH2_srl_35_26_g1214 ( .a(cordic_SH2_srl_35_26_n_3), .b(cordic_SH2_srl_35_26_n_0), .c(cordic_X_15_), .o(cordic_SH2_srl_35_26_n_41) );
fflopd Config_Reg_reg_25_ ( .CK(newNet_936), .D(n_671), .Q(Config_Reg_25_) );
NOR2_Z1 cordic_g450 ( .a(cordic_n_9), .b(Issue_Rst), .o(cordic_n_57) );
NAND2_Z01 cordic_Add0_MUX_0_g258 ( .a(cordic_Add0_MUX_0_n_23), .b(cordic_Add0_MUX_0_n_5), .o(cordic_Add0_Atemp_12_) );
NAND2_Z01 g15247 ( .a(n_317), .b(n_318), .o(n_413) );
XNOR2_X1 cordic_AddY_Compl_g366 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_3_), .o(cordic_AddY_Compl_n_16) );
NAND2_Z01 cordic_g444 ( .a(cordic_SumAngle_6_), .b(cordic_n_7), .o(cordic_n_63) );
NAND2_Z01 cordic_AddY_MUX_0_g311 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_8_), .o(cordic_AddY_MUX_0_n_10) );
NAND2_Z01 g15241 ( .a(n_274), .b(Access_Address_1_29_), .o(n_419) );
NAND2_Z01 g14901 ( .a(n_620), .b(n_549), .o(n_673) );
NAND2_Z01 cordic_SH1_srl_35_26_g1166 ( .a(cordic_SH1_srl_35_26_n_56), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_86) );
NAND2_Z01 g15233 ( .a(n_274), .b(Access_Address_1_20_), .o(n_427) );
BUF_X2 newInst_121 ( .a(newNet_120), .o(newNet_121) );
INV_X2 cordic_SH1_srl_35_26_g1252 ( .a(cordic_iteration_0_), .o(cordic_SH1_srl_35_26_n_0) );
NAND3_Z1 g15107 ( .a(n_442), .b(n_443), .c(n_10), .o(n_501) );
NAND2_Z01 cordic_g449 ( .a(cordic_SumAngle_9_), .b(cordic_n_7), .o(cordic_n_58) );
BUF_X2 newInst_818 ( .a(newNet_817), .o(newNet_818) );
BUF_X2 newInst_654 ( .a(newNet_653), .o(newNet_654) );
NAND2_Z01 g13510 ( .a(Idsel), .b(Config_Reg_20_), .o(n_776) );
AND4_X1 g14946 ( .a(Access_Address_1_29_), .b(n_20), .c(n_561), .d(Access_Address_1_27_), .o(n_628) );
NAND2_Z01 g15514 ( .a(n_118), .b(First_Entry), .o(n_147) );
NAND2_Z01 g13535 ( .a(Idsel), .b(Config_Reg_23_), .o(n_751) );
NAND2_Z01 cordic_AddX_MUX_0_g315 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_11_), .o(cordic_AddX_MUX_0_n_6) );
NAND2_Z01 g15100 ( .a(n_473), .b(PI_AD_14), .o(n_508) );
INV_X1 g13465 ( .a(PAR_Int_d), .o(n_817) );
fflopd CBE_par_reg_2_ ( .CK(newNet_1078), .D(n_351), .Q(CBE_par_2_) );
NAND2_Z01 g13533 ( .a(Idsel), .b(Config_Reg_0_), .o(n_753) );
NAND2_Z01 cordic_g395 ( .a(cordic_n_70), .b(cordic_n_92), .o(cordic_n_112) );
BUF_X2 newInst_721 ( .a(newNet_720), .o(newNet_721) );
NAND2_Z01 cordic_AddX_MUX_0_g317 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_5_), .o(cordic_AddX_MUX_0_n_4) );
XOR2_X1 cordic_AddY_Compl_g346 ( .a(cordic_AddY_Compl_n_33), .b(cordic_AddY_Compl_n_9), .o(CoreOutput_10_) );
NAND2_Z01 cordic_AddX_Add_g721 ( .a(cordic_AddX_Btemp1_10_), .b(cordic_AddX_Atemp_10_), .o(cordic_AddX_Add_n_13) );
NAND2_Z01 cordic_SH2_srl_35_26_g1172 ( .a(cordic_SH2_srl_35_26_n_47), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_80) );
BUF_X2 newInst_999 ( .a(newNet_998), .o(newNet_999) );
BUF_X2 newInst_656 ( .a(newNet_27), .o(newNet_656) );
NOR2_Z1 g13440 ( .a(n_806), .b(n_710), .o(n_842) );
XOR2_X1 cordic_AddY_Add_g692 ( .a(cordic_AddY_Add_n_40), .b(cordic_AddY_Add_n_24), .o(cordic_AddY_Stemp_3_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1247 ( .a(cordic_SH1_srl_35_26_n_1), .b(cordic_iteration_2_), .o(cordic_SH1_srl_35_26_n_20) );
BUF_X2 newInst_179 ( .a(newNet_106), .o(newNet_179) );
NAND2_Z01 cordic_Add0_MUX_0_g284 ( .a(cordic_tanangle_2_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_19) );
fflopd CoreOutputReg_reg_3_ ( .CK(newNet_585), .D(n_379), .Q(CoreOutputReg_3_) );
NAND2_Z01 g14907 ( .a(n_614), .b(n_542), .o(n_667) );
AND2_X1 g15437 ( .a(n_185), .b(System_Busy), .o(n_271) );
NAND2_Z01 g15325 ( .a(n_213), .b(Trdy_Wait_Cnt_3_), .o(n_336) );
NAND2_Z01 cordic_SH2_srl_35_26_g1193 ( .a(cordic_SH2_srl_35_26_n_40), .b(cordic_SH2_srl_35_26_n_20), .o(cordic_SH2_srl_35_26_n_59) );
XOR2_X1 cordic_AddX_Add_g712 ( .a(cordic_AddX_Btemp1_14_), .b(cordic_AddX_Atemp_14_), .o(cordic_AddX_Add_n_22) );
INV_X2 newInst_939 ( .a(newNet_938), .o(newNet_939) );
BUF_X2 newInst_493 ( .a(newNet_492), .o(newNet_493) );
BUF_X2 newInst_749 ( .a(newNet_748), .o(newNet_749) );
NAND2_Z01 g15263 ( .a(n_284), .b(n_285), .o(n_397) );
INV_X2 newInst_704 ( .a(newNet_703), .o(newNet_704) );
fflopd CoreOutputReg_reg_1_ ( .CK(newNet_670), .D(n_402), .Q(CoreOutputReg_1_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1139 ( .a(cordic_SH2_srl_35_26_n_93), .b(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_113) );
NAND2_Z01 cordic_SH1_srl_35_26_g1216 ( .a(cordic_iteration_0_), .b(cordic_Y_13_), .o(cordic_SH1_srl_35_26_n_36) );
BUF_X2 newInst_272 ( .a(newNet_271), .o(newNet_272) );
NOR2_Z1 cordic_pla_g281 ( .a(cordic_pla_n_5), .b(cordic_pla_n_15), .o(cordic_tanangle_11_) );
NAND2_Z01 g14995 ( .a(n_572), .b(Config_Reg_13_), .o(n_582) );
XOR2_X1 g15486 ( .a(n_85), .b(n_86), .o(n_177) );
NAND2_Z01 g15340 ( .a(n_184), .b(PI_AD_25), .o(n_321) );
NAND2_Z01 g15376 ( .a(n_214), .b(CoreOutputReg_24_), .o(n_285) );
BUF_X2 newInst_201 ( .a(newNet_200), .o(newNet_201) );
INV_X1 cordic_g492 ( .a(CoreOutput_30_), .o(cordic_n_15) );
INV_X1 cordic_g489 ( .a(CoreOutput_27_), .o(cordic_n_18) );
NAND2_Z01 cordic_AddY_MUX_0_g283 ( .a(cordic_AddY_MUX_0_n_31), .b(cordic_AddY_MUX_0_n_9), .o(cordic_AddY_Atemp_14_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1108 ( .a(cordic_SH1_srl_35_26_n_128), .b(cordic_iteration_3_), .o(cordic_SH1_srl_35_26_n_144) );
BUF_X2 newInst_677 ( .a(newNet_676), .o(newNet_677) );
NAND2_Z01 g15296 ( .a(n_272), .b(PI_CBE_L_0), .o(n_359) );
BUF_X2 newInst_400 ( .a(newNet_282), .o(newNet_400) );
fflopd First_Entry_reg ( .CK(newNet_476), .D(n_693), .Q(First_Entry) );
BUF_X2 newInst_1009 ( .a(newNet_1008), .o(newNet_1009) );
NAND2_Z01 g13515 ( .a(Idsel), .b(Config_Reg_29_), .o(n_771) );
NOR2_Z1 cordic_SH2_srl_35_26_g1150 ( .a(cordic_SH2_srl_35_26_n_89), .b(cordic_iteration_3_), .o(cordic_BS2_14_) );
fflopd Config_Reg_reg_17_ ( .CK(newNet_995), .D(n_680), .Q(Config_Reg_17_) );
fflopd Config_Reg_reg_4_ ( .CK(newNet_885), .D(n_663), .Q(Config_Reg_4_) );
XOR2_X1 cordic_AddX_g212 ( .a(cordic_AddX_Btemp_1_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_1_) );
NAND2_Z01 cordic_AddY_Add_g670 ( .a(cordic_AddY_Add_n_62), .b(cordic_AddY_Add_n_13), .o(cordic_AddY_Add_n_64) );
BUF_X2 newInst_1041 ( .a(newNet_1040), .o(newNet_1041) );
NAND2_Z01 cordic_AddX_MUX_1_g276 ( .a(cordic_AddX_MUX_1_n_14), .b(cordic_AddX_MUX_1_n_29), .o(cordic_AddX_Btemp_2_) );
BUF_X2 newInst_256 ( .a(newNet_255), .o(newNet_256) );
INV_X1 cordic_g497 ( .a(CoreOutput_12_), .o(cordic_n_10) );
NAND2_Z01 cordic_AddY_Add_g687 ( .a(cordic_AddY_Add_n_46), .b(cordic_AddY_Add_n_31), .o(cordic_AddY_Add_n_47) );
fflopd Config_Reg_reg_26_ ( .CK(newNet_929), .D(n_670), .Q(Config_Reg_26_) );
BUF_X2 newInst_586 ( .a(newNet_521), .o(newNet_586) );
INV_X1 g15549 ( .a(n_112), .o(n_111) );
NAND2_Z01 cordic_SH2_srl_35_26_g1248 ( .a(cordic_SH2_srl_35_26_n_1), .b(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_19) );
NAND2_Z01 g13479 ( .a(n_723), .b(n_759), .o(n_805) );
NAND2_Z01 cordic_AddX_MUX_1_g311 ( .a(cordic_BS1_8_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_10) );
NAND2_Z01 g15122 ( .a(n_439), .b(n_93), .o(n_487) );
BUF_X2 newInst_500 ( .a(newNet_499), .o(newNet_500) );
XOR2_X1 g15493 ( .a(n_80), .b(n_67), .o(n_170) );
BUF_X2 newInst_1022 ( .a(newNet_1021), .o(newNet_1022) );
BUF_X2 newInst_607 ( .a(newNet_312), .o(newNet_607) );
NAND3_Z1 g15484 ( .a(n_43), .b(n_110), .c(n_10), .o(n_183) );
XOR2_X1 g15608 ( .a(PI_AD_52), .b(PI_AD_51), .o(n_57) );
BUF_X2 newInst_195 ( .a(newNet_194), .o(newNet_195) );
NAND2_Z01 g15358 ( .a(n_208), .b(n_138), .o(n_303) );
NAND2_Z01 g14925 ( .a(n_597), .b(n_526), .o(n_649) );
NAND2_Z01 g15051 ( .a(n_485), .b(Set_Data_Parity), .o(n_557) );
BUF_X2 newInst_557 ( .a(newNet_556), .o(newNet_557) );
XOR2_X1 cordic_AddY_Add_g710 ( .a(cordic_AddY_Btemp1_3_), .b(cordic_AddY_Atemp_3_), .o(cordic_AddY_Add_n_24) );
NAND2_Z01 cordic_SH1_srl_35_26_g1208 ( .a(cordic_SH1_srl_35_26_n_4), .b(cordic_SH1_srl_35_26_n_24), .o(cordic_SH1_srl_35_26_n_46) );
NAND2_Z01 cordic_AddX_MUX_1_g300 ( .a(cordic_AddX_Y_1), .b(cordic_X_5_), .o(cordic_AddX_MUX_1_n_21) );
BUF_X2 newInst_429 ( .a(newNet_428), .o(newNet_429) );
BUF_X2 newInst_990 ( .a(newNet_989), .o(newNet_990) );
BUF_X2 newInst_203 ( .a(newNet_132), .o(newNet_203) );
NAND2_Z01 cordic_SH1_srl_35_26_g1235 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_5_), .o(cordic_SH1_srl_35_26_n_14) );
NAND2_Z01 g15362 ( .a(CoreOutput_18_), .b(n_2), .o(n_299) );
BUF_X2 newInst_993 ( .a(newNet_992), .o(newNet_993) );
BUF_X2 newInst_921 ( .a(newNet_920), .o(newNet_921) );
BUF_X2 newInst_728 ( .a(newNet_727), .o(newNet_728) );
BUF_X2 newInst_1172 ( .a(newNet_891), .o(newNet_1172) );
XOR2_X1 g15001 ( .a(n_560), .b(n_166), .o(n_576) );
fflopd Config_Reg_reg_20_ ( .CK(newNet_980), .D(n_676), .Q(Config_Reg_20_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1238 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_12_), .o(cordic_SH1_srl_35_26_n_11) );
NOR2_Z1 g14839 ( .a(n_681), .b(n_231), .o(n_684) );
NOR2_Z1 cordic_pla_g289 ( .a(cordic_pla_n_5), .b(cordic_pla_n_12), .o(cordic_tanangle_12_) );
XOR2_X1 cordic_AddX_Compl_g358 ( .a(cordic_AddX_Compl_n_21), .b(cordic_AddX_Compl_n_7), .o(CoreOutput_21_) );
NAND2_Z01 g15552 ( .a(n_45), .b(First_Entry), .o(n_104) );
BUF_X2 newInst_155 ( .a(newNet_154), .o(newNet_155) );
BUF_X2 newInst_479 ( .a(newNet_478), .o(newNet_479) );
XOR2_X1 cordic_AddY_Add_g714 ( .a(cordic_AddY_Btemp1_2_), .b(cordic_AddY_Atemp_2_), .o(cordic_AddY_Add_n_20) );
XOR2_X1 cordic_Add0_Compl_g360 ( .a(cordic_Add0_Compl_n_19), .b(cordic_Add0_Compl_n_16), .o(cordic_SumAngle_3_) );
BUF_X2 newInst_1050 ( .a(newNet_1049), .o(newNet_1050) );
fflopd CoreOutputReg_reg_11_ ( .CK(newNet_719), .D(n_412), .Q(CoreOutputReg_11_) );
XOR2_X1 cordic_AddX_g205 ( .a(cordic_AddX_Btemp_5_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_5_) );
BUF_X2 newInst_1090 ( .a(newNet_866), .o(newNet_1090) );
NAND2_Z01 g14910 ( .a(n_610), .b(n_538), .o(n_664) );
BUF_X2 newInst_699 ( .a(newNet_698), .o(newNet_699) );
NAND2_Z01 cordic_SH2_srl_35_26_g1166 ( .a(cordic_SH2_srl_35_26_n_56), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_86) );
NAND2_Z01 g14950 ( .a(n_572), .b(Config_Reg_18_), .o(n_627) );
NAND2_Z01 cordic_SH2_srl_35_26_g1135 ( .a(cordic_SH2_srl_35_26_n_92), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_117) );
NAND2_Z01 g15389 ( .a(n_214), .b(CoreOutputReg_28_), .o(n_261) );
NAND2_Z01 cordic_Add0_MUX_0_g264 ( .a(cordic_Add0_MUX_0_n_27), .b(cordic_Add0_MUX_0_n_10), .o(cordic_Add0_Atemp_6_) );
BUF_X2 newInst_1161 ( .a(newNet_430), .o(newNet_1161) );
XOR2_X1 cordic_AddY_g204 ( .a(cordic_AddY_Btemp_6_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_6_) );
fflopd Trdy_Wait_Cnt_reg_2_ ( .CK(newNet_310), .D(n_366), .Q(Trdy_Wait_Cnt_2_) );
BUF_X2 newInst_859 ( .a(newNet_858), .o(newNet_859) );
BUF_X2 newInst_100 ( .a(newNet_6), .o(newNet_100) );
XOR2_X1 cordic_AddX_Add_g677 ( .a(cordic_AddX_Add_n_55), .b(cordic_AddX_Add_n_17), .o(cordic_AddX_Stemp_8_) );
BUF_X2 newInst_756 ( .a(newNet_755), .o(newNet_756) );
BUF_X2 newInst_523 ( .a(newNet_522), .o(newNet_523) );
fflopd CBE_par_reg_1_ ( .CK(newNet_1089), .D(n_350), .Q(CBE_par_1_) );
BUF_X2 newInst_890 ( .a(newNet_889), .o(newNet_890) );
NAND3_Z1 g15440 ( .a(Dual_Cycle), .b(n_139), .c(n_10), .o(n_219) );
BUF_X2 newInst_1000 ( .a(newNet_999), .o(newNet_1000) );
NAND2_Z01 cordic_SH2_srl_35_26_g1142 ( .a(cordic_SH2_srl_35_26_n_91), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_110) );
BUF_X2 newInst_683 ( .a(newNet_682), .o(newNet_683) );
XOR2_X1 g13395 ( .a(n_884), .b(PO_AD_20), .o(n_885) );
NAND2_Z01 cordic_SH1_srl_35_26_g1162 ( .a(cordic_SH1_srl_35_26_n_80), .b(cordic_SH1_srl_35_26_n_62), .o(cordic_SH1_srl_35_26_n_90) );
XOR2_X1 cordic_Add0_Compl_g358 ( .a(cordic_Add0_Compl_n_21), .b(cordic_Add0_Compl_n_7), .o(cordic_SumAngle_4_) );
BUF_X2 newInst_235 ( .a(newNet_55), .o(newNet_235) );
XOR2_X1 cordic_AddX_Compl_g354 ( .a(cordic_AddX_Compl_n_25), .b(cordic_AddX_Compl_n_4), .o(CoreOutput_23_) );
BUF_X2 newInst_600 ( .a(newNet_599), .o(newNet_600) );
NAND3_Z1 g15131 ( .a(n_328), .b(n_423), .c(n_10), .o(n_479) );
fflopd CoreOutputReg_reg_24_ ( .CK(newNet_635), .D(n_397), .Q(CoreOutputReg_24_) );
NAND2_Z01 cordic_AddY_MUX_1_g318 ( .a(cordic_BS2_13_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_3) );
BUF_X2 newInst_40 ( .a(newNet_28), .o(newNet_40) );
AND3_X1 g15573 ( .a(Trdy_Wait_Cnt_2_), .b(Trdy_Wait_Cnt_1_), .c(Trdy_Wait_Cnt_3_), .o(n_92) );
NOR2_Z1 g13433 ( .a(n_816), .b(n_710), .o(n_849) );
NAND2_Z01 cordic_AddX_Add_g664 ( .a(cordic_AddX_Add_n_68), .b(cordic_AddX_Add_n_4), .o(cordic_AddX_Add_n_70) );
NAND2_Z01 cordic_SH2_srl_35_26_g1187 ( .a(cordic_SH2_srl_35_26_n_54), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_65) );
BUF_X2 newInst_118 ( .a(newNet_13), .o(newNet_118) );
fflopd Config_Reg_reg_5_ ( .CK(newNet_874), .D(n_661), .Q(Config_Reg_5_) );
INV_Z1 cordic_AddX_MUX_0_g321 ( .a(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_0) );
NAND2_Z01 g14957 ( .a(n_572), .b(Config_Reg_23_), .o(n_620) );
BUF_X2 newInst_535 ( .a(newNet_486), .o(newNet_535) );
BUF_X2 newInst_342 ( .a(newNet_341), .o(newNet_342) );
NAND2_Z01 cordic_AddX_MUX_1_g308 ( .a(cordic_BS1_1_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_13) );
BUF_X2 newInst_783 ( .a(newNet_756), .o(newNet_783) );
BUF_X2 newInst_462 ( .a(newNet_461), .o(newNet_462) );
BUF_X2 newInst_279 ( .a(newNet_278), .o(newNet_279) );
BUF_X2 newInst_514 ( .a(newNet_513), .o(newNet_514) );
NAND2_Z01 g15346 ( .a(CoreOutput_11_), .b(n_2), .o(n_315) );
BUF_X2 newInst_189 ( .a(newNet_103), .o(newNet_189) );
NAND2_Z01 cordic_AddY_MUX_1_g291 ( .a(cordic_AddY_Y_1), .b(cordic_Y_9_), .o(cordic_AddY_MUX_1_n_30) );
NAND2_Z01 g15424 ( .a(n_184), .b(PI_AD_16), .o(n_229) );
XNOR2_X1 cordic_Add0_Compl_g377 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_5_), .o(cordic_Add0_Compl_n_5) );
XOR2_X1 g13411 ( .a(n_868), .b(PO_AD_11), .o(n_869) );
BUF_X2 newInst_507 ( .a(newNet_506), .o(newNet_507) );
BUF_X2 newInst_182 ( .a(newNet_181), .o(newNet_182) );
NOR2_Z4 g15146 ( .a(n_445), .b(n_132), .o(n_473) );
NAND3_Z1 g15314 ( .a(n_190), .b(n_212), .c(n_189), .o(n_381) );
BUF_X2 newInst_1082 ( .a(newNet_1081), .o(newNet_1082) );
NAND2_Z01 g15558 ( .a(n_34), .b(n_29), .o(n_101) );
BUF_X2 newInst_1095 ( .a(newNet_1094), .o(newNet_1095) );
INV_X1 drc_bufs15666 ( .a(n_184), .o(n_6) );
BUF_X2 newInst_633 ( .a(newNet_632), .o(newNet_633) );
NAND2_Z01 cordic_AddY_Add_g719 ( .a(cordic_AddY_Btemp1_7_), .b(cordic_AddY_Atemp_7_), .o(cordic_AddY_Add_n_15) );
NAND2_Z01 cordic_SH2_srl_35_26_g1237 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_9_), .o(cordic_SH2_srl_35_26_n_12) );
NOR4_Z1 g15543 ( .a(Trdy_Cnt_En), .b(System_Busy), .c(n_22), .d(RESET), .o(n_129) );
NAND2_Z01 cordic_SH1_srl_35_26_g1207 ( .a(cordic_SH1_srl_35_26_n_15), .b(cordic_SH1_srl_35_26_n_23), .o(cordic_SH1_srl_35_26_n_39) );
BUF_X2 newInst_499 ( .a(newNet_498), .o(newNet_499) );
INV_X1 g15548 ( .a(n_113), .o(n_114) );
BUF_X2 newInst_1121 ( .a(newNet_1120), .o(newNet_1121) );
BUF_X2 newInst_941 ( .a(newNet_940), .o(newNet_941) );
NAND2_Z01 cordic_AddY_MUX_0_g291 ( .a(cordic_BS2_9_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_30) );
NAND2_Z01 g15278 ( .a(n_324), .b(n_245), .o(n_377) );
BUF_X2 newInst_942 ( .a(newNet_941), .o(newNet_942) );
AND2_X1 cordic_Add0_Compl_g355 ( .a(cordic_Add0_Compl_n_25), .b(cordic_Add0_Compl_n_4), .o(cordic_Add0_Compl_n_27) );
NAND2_Z01 cordic_SH1_srl_35_26_g1188 ( .a(cordic_SH1_srl_35_26_n_44), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_64) );
NAND2_Z01 g15006 ( .a(n_565), .b(n_558), .o(n_573) );
XOR2_X1 cordic_AddX_Add_g698 ( .a(cordic_AddX_Add_n_34), .b(cordic_AddX_Add_n_18), .o(cordic_AddX_Stemp_1_) );
NAND3_Z1 g13422 ( .a(Check_Data_Parity), .b(n_1047), .c(n_10), .o(n_859) );
NAND2_Z01 cordic_AddX_MUX_1_g312 ( .a(cordic_BS1_14_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_9) );
AND2_X1 g15522 ( .a(n_106), .b(RESET), .o(n_155) );
XOR2_X1 cordic_AddX_Add_g683 ( .a(cordic_AddX_Add_n_49), .b(cordic_AddX_Add_n_28), .o(cordic_AddX_Stemp_6_) );
NAND2_Z01 g15369 ( .a(n_214), .b(CoreOutputReg_21_), .o(n_292) );
NAND2_Z01 g13494 ( .a(n_722), .b(n_756), .o(n_790) );
BUF_X2 newInst_428 ( .a(newNet_427), .o(newNet_428) );
BUF_X2 newInst_32 ( .a(newNet_31), .o(newNet_32) );
BUF_X2 newInst_1012 ( .a(newNet_1011), .o(newNet_1012) );
NAND2_Z01 g15253 ( .a(n_303), .b(n_205), .o(n_407) );
XOR2_X1 cordic_AddX_Compl_g362 ( .a(cordic_AddX_Compl_n_17), .b(cordic_AddX_Compl_n_14), .o(CoreOutput_19_) );
BUF_X2 newInst_79 ( .a(newNet_78), .o(newNet_79) );
NAND2_Z01 cordic_SH1_srl_35_26_g1107 ( .a(cordic_SH1_srl_35_26_n_130), .b(cordic_iteration_3_), .o(cordic_SH1_srl_35_26_n_145) );
NAND2_Z01 cordic_Add0_Add_g656 ( .a(cordic_Add0_Add_n_50), .b(cordic_Add0_Add_n_29), .o(cordic_Add0_Add_n_51) );
NAND2_Z01 cordic_SH1_srl_35_26_g1229 ( .a(cordic_iteration_0_), .b(cordic_Y_2_), .o(cordic_SH1_srl_35_26_n_23) );
NAND2_Z01 cordic_AddY_MUX_0_g298 ( .a(cordic_BS2_11_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_23) );
NAND2_Z01 cordic_AddY_MUX_0_g292 ( .a(cordic_BS2_2_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_29) );
NAND2_Z01 cordic_AddY_Add_g666 ( .a(cordic_AddY_Add_n_67), .b(cordic_AddY_Add_n_19), .o(cordic_AddY_Add_n_68) );
NAND2_Z01 cordic_SH2_srl_35_26_g1223 ( .a(cordic_iteration_0_), .b(cordic_X_3_), .o(cordic_SH2_srl_35_26_n_29) );
NAND2_Z01 g13569 ( .a(n_712), .b(CoreOutputReg_5_), .o(n_718) );
NAND2_Z01 cordic_AddX_MUX_0_g298 ( .a(cordic_BS1_11_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_23) );
NAND2_Z01 cordic_pla_g277 ( .a(cordic_pla_n_24), .b(cordic_pla_n_26), .o(cordic_tanangle_9_) );
BUF_X2 newInst_1045 ( .a(newNet_1044), .o(newNet_1045) );
fflopd cordic_X_reg_12_ ( .CK(newNet_45), .D(cordic_n_33), .Q(cordic_X_12_) );
BUF_X2 newInst_826 ( .a(newNet_825), .o(newNet_826) );
NAND2_Z01 cordic_SH2_srl_35_26_g1157 ( .a(cordic_SH2_srl_35_26_n_84), .b(cordic_SH2_srl_35_26_n_66), .o(cordic_SH2_srl_35_26_n_96) );
BUF_X2 newInst_60 ( .a(newNet_59), .o(newNet_60) );
NAND2_Z01 g15276 ( .a(n_248), .b(n_249), .o(n_379) );
NOR2_Z1 g15421 ( .a(n_207), .b(n_143), .o(n_231) );
XOR2_X1 cordic_Add0_Add_g664 ( .a(cordic_Add0_Add_n_41), .b(cordic_Add0_Add_n_25), .o(cordic_Add0_Stemp_4_) );
NAND2_Z01 g14986 ( .a(n_0), .b(CoreInput_5_), .o(n_591) );
BUF_X2 newInst_1078 ( .a(newNet_1077), .o(newNet_1078) );
INV_X1 g15613 ( .a(n_50), .o(n_49) );
INV_Z1 g8016 ( .a(Access_Type_1_3_), .o(n_897) );
NAND2_Z01 cordic_Add0_MUX_1_g294 ( .a(cordic_tanangle_5_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_7) );
XOR2_X1 g15592 ( .a(PI_AD_63), .b(PI_AD_32), .o(n_73) );
fflopd PO_DEVSEL_L_reg ( .CK(newNet_440), .D(n_704), .Q(PO_DEVSEL_L) );
fflopd Core_Cnt_reg_0_ ( .CK(newNet_549), .D(n_97), .Q(Core_Cnt_0_) );
BUF_X2 newInst_218 ( .a(newNet_140), .o(newNet_218) );
NAND3_Z1 g14816 ( .a(n_440), .b(n_694), .c(n_10), .o(n_703) );
AND2_X1 cordic_g476 ( .a(CoreOutput_24_), .b(Issue_Rst), .o(cordic_n_31) );
AND2_X1 g43 ( .a(n_848), .b(n_856), .o(PO_AD_21) );
XNOR2_X1 cordic_AddY_Compl_g367 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_9_), .o(cordic_AddY_Compl_n_15) );
XOR2_X1 cordic_AddX_Compl_g346 ( .a(cordic_AddX_Compl_n_33), .b(cordic_AddX_Compl_n_9), .o(CoreOutput_27_) );
NAND2_Z01 cordic_AddY_MUX_1_g302 ( .a(cordic_AddY_Y_1), .b(cordic_Y_10_), .o(cordic_AddY_MUX_1_n_19) );
BUF_X2 newInst_744 ( .a(newNet_80), .o(newNet_744) );
NAND2_Z01 g13552 ( .a(n_712), .b(CoreOutputReg_11_), .o(n_734) );
BUF_X2 newInst_26 ( .a(newNet_25), .o(newNet_26) );
NAND2_Z01 g15472 ( .a(n_135), .b(n_14), .o(n_190) );
NAND2_Z01 cordic_SH1_srl_35_26_g1122 ( .a(cordic_SH1_srl_35_26_n_113), .b(cordic_SH1_srl_35_26_n_88), .o(cordic_SH1_srl_35_26_n_130) );
NAND2_Z01 g15624 ( .a(n_25), .b(DevSel_Wait_Cnt_2_), .o(n_41) );
BUF_X2 newInst_619 ( .a(newNet_618), .o(newNet_619) );
fflopd CoreOutputReg_reg_13_ ( .CK(newNet_707), .D(n_410), .Q(CoreOutputReg_13_) );
BUF_X2 newInst_16 ( .a(newNet_15), .o(newNet_16) );
NAND4_Z1 g15538 ( .a(PI_CBE_L_3), .b(PI_CBE_L_0), .c(n_9), .d(PI_CBE_L_2), .o(n_133) );
NAND2_Z01 cordic_Add0_MUX_1_g281 ( .a(cordic_AngleCin), .b(cordic_Angle_9_), .o(cordic_Add0_MUX_1_n_20) );
NAND2_Z01 cordic_Add0_MUX_1_g276 ( .a(cordic_AngleCin), .b(cordic_Angle_10_), .o(cordic_Add0_MUX_1_n_25) );
NAND2_Z01 cordic_Add0_MUX_1_g257 ( .a(cordic_Add0_MUX_1_n_11), .b(cordic_Add0_MUX_1_n_32), .o(cordic_Add0_Btemp_11_) );
BUF_X2 newInst_441 ( .a(newNet_314), .o(newNet_441) );
BUF_X2 newInst_169 ( .a(newNet_168), .o(newNet_169) );
NAND2_Z01 g15332 ( .a(n_3), .b(PI_AD_23), .o(n_329) );
BUF_X2 newInst_1162 ( .a(newNet_1161), .o(newNet_1162) );
BUF_X2 newInst_549 ( .a(newNet_548), .o(newNet_549) );
NAND2_Z01 g15406 ( .a(n_214), .b(CoreOutputReg_6_), .o(n_244) );
BUF_X2 newInst_37 ( .a(newNet_36), .o(newNet_37) );
XOR2_X1 cordic_AddY_Compl_g342 ( .a(cordic_AddY_Compl_n_37), .b(cordic_AddY_Compl_n_12), .o(CoreOutput_12_) );
XOR2_X1 g15600 ( .a(PI_CBE_L_7), .b(PI_CBE_L_4), .o(n_65) );
NAND2_Z01 g15245 ( .a(n_274), .b(Access_Address_1_31_), .o(n_415) );
NAND2_Z01 cordic_SH1_srl_35_26_g1134 ( .a(cordic_SH1_srl_35_26_n_98), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_118) );
NAND2_Z01 cordic_AddX_MUX_0_g310 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_12_), .o(cordic_AddX_MUX_0_n_11) );
INV_X1 g15195 ( .a(n_445), .o(n_444) );
BUF_X2 newInst_613 ( .a(newNet_612), .o(newNet_613) );
NAND2_Z01 g15345 ( .a(n_214), .b(CoreOutputReg_11_), .o(n_316) );
XOR2_X1 cordic_AddX_Add_g695 ( .a(cordic_AddX_Add_n_37), .b(cordic_AddX_Add_n_20), .o(cordic_AddX_Stemp_2_) );
XOR2_X1 cordic_AddY_g200 ( .a(cordic_AddY_Btemp_8_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_8_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1243 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_4_), .o(cordic_SH1_srl_35_26_n_6) );
BUF_X2 newInst_207 ( .a(newNet_206), .o(newNet_207) );
NAND2_Z01 cordic_SH2_srl_35_26_g1184 ( .a(cordic_SH2_srl_35_26_n_43), .b(cordic_SH2_srl_35_26_n_55), .o(cordic_SH2_srl_35_26_n_68) );
NAND2_Z01 g14968 ( .a(n_572), .b(Config_Reg_4_), .o(n_609) );
BUF_X2 newInst_627 ( .a(newNet_626), .o(newNet_627) );
NAND3_Z1 g14840 ( .a(n_631), .b(n_567), .c(n_10), .o(n_683) );
NAND2_Z01 g15060 ( .a(n_473), .b(PI_AD_24), .o(n_548) );
AND2_X1 cordic_Add0_Compl_g353 ( .a(cordic_Add0_Compl_n_27), .b(cordic_Add0_Compl_n_6), .o(cordic_Add0_Compl_n_29) );
INV_X1 g15526 ( .a(n_131), .o(n_130) );
AND2_X1 g15565 ( .a(n_48), .b(Trdy_Wait_Cnt_0_), .o(n_96) );
BUF_X2 newInst_459 ( .a(newNet_458), .o(newNet_459) );
BUF_X2 newInst_649 ( .a(newNet_648), .o(newNet_649) );
NAND2_Z01 g15411 ( .a(CoreOutput_8_), .b(n_188), .o(n_239) );
XOR2_X1 g15585 ( .a(PI_AD_12), .b(PI_AD_6), .o(n_80) );
BUF_X2 newInst_918 ( .a(newNet_917), .o(newNet_918) );
XOR2_X1 g15492 ( .a(n_63), .b(n_78), .o(n_171) );
XOR2_X1 cordic_Add0_Add_g631 ( .a(cordic_Add0_Add_n_74), .b(cordic_Add0_Add_n_24), .o(cordic_Add0_Stemp_15_) );
BUF_X2 newInst_409 ( .a(newNet_408), .o(newNet_409) );
BUF_X2 newInst_364 ( .a(newNet_335), .o(newNet_364) );
BUF_X2 newInst_669 ( .a(newNet_668), .o(newNet_669) );
BUF_X2 newInst_864 ( .a(newNet_863), .o(newNet_864) );
INV_X1 g15381 ( .a(n_277), .o(n_278) );
NAND3_Z1 cordic_SH2_srl_35_26_g1163 ( .a(cordic_SH2_srl_35_26_n_3), .b(cordic_SH2_srl_35_26_n_46), .c(cordic_iteration_2_), .o(cordic_SH2_srl_35_26_n_88) );
NAND2_Z01 g15451 ( .a(n_156), .b(TAR_TRI_P), .o(n_204) );
BUF_X2 newInst_1145 ( .a(newNet_1144), .o(newNet_1145) );
INV_X1 g15382 ( .a(n_271), .o(n_270) );
NOR2_Z1 cordic_g430 ( .a(cordic_n_28), .b(Issue_Rst), .o(cordic_n_77) );
BUF_X2 newInst_955 ( .a(newNet_954), .o(newNet_955) );
NAND2_Z01 cordic_AddY_MUX_0_g314 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_15_), .o(cordic_AddY_MUX_0_n_7) );
INV_X1 cordic_g503 ( .a(CoreOutput_10_), .o(cordic_n_4) );
BUF_X2 newInst_520 ( .a(newNet_519), .o(newNet_520) );
NAND2_Z01 cordic_g411 ( .a(Issue_Rst), .b(CoreInput_11_), .o(cordic_n_96) );
NOR2_Z1 cordic_AddY_g67 ( .a(cordic_AngleCin), .b(cordic_Ysign), .o(cordic_AddY_n_1) );
NAND2_Z01 g14932 ( .a(n_589), .b(n_519), .o(n_642) );
BUF_X2 newInst_404 ( .a(newNet_403), .o(newNet_404) );
NAND2_Z01 g13542 ( .a(n_712), .b(CoreOutputReg_16_), .o(n_744) );
INV_X1 cordic_g486 ( .a(CoreOutput_3_), .o(cordic_n_21) );
BUF_X2 newInst_770 ( .a(newNet_769), .o(newNet_770) );
NAND2_Z01 cordic_AddY_Add_g723 ( .a(cordic_AddY_Btemp1_5_), .b(cordic_AddY_Atemp_5_), .o(cordic_AddY_Add_n_11) );
NAND2_Z01 g14972 ( .a(n_572), .b(Config_Reg_8_), .o(n_605) );
BUF_X2 newInst_966 ( .a(newNet_965), .o(newNet_966) );
BUF_X2 newInst_341 ( .a(newNet_132), .o(newNet_341) );
BUF_X2 newInst_291 ( .a(newNet_253), .o(newNet_291) );
NAND2_Z01 cordic_pla_g285 ( .a(cordic_pla_n_4), .b(cordic_pla_n_6), .o(cordic_pla_n_26) );
XOR2_X1 g15498 ( .a(n_105), .b(Core_Cnt_3_), .o(n_165) );
NAND2_Z01 g15259 ( .a(n_293), .b(n_294), .o(n_401) );
AND2_X1 cordic_AddX_Compl_g357 ( .a(cordic_AddX_Compl_n_23), .b(cordic_AddX_Compl_n_5), .o(cordic_AddX_Compl_n_25) );
BUF_X2 newInst_48 ( .a(newNet_47), .o(newNet_48) );
BUF_X2 newInst_660 ( .a(newNet_659), .o(newNet_660) );
NOR2_Z1 cordic_g456 ( .a(cordic_n_1), .b(Issue_Rst), .o(cordic_n_51) );
BUF_X2 newInst_817 ( .a(newNet_816), .o(newNet_817) );
BUF_X2 newInst_171 ( .a(newNet_170), .o(newNet_171) );
NAND2_Z01 cordic_SH1_srl_35_26_g1130 ( .a(cordic_SH1_srl_35_26_n_97), .b(cordic_SH1_srl_35_26_n_21), .o(cordic_SH1_srl_35_26_n_122) );
XOR2_X1 cordic_AddY_Add_g668 ( .a(cordic_AddY_Add_n_64), .b(cordic_AddY_Add_n_29), .o(cordic_AddY_Stemp_11_) );
NAND2_Z01 g13558 ( .a(n_712), .b(CoreOutputReg_18_), .o(n_729) );
NAND2_Z01 cordic_Add0_MUX_0_g283 ( .a(cordic_tanangle_3_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_20) );
XOR2_X1 cordic_AddX_Add_g708 ( .a(cordic_AddX_Btemp1_4_), .b(cordic_AddX_Atemp_4_), .o(cordic_AddX_Add_n_26) );
NAND2_Z01 g15622 ( .a(n_967), .b(n_10), .o(n_46) );
NAND2_Z01 cordic_Add0_Add_g693 ( .a(cordic_Add0_n_12), .b(cordic_Add0_Atemp_11_), .o(cordic_Add0_Add_n_14) );
BUF_X2 newInst_301 ( .a(newNet_122), .o(newNet_301) );
BUF_X2 newInst_55 ( .a(newNet_54), .o(newNet_55) );
NOR2_Z1 cordic_AddX_g67 ( .a(cordic_n_144), .b(cordic_Xsign), .o(cordic_AddX_n_1) );
BUF_X2 newInst_213 ( .a(newNet_96), .o(newNet_213) );
BUF_X2 newInst_6 ( .a(newNet_2), .o(newNet_6) );
NAND2_Z01 g14914 ( .a(n_607), .b(n_535), .o(n_660) );
fflopd CoreInput_reg_11_ ( .CK(newNet_815), .D(n_654), .Q(CoreInput_11_) );
NAND2_Z01 cordic_Add0_MUX_1_g263 ( .a(cordic_Add0_MUX_1_n_7), .b(cordic_Add0_MUX_1_n_24), .o(cordic_Add0_Btemp_5_) );
BUF_X2 newInst_623 ( .a(newNet_331), .o(newNet_623) );
BUF_X2 newInst_734 ( .a(newNet_733), .o(newNet_734) );
BUF_X2 newInst_581 ( .a(newNet_580), .o(newNet_581) );
NAND2_Z01 cordic_AddX_MUX_0_g274 ( .a(cordic_AddX_MUX_0_n_28), .b(cordic_AddX_MUX_0_n_11), .o(cordic_AddX_Atemp_12_) );
BUF_X2 newInst_267 ( .a(newNet_266), .o(newNet_267) );
NAND2_Z01 cordic_AddY_Add_g685 ( .a(cordic_AddY_Add_n_47), .b(cordic_AddY_Add_n_11), .o(cordic_AddY_Add_n_49) );
BUF_X2 newInst_606 ( .a(newNet_605), .o(newNet_606) );
NAND2_Z01 g13519 ( .a(Idsel), .b(Config_Reg_27_), .o(n_767) );
NAND3_Z1 cordic_SH1_srl_35_26_g1115 ( .a(cordic_SH1_srl_35_26_n_115), .b(cordic_SH1_srl_35_26_n_118), .c(cordic_SH1_srl_35_26_n_59), .o(cordic_BS1_7_) );
NAND2_Z01 cordic_pla_g299 ( .a(cordic_pla_n_3), .b(cordic_iteration_0_), .o(cordic_pla_n_12) );
XOR2_X1 g13401 ( .a(n_878), .b(PO_AD_6), .o(n_879) );
NAND2_Z01 cordic_AddX_MUX_0_g297 ( .a(cordic_BS1_7_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_24) );
NAND3_Z1 cordic_SH2_srl_35_26_g1117 ( .a(cordic_SH2_srl_35_26_n_110), .b(cordic_SH2_srl_35_26_n_111), .c(cordic_SH2_srl_35_26_n_109), .o(cordic_BS2_5_) );
AND2_X1 g348 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_46) );
XNOR2_X1 cordic_AddY_Compl_g375 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_4_), .o(cordic_AddY_Compl_n_7) );
BUF_X2 newInst_643 ( .a(newNet_642), .o(newNet_643) );
BUF_X2 newInst_452 ( .a(newNet_451), .o(newNet_452) );
BUF_X2 newInst_145 ( .a(newNet_144), .o(newNet_145) );
INV_X2 newInst_93 ( .a(newNet_92), .o(newNet_93) );
NAND2_Z01 g14915 ( .a(n_606), .b(n_546), .o(n_659) );
BUF_X2 newInst_347 ( .a(newNet_346), .o(newNet_347) );
XOR2_X1 cordic_AddY_g210 ( .a(cordic_AddY_Btemp_9_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_9_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1146 ( .a(cordic_SH2_srl_35_26_n_91), .b(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_106) );
BUF_X2 newInst_1132 ( .a(newNet_583), .o(newNet_1132) );
XOR2_X1 g15023 ( .a(n_449), .b(n_450), .o(n_559) );
fflopd System_Busy_reg ( .CK(newNet_371), .D(n_630), .Q(System_Busy) );
NAND2_Z01 cordic_SH2_srl_35_26_g1127 ( .a(cordic_SH2_srl_35_26_n_95), .b(cordic_iteration_2_), .o(cordic_SH2_srl_35_26_n_125) );
NAND2_Z01 cordic_AddY_MUX_1_g277 ( .a(cordic_AddY_MUX_1_n_10), .b(cordic_AddY_MUX_1_n_26), .o(cordic_AddY_Btemp_8_) );
AND2_X1 cordic_pla_g295 ( .a(cordic_pla_n_9), .b(cordic_iteration_0_), .o(cordic_pla_n_16) );
NAND2_Z01 cordic_AddY_Add_g678 ( .a(cordic_AddY_Add_n_55), .b(cordic_AddY_Add_n_17), .o(cordic_AddY_Add_n_56) );
INV_Z1 cordic_Add0_MUX_1_g299 ( .a(cordic_AngleCin), .o(cordic_Add0_MUX_1_n_2) );
fflopd TAR_TRI_E_reg ( .CK(newNet_362), .D(n_684), .Q(TAR_TRI_E) );
NAND2_Z01 g15433 ( .a(n_6), .b(n_155), .o(n_272) );
AND2_X1 cordic_Add0_Compl_g347 ( .a(cordic_Add0_Compl_n_33), .b(cordic_Add0_Compl_n_9), .o(cordic_Add0_Compl_n_35) );
BUF_X2 newInst_888 ( .a(newNet_887), .o(newNet_888) );
NOR2_Z1 cordic_SH2_srl_35_26_g1110 ( .a(cordic_SH2_srl_35_26_n_131), .b(cordic_iteration_3_), .o(cordic_BS2_10_) );
AND2_X1 g58 ( .a(n_821), .b(n_856), .o(PO_AD_6) );
NAND2_Z01 g15375 ( .a(CoreOutput_23_), .b(n_188), .o(n_286) );
NAND2_Z01 g15085 ( .a(n_494), .b(PI_AD_3), .o(n_523) );
NAND2_Z01 cordic_AddX_Add_g673 ( .a(cordic_AddX_Add_n_59), .b(cordic_AddX_Add_n_5), .o(cordic_AddX_Add_n_61) );
BUF_X2 newInst_732 ( .a(newNet_731), .o(newNet_732) );
BUF_X1 drc_bufs15692 ( .a(n_571), .o(n_0) );
BUF_X2 newInst_1030 ( .a(newNet_1029), .o(newNet_1030) );
BUF_X2 newInst_853 ( .a(newNet_852), .o(newNet_853) );
NAND2_Z01 g15286 ( .a(n_274), .b(Access_Address_1_18_), .o(n_369) );
NAND2_Z01 g14936 ( .a(n_584), .b(n_512), .o(n_638) );
NAND2_Z01 g15101 ( .a(n_473), .b(PI_AD_15), .o(n_507) );
NAND3_Z1 g15157 ( .a(n_137), .b(n_386), .c(DWord_Trans), .o(n_455) );
XNOR2_X1 g15578 ( .a(Core_Cnt_0_), .b(Core_Cnt_1_), .o(n_87) );
BUF_X2 newInst_435 ( .a(newNet_434), .o(newNet_435) );
NOR2_Z1 cordic_SH2_srl_35_26_g1114 ( .a(cordic_SH2_srl_35_26_n_127), .b(cordic_iteration_3_), .o(cordic_BS2_11_) );
BUF_X2 newInst_833 ( .a(newNet_832), .o(newNet_833) );
BUF_X2 newInst_465 ( .a(newNet_464), .o(newNet_465) );
BUF_X2 newInst_70 ( .a(newNet_69), .o(newNet_70) );
NAND2_Z01 cordic_SH2_srl_35_26_g1180 ( .a(cordic_SH2_srl_35_26_n_42), .b(cordic_SH2_srl_35_26_n_49), .o(cordic_SH2_srl_35_26_n_72) );
NAND2_Z01 cordic_SH2_srl_35_26_g1177 ( .a(cordic_SH2_srl_35_26_n_51), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_75) );
NAND2_Z01 g13532 ( .a(Idsel), .b(Config_Reg_24_), .o(n_754) );
NAND2_Z01 cordic_Add0_Add_g695 ( .a(cordic_Add0_n_14), .b(cordic_Add0_Atemp_13_), .o(cordic_Add0_Add_n_12) );
fflopd Config_Reg_reg_18_ ( .CK(newNet_986), .D(n_679), .Q(Config_Reg_18_) );
BUF_X2 newInst_1152 ( .a(newNet_145), .o(newNet_1152) );
NAND4_Z1 g15216 ( .a(Access_Address_1_22_), .b(Access_Address_1_23_), .c(n_180), .d(Access_Address_1_21_), .o(n_437) );
XOR2_X1 g15595 ( .a(PI_AD_27), .b(PI_AD_15), .o(n_70) );
NAND2_Z01 cordic_AddY_Add_g663 ( .a(cordic_AddY_Add_n_70), .b(cordic_AddY_Add_n_23), .o(cordic_AddY_Add_n_71) );
BUF_X2 newInst_247 ( .a(newNet_246), .o(newNet_247) );
NOR2_Z1 g13456 ( .a(n_789), .b(n_710), .o(n_826) );
INV_X1 cordic_g498 ( .a(CoreOutput_5_), .o(cordic_n_9) );
NAND2_Z01 g15138 ( .a(n_444), .b(n_35), .o(n_474) );
NAND2_Z01 cordic_Add0_MUX_0_g277 ( .a(cordic_tanangle_10_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_26) );
fflopd Config_Reg_reg_30_ ( .CK(newNet_894), .D(n_665), .Q(Config_Reg_30_) );
INV_X1 cordic_g481 ( .a(CoreOutput_15_), .o(cordic_n_26) );
NAND2_Z01 cordic_SH2_srl_35_26_g1228 ( .a(cordic_iteration_0_), .b(cordic_X_15_), .o(cordic_SH2_srl_35_26_n_24) );
NAND2_Z01 g15344 ( .a(CoreOutput_10_), .b(n_188), .o(n_317) );
NAND2_Z01 cordic_SH1_srl_35_26_g1222 ( .a(cordic_iteration_0_), .b(cordic_Y_5_), .o(cordic_SH1_srl_35_26_n_30) );
NAND2_Z01 g15366 ( .a(CoreOutput_1_), .b(n_188), .o(n_295) );
NAND3_Z1 cordic_SH1_srl_35_26_g1212 ( .a(cordic_iteration_1_), .b(cordic_SH1_srl_35_26_n_0), .c(cordic_Y_15_), .o(cordic_SH1_srl_35_26_n_38) );
fflopd Config_Reg_reg_29_ ( .CK(newNet_909), .D(n_667), .Q(Config_Reg_29_) );
NAND3_Z1 g13503 ( .a(State_0_), .b(n_898), .c(State_1_), .o(n_798) );
NAND2_Z01 g15097 ( .a(n_473), .b(PI_AD_12), .o(n_511) );
BUF_X2 newInst_11 ( .a(newNet_10), .o(newNet_11) );
NAND2_Z01 g13539 ( .a(n_712), .b(CoreOutputReg_30_), .o(n_747) );
BUF_X2 newInst_1037 ( .a(newNet_1036), .o(newNet_1037) );
INV_X1 cordic_Add0_MUX_1_g301 ( .a(cordic_Angle_15_), .o(cordic_Add0_MUX_1_n_0) );
XOR2_X1 cordic_AddX_Add_g680 ( .a(cordic_AddX_Add_n_52), .b(cordic_AddX_Add_n_30), .o(cordic_AddX_Stemp_7_) );
NAND2_Z01 g15513 ( .a(n_108), .b(n_51), .o(n_148) );
NAND2_Z01 cordic_SH1_srl_35_26_g1219 ( .a(cordic_iteration_0_), .b(cordic_Y_12_), .o(cordic_SH1_srl_35_26_n_33) );
BUF_X2 newInst_712 ( .a(newNet_711), .o(newNet_712) );
INV_X2 newInst_751 ( .a(newNet_750), .o(newNet_751) );
XNOR2_X1 cordic_Add0_Compl_g374 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_13_), .o(cordic_Add0_Compl_n_8) );
NAND2_Z01 g14991 ( .a(n_572), .b(Config_Reg_0_), .o(n_586) );
AND2_X1 g35 ( .a(n_843), .b(n_856), .o(PO_AD_29) );
NAND2_Z01 cordic_SH2_srl_35_26_g1238 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_12_), .o(cordic_SH2_srl_35_26_n_11) );
NAND2_Z01 cordic_AddY_MUX_1_g284 ( .a(cordic_AddY_MUX_1_n_3), .b(cordic_AddY_MUX_1_n_20), .o(cordic_AddY_Btemp_13_) );
NAND2_Z01 g14835 ( .a(n_685), .b(n_130), .o(n_686) );
NAND2_Z01 g15629 ( .a(Access_Type_1_2_), .b(Access_Type_1_3_), .o(n_30) );
BUF_X2 newInst_972 ( .a(newNet_971), .o(newNet_972) );
BUF_X2 newInst_1110 ( .a(newNet_1109), .o(newNet_1110) );
BUF_X2 newInst_970 ( .a(newNet_969), .o(newNet_970) );
AND2_X1 g15636 ( .a(Check_Add_Parity), .b(Check_Attr_Parity), .o(n_33) );
NAND2_Z01 g15295 ( .a(n_276), .b(n_126), .o(n_360) );
NOR2_Z1 g15435 ( .a(n_179), .b(n_116), .o(n_223) );
NOR2_Z1 g13437 ( .a(n_811), .b(n_710), .o(n_845) );
fflopd cordic_Angle_reg_2_ ( .CK(newNet_238), .D(cordic_n_109), .Q(cordic_Angle_2_) );
NAND2_Z01 cordic_AddX_MUX_1_g284 ( .a(cordic_AddX_MUX_1_n_3), .b(cordic_AddX_MUX_1_n_20), .o(cordic_AddX_Btemp_13_) );
BUF_X2 newInst_932 ( .a(newNet_931), .o(newNet_932) );
XOR2_X1 cordic_AddY_Compl_g362 ( .a(cordic_AddY_Compl_n_17), .b(cordic_AddY_Compl_n_14), .o(CoreOutput_2_) );
BUF_X2 newInst_1117 ( .a(newNet_1116), .o(newNet_1117) );
NAND2_Z01 cordic_AddY_MUX_1_g317 ( .a(cordic_BS2_5_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_4) );
NAND2_Z01 g15618 ( .a(n_12), .b(Trdy_Wait_Cnt_3_), .o(n_42) );
AND2_X1 cordic_AddX_Compl_g347 ( .a(cordic_AddX_Compl_n_33), .b(cordic_AddX_Compl_n_9), .o(cordic_AddX_Compl_n_35) );
BUF_X2 newInst_961 ( .a(newNet_960), .o(newNet_961) );
NAND2_Z01 cordic_AddY_MUX_1_g278 ( .a(cordic_AddY_MUX_1_n_13), .b(cordic_AddY_MUX_1_n_27), .o(cordic_AddY_Btemp_1_) );
NOR2_Z1 g13452 ( .a(n_800), .b(n_710), .o(n_830) );
BUF_X2 newInst_695 ( .a(newNet_694), .o(newNet_695) );
INV_X1 g15443 ( .a(n_216), .o(n_215) );
fflopd cordic_Y_reg_12_ ( .CK(newNet_86), .D(cordic_n_44), .Q(cordic_Y_12_) );
XOR2_X1 cordic_Add0_Add_g683 ( .a(cordic_Add0_n_16), .b(cordic_Add0_Atemp_15_), .o(cordic_Add0_Add_n_24) );
BUF_X2 newInst_831 ( .a(newNet_830), .o(newNet_831) );
BUF_X2 newInst_894 ( .a(newNet_71), .o(newNet_894) );
NAND2_Z01 g15518 ( .a(n_101), .b(Access_Type_1_3_), .o(n_144) );
XOR2_X1 g3 ( .a(n_892), .b(PO_AD_31), .o(n_1062) );
NAND2_Z01 cordic_AddY_MUX_0_g287 ( .a(cordic_AddY_MUX_0_n_18), .b(cordic_AddY_MUX_0_n_2), .o(cordic_AddY_Atemp_4_) );
XOR2_X1 g15318 ( .a(n_171), .b(n_172), .o(n_342) );
BUF_X2 newInst_158 ( .a(newNet_157), .o(newNet_158) );
NOR2_Z1 g13449 ( .a(n_793), .b(n_710), .o(n_833) );
BUF_X2 newInst_90 ( .a(newNet_67), .o(newNet_90) );
BUF_X2 newInst_687 ( .a(newNet_686), .o(newNet_687) );
AND2_X1 g62 ( .a(n_847), .b(n_856), .o(PO_AD_2) );
BUF_X2 newInst_357 ( .a(newNet_356), .o(newNet_357) );
NAND2_Z01 cordic_Add0_Add_g702 ( .a(cordic_Add0_n_10), .b(cordic_Add0_Atemp_9_), .o(cordic_Add0_Add_n_5) );
NAND2_Z01 g15065 ( .a(n_473), .b(PI_AD_28), .o(n_543) );
NAND2_Z01 g15104 ( .a(n_494), .b(PI_AD_16), .o(n_504) );
NAND2_Z01 cordic_SH2_srl_35_26_g1131 ( .a(cordic_SH2_srl_35_26_n_99), .b(cordic_SH2_srl_35_26_n_2), .o(cordic_SH2_srl_35_26_n_121) );
AND2_X1 cordic_Add0_Compl_g341 ( .a(cordic_Add0_Compl_n_39), .b(cordic_Add0_Compl_n_8), .o(cordic_Add0_Compl_n_41) );
fflopd cordic_X_reg_10_ ( .CK(newNet_172), .D(cordic_n_59), .Q(cordic_X_10_) );
BUF_X2 newInst_1176 ( .a(newNet_1175), .o(newNet_1176) );
NAND2_Z01 cordic_SH2_srl_35_26_g1196 ( .a(cordic_SH2_srl_35_26_n_12), .b(cordic_SH2_srl_35_26_n_37), .o(cordic_SH2_srl_35_26_n_56) );
NAND2_Z01 g15269 ( .a(n_257), .b(n_256), .o(n_391) );
XOR2_X1 cordic_AddY_Compl_g337 ( .a(cordic_AddY_Compl_n_43), .b(cordic_AddY_Compl_n_2), .o(CoreOutput_15_) );
BUF_X2 newInst_1186 ( .a(newNet_223), .o(newNet_1186) );
INV_X2 drc_bufs15677 ( .a(n_1), .o(n_2) );
BUF_X2 newInst_229 ( .a(newNet_157), .o(newNet_229) );
BUF_X2 newInst_983 ( .a(newNet_982), .o(newNet_983) );
NOR2_Z1 cordic_g459 ( .a(cordic_n_19), .b(Issue_Rst), .o(cordic_n_48) );
BUF_X2 newInst_192 ( .a(newNet_191), .o(newNet_192) );
fflopd PAR64_Int_reg ( .CK(newNet_454), .D(n_682), .Q(PAR64_Int) );
fflopd CoreOutputReg_reg_16_ ( .CK(newNet_693), .D(n_406), .Q(CoreOutputReg_16_) );
BUF_X2 newInst_511 ( .a(newNet_510), .o(newNet_511) );
BUF_X2 newInst_352 ( .a(newNet_79), .o(newNet_352) );
BUF_X2 newInst_1028 ( .a(newNet_1027), .o(newNet_1028) );
NAND2_Z01 cordic_SH1_srl_35_26_g1157 ( .a(cordic_SH1_srl_35_26_n_84), .b(cordic_SH1_srl_35_26_n_66), .o(cordic_SH1_srl_35_26_n_96) );
BUF_X2 newInst_1104 ( .a(newNet_1103), .o(newNet_1104) );
NOR2_Z1 cordic_g451 ( .a(cordic_n_15), .b(Issue_Rst), .o(cordic_n_56) );
XOR2_X1 cordic_Add0_Add_g643 ( .a(cordic_Add0_Add_n_62), .b(cordic_Add0_Add_n_31), .o(cordic_Add0_Stemp_11_) );
BUF_X2 newInst_625 ( .a(newNet_624), .o(newNet_625) );
NAND2_Z01 g15074 ( .a(n_473), .b(PI_AD_8), .o(n_534) );
NAND2_Z01 cordic_AddX_MUX_1_g301 ( .a(cordic_AddX_Y_1), .b(cordic_X_13_), .o(cordic_AddX_MUX_1_n_20) );
NAND2_Z01 cordic_AddX_MUX_1_g304 ( .a(cordic_AddX_Y_1), .b(cordic_X_3_), .o(cordic_AddX_MUX_1_n_17) );
BUF_X2 newInst_251 ( .a(newNet_250), .o(newNet_251) );
NAND2_Z01 cordic_Add0_MUX_1_g286 ( .a(cordic_tanangle_8_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_15) );
NAND2_Z01 cordic_AddX_MUX_1_g315 ( .a(cordic_BS1_11_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_6) );
BUF_X2 newInst_708 ( .a(newNet_332), .o(newNet_708) );
BUF_X2 newInst_194 ( .a(newNet_193), .o(newNet_194) );
BUF_X2 newInst_389 ( .a(newNet_388), .o(newNet_389) );
NAND2_Z01 g14975 ( .a(n_0), .b(CoreInput_10_), .o(n_602) );
BUF_X2 newInst_653 ( .a(newNet_652), .o(newNet_653) );
BUF_X2 newInst_310 ( .a(newNet_309), .o(newNet_310) );
fflopd Issue_Rst_reg ( .CK(newNet_460), .D(n_569), .Q(Issue_Rst) );
NAND2_Z01 g14963 ( .a(n_572), .b(Config_Reg_29_), .o(n_614) );
BUF_X2 newInst_931 ( .a(newNet_930), .o(newNet_931) );
BUF_X2 newInst_393 ( .a(newNet_392), .o(newNet_393) );
NAND2_Z01 cordic_SH1_srl_35_26_g1179 ( .a(cordic_SH1_srl_35_26_n_42), .b(cordic_SH1_srl_35_26_n_39), .o(cordic_SH1_srl_35_26_n_73) );
BUF_X2 newInst_115 ( .a(newNet_114), .o(newNet_115) );
NAND2_Z01 cordic_SH1_srl_35_26_g1186 ( .a(cordic_SH1_srl_35_26_n_47), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_66) );
BUF_X2 newInst_531 ( .a(newNet_530), .o(newNet_531) );
BUF_X2 newInst_1109 ( .a(newNet_1108), .o(newNet_1109) );
NAND2_Z01 g14894 ( .a(n_626), .b(n_556), .o(n_680) );
NAND2_Z01 g14979 ( .a(n_571), .b(CoreInput_14_), .o(n_598) );
NOR2_Z1 g13457 ( .a(n_788), .b(n_710), .o(n_825) );
BUF_X2 newInst_790 ( .a(newNet_789), .o(newNet_790) );
NAND2_Z01 g14921 ( .a(n_600), .b(n_530), .o(n_653) );
XNOR2_X1 cordic_Add0_Compl_g369 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_14_), .o(cordic_Add0_Compl_n_13) );
NAND2_Z01 cordic_Add0_MUX_0_g270 ( .a(cordic_Add0_MUX_0_n_19), .b(cordic_Add0_MUX_0_n_18), .o(cordic_Add0_Atemp_2_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1112 ( .a(cordic_SH1_srl_35_26_n_129), .b(cordic_iteration_3_), .o(cordic_BS1_9_) );
NOR2_Z1 cordic_g466 ( .a(cordic_n_26), .b(Issue_Rst), .o(cordic_n_41) );
NAND2_Z01 g15372 ( .a(n_214), .b(CoreOutputReg_22_), .o(n_289) );
BUF_X2 newInst_1139 ( .a(newNet_1138), .o(newNet_1139) );
XNOR2_X1 cordic_Add0_Compl_g372 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_8_), .o(cordic_Add0_Compl_n_10) );
NAND2_Z01 cordic_SH2_srl_35_26_g1243 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_4_), .o(cordic_SH2_srl_35_26_n_6) );
NAND2_Z01 cordic_SH1_srl_35_26_g1184 ( .a(cordic_SH1_srl_35_26_n_43), .b(cordic_SH1_srl_35_26_n_55), .o(cordic_SH1_srl_35_26_n_68) );
BUF_X2 newInst_928 ( .a(newNet_927), .o(newNet_928) );
BUF_X2 newInst_1066 ( .a(newNet_116), .o(newNet_1066) );
BUF_X2 newInst_475 ( .a(newNet_474), .o(newNet_475) );
NOR2_Z1 g15307 ( .a(n_223), .b(RESET), .o(n_386) );
XOR2_X1 g15588 ( .a(PI_AD_11), .b(PI_AD_5), .o(n_77) );
NAND2_Z01 cordic_AddY_MUX_1_g295 ( .a(cordic_AddY_Y_1), .b(cordic_Y_8_), .o(cordic_AddY_MUX_1_n_26) );
XOR2_X1 cordic_AddY_Add_g695 ( .a(cordic_AddY_Add_n_37), .b(cordic_AddY_Add_n_20), .o(cordic_AddY_Stemp_2_) );
XOR2_X1 g15604 ( .a(PI_AD_62), .b(PI_AD_33), .o(n_61) );
NAND2_Z01 cordic_g396 ( .a(cordic_n_69), .b(cordic_n_91), .o(cordic_n_111) );
NAND2_Z01 cordic_g416 ( .a(Issue_Rst), .b(CoreInput_16_), .o(cordic_n_91) );
BUF_X2 newInst_239 ( .a(newNet_168), .o(newNet_239) );
NAND2_Z01 cordic_g423 ( .a(Issue_Rst), .b(CoreInput_8_), .o(cordic_n_84) );
NAND2_Z01 cordic_g403 ( .a(cordic_n_62), .b(cordic_n_84), .o(cordic_n_104) );
BUF_X2 newInst_372 ( .a(newNet_200), .o(newNet_372) );
BUF_X2 newInst_275 ( .a(newNet_274), .o(newNet_275) );
NAND2_Z01 cordic_AddY_MUX_1_g283 ( .a(cordic_AddY_MUX_1_n_9), .b(cordic_AddY_MUX_1_n_31), .o(cordic_AddY_Btemp_14_) );
XOR2_X1 g15575 ( .a(PI_CBE_L_2), .b(PI_CBE_L_1), .o(n_90) );
NAND2_Z01 cordic_AddX_Add_g724 ( .a(cordic_AddX_Btemp1_14_), .b(cordic_AddX_Atemp_14_), .o(cordic_AddX_Add_n_10) );
INV_X1 cordic_SH1_srl_35_26_g1231 ( .a(cordic_SH1_srl_35_26_n_19), .o(cordic_SH1_srl_35_26_n_18) );
NAND2_Z01 g15336 ( .a(n_214), .b(CoreOutputReg_9_), .o(n_325) );
NAND2_Z01 cordic_AddX_MUX_1_g297 ( .a(cordic_AddX_Y_1), .b(cordic_X_7_), .o(cordic_AddX_MUX_1_n_24) );
fflopd Par64_Sgnl_reg ( .CK(newNet_406), .D(n_562), .Q(Par64_Sgnl) );
NAND2_Z01 cordic_Add0_MUX_0_g259 ( .a(cordic_Add0_MUX_0_n_32), .b(cordic_Add0_MUX_0_n_13), .o(cordic_Add0_Atemp_11_) );
BUF_X2 newInst_471 ( .a(newNet_470), .o(newNet_471) );
XOR2_X1 g13410 ( .a(n_869), .b(PO_AD_5), .o(n_870) );
BUF_X2 newInst_346 ( .a(newNet_345), .o(newNet_346) );
NAND2_Z01 cordic_Add0_MUX_0_g286 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_8_), .o(cordic_Add0_MUX_0_n_17) );
NAND2_Z01 cordic_SH1_srl_35_26_g1195 ( .a(cordic_SH1_srl_35_26_n_10), .b(cordic_SH1_srl_35_26_n_33), .o(cordic_SH1_srl_35_26_n_57) );
BUF_X2 newInst_529 ( .a(newNet_528), .o(newNet_529) );
BUF_X2 newInst_325 ( .a(newNet_324), .o(newNet_325) );
INV_X1 g15524 ( .a(n_139), .o(n_138) );
BUF_X2 newInst_571 ( .a(newNet_570), .o(newNet_571) );
NAND2_Z01 cordic_SH2_srl_35_26_g1169 ( .a(cordic_SH2_srl_35_26_n_44), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_83) );
NAND2_Z01 g14920 ( .a(n_601), .b(n_531), .o(n_654) );
NAND2_Z01 g15329 ( .a(n_184), .b(PI_AD_30), .o(n_332) );
NAND2_Z01 cordic_SH1_srl_35_26_g1234 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_1_), .o(cordic_SH1_srl_35_26_n_15) );
XNOR2_X1 cordic_AddX_Compl_g373 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_10_), .o(cordic_AddX_Compl_n_9) );
XOR2_X1 g13415 ( .a(n_864), .b(PO_AD_15), .o(n_865) );
XNOR2_X1 cordic_AddY_Compl_g380 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_11_), .o(cordic_AddY_Compl_n_3) );
NAND2_Z01 g13474 ( .a(n_739), .b(n_776), .o(n_810) );
AND2_X1 g53 ( .a(n_839), .b(n_856), .o(PO_AD_11) );
INV_X1 g15645 ( .a(Access_Address_1_28_), .o(n_20) );
BUF_X2 newInst_392 ( .a(newNet_391), .o(newNet_392) );
BUF_X2 newInst_412 ( .a(newNet_411), .o(newNet_412) );
BUF_X2 newInst_1055 ( .a(newNet_1054), .o(newNet_1055) );
BUF_X2 newInst_199 ( .a(newNet_5), .o(newNet_199) );
BUF_X2 newInst_483 ( .a(newNet_482), .o(newNet_483) );
BUF_X2 newInst_44 ( .a(newNet_43), .o(newNet_44) );
XOR2_X1 cordic_AddY_g207 ( .a(cordic_AddY_Btemp_10_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_10_) );
XOR2_X1 cordic_AddY_Add_g707 ( .a(cordic_AddY_Btemp1_10_), .b(cordic_AddY_Atemp_10_), .o(cordic_AddY_Add_n_27) );
NAND2_Z01 g14944 ( .a(n_577), .b(n_7), .o(n_630) );
AND2_X1 g64 ( .a(n_824), .b(n_856), .o(PO_AD_0) );
NOR2_Z1 g13444 ( .a(n_797), .b(n_710), .o(n_838) );
BUF_X2 newInst_797 ( .a(newNet_796), .o(newNet_797) );
BUF_X2 newInst_299 ( .a(newNet_298), .o(newNet_299) );
XOR2_X1 g15609 ( .a(PI_AD_61), .b(PI_AD_35), .o(n_56) );
NAND2_Z01 cordic_Add0_MUX_0_g268 ( .a(cordic_Add0_MUX_0_n_31), .b(cordic_Add0_MUX_0_n_17), .o(cordic_Add0_Atemp_8_) );
BUF_X2 newInst_871 ( .a(newNet_870), .o(newNet_871) );
BUF_X2 newInst_850 ( .a(newNet_849), .o(newNet_850) );
NAND2_Z01 g15401 ( .a(n_214), .b(CoreOutputReg_3_), .o(n_249) );
NAND2_Z01 g14953 ( .a(n_572), .b(Config_Reg_1_), .o(n_624) );
NAND2_Z01 g15081 ( .a(n_494), .b(PI_AD_14), .o(n_527) );
XOR2_X1 cordic_AddX_Add_g716 ( .a(cordic_AddX_Btemp1_1_), .b(cordic_AddX_Atemp_1_), .o(cordic_AddX_Add_n_18) );
XOR2_X1 cordic_AddX_g199 ( .a(cordic_AddX_Btemp_12_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_12_) );
BUF_X2 newInst_503 ( .a(newNet_502), .o(newNet_503) );
NAND2_Z01 cordic_SH1_srl_35_26_g1197 ( .a(cordic_SH1_srl_35_26_n_8), .b(cordic_SH1_srl_35_26_n_35), .o(cordic_SH1_srl_35_26_n_55) );
BUF_X2 newInst_849 ( .a(newNet_440), .o(newNet_849) );
BUF_X2 newInst_725 ( .a(newNet_724), .o(newNet_725) );
NAND2_Z01 cordic_SH2_srl_35_26_g1240 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_0_), .o(cordic_SH2_srl_35_26_n_9) );
BUF_X2 newInst_958 ( .a(newNet_957), .o(newNet_958) );
NAND2_Z01 g15273 ( .a(n_250), .b(n_251), .o(n_387) );
NAND2_Z01 cordic_pla_g302 ( .a(cordic_pla_n_1), .b(cordic_iteration_2_), .o(cordic_pla_n_9) );
NAND2_Z01 cordic_SH1_srl_35_26_g1148 ( .a(cordic_SH1_srl_35_26_n_90), .b(cordic_SH1_srl_35_26_n_18), .o(cordic_SH1_srl_35_26_n_104) );
BUF_X2 newInst_185 ( .a(newNet_184), .o(newNet_185) );
XOR2_X1 cordic_Add0_Add_g689 ( .a(cordic_Add0_n_2), .b(cordic_Add0_Atemp_1_), .o(cordic_Add0_Add_n_18) );
BUF_X2 newInst_321 ( .a(newNet_320), .o(newNet_321) );
BUF_X2 newInst_994 ( .a(newNet_993), .o(newNet_994) );
BUF_X2 newInst_714 ( .a(newNet_713), .o(newNet_714) );
NAND2_Z01 g13521 ( .a(Idsel), .b(Config_Reg_16_), .o(n_765) );
fflopd cordic_Angle_reg_0_ ( .CK(newNet_262), .D(cordic_n_115), .Q(cordic_Angle_0_) );
AND2_X1 g50 ( .a(n_830), .b(n_856), .o(PO_AD_14) );
fflopd Par_Sgnl_reg ( .CK(newNet_399), .D(n_501), .Q(Par_Sgnl) );
BUF_X2 newInst_1007 ( .a(newNet_1006), .o(newNet_1007) );
BUF_X2 newInst_252 ( .a(newNet_61), .o(newNet_252) );
fflopd Access_Address_1_reg_19_ ( .CK(newNet_1185), .D(n_456), .Q(Access_Address_1_19_) );
AND2_X1 g15634 ( .a(Access_Type_1_1_), .b(Access_Type_1_2_), .o(n_34) );
BUF_X2 newInst_976 ( .a(newNet_975), .o(newNet_976) );
AND2_X1 g360 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_34) );
NAND2_Z01 g15088 ( .a(n_4), .b(PI_AD_6), .o(n_520) );
BUF_X2 newInst_822 ( .a(newNet_821), .o(newNet_822) );
BUF_X2 newInst_589 ( .a(newNet_588), .o(newNet_589) );
BUF_X2 newInst_211 ( .a(newNet_210), .o(newNet_211) );
BUF_X2 newInst_305 ( .a(newNet_304), .o(newNet_305) );
INV_Z1 cordic_Add0_g57 ( .a(cordic_Add0_Btemp_4_), .o(cordic_Add0_n_5) );
BUF_X2 newInst_948 ( .a(newNet_947), .o(newNet_948) );
XNOR2_X1 cordic_AddY_Compl_g379 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_6_), .o(cordic_AddY_Compl_n_4) );
fflopd CoreOutputReg_reg_25_ ( .CK(newNet_629), .D(n_396), .Q(CoreOutputReg_25_) );
BUF_X2 newInst_842 ( .a(newNet_841), .o(newNet_842) );
fflopd CoreInput_reg_0_ ( .CK(newNet_833), .D(n_656), .Q(CoreInput_0_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1191 ( .a(cordic_SH1_srl_35_26_n_56), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_61) );
BUF_X2 newInst_217 ( .a(newNet_216), .o(newNet_217) );
BUF_X2 newInst_268 ( .a(newNet_267), .o(newNet_268) );
BUF_X2 newInst_74 ( .a(newNet_73), .o(newNet_74) );
NAND2_Z01 g15349 ( .a(CoreOutput_32_), .b(n_2), .o(n_312) );
BUF_X2 newInst_791 ( .a(newNet_790), .o(newNet_791) );
BUF_X2 newInst_68 ( .a(newNet_67), .o(newNet_68) );
BUF_X2 newInst_938 ( .a(newNet_937), .o(newNet_938) );
BUF_X2 newInst_998 ( .a(newNet_997), .o(newNet_998) );
BUF_X2 newInst_779 ( .a(newNet_778), .o(newNet_779) );
XOR2_X1 cordic_AddX_Add_g705 ( .a(cordic_AddX_Btemp1_11_), .b(cordic_AddX_Atemp_11_), .o(cordic_AddX_Add_n_29) );
XOR2_X1 g15500 ( .a(n_60), .b(n_61), .o(n_163) );
AND2_X1 g331 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_63) );
NAND2_Z01 g15103 ( .a(n_496), .b(n_276), .o(n_505) );
INV_X2 newInst_798 ( .a(newNet_99), .o(newNet_798) );
BUF_X2 newInst_985 ( .a(newNet_984), .o(newNet_985) );
INV_X1 g15506 ( .a(n_155), .o(n_154) );
NAND2_Z01 cordic_AddX_MUX_1_g298 ( .a(cordic_AddX_Y_1), .b(cordic_X_11_), .o(cordic_AddX_MUX_1_n_23) );
XOR2_X1 cordic_AddY_Add_g716 ( .a(cordic_AddY_Btemp1_1_), .b(cordic_AddY_Atemp_1_), .o(cordic_AddY_Add_n_18) );
NAND2_Z01 g13516 ( .a(Idsel), .b(Config_Reg_11_), .o(n_770) );
XOR2_X1 g13406 ( .a(n_873), .b(PO_AD_28), .o(n_874) );
NOR2_Z1 g15535 ( .a(n_108), .b(RESET), .o(n_135) );
XOR2_X1 g13399 ( .a(n_880), .b(PO_AD_4), .o(n_881) );
BUF_X2 newInst_1089 ( .a(newNet_1088), .o(newNet_1089) );
NAND2_Z01 cordic_AddX_g63 ( .a(cordic_AddX_n_3), .b(cordic_AddX_n_2), .o(CoreOutput_33_) );
NAND2_Z01 cordic_Add0_Add_g648 ( .a(cordic_Add0_Add_n_57), .b(cordic_Add0_Add_n_5), .o(cordic_Add0_Add_n_59) );
BUF_X2 newInst_2 ( .a(newNet_1), .o(newNet_2) );
INV_X1 g15649 ( .a(Dual_Cycle), .o(n_16) );
fflopd TAR_TRI_P_reg ( .CK(newNet_351), .D(n_337), .Q(TAR_TRI_P) );
NAND3_Z1 g15135 ( .a(n_327), .b(n_420), .c(n_10), .o(n_476) );
NAND2_Z01 g15449 ( .a(n_156), .b(Burst_Trans), .o(n_205) );
XNOR2_X1 cordic_AddY_Compl_g370 ( .a(cordic_AddY_Y_4), .b(cordic_AddY_Stemp_12_), .o(cordic_AddY_Compl_n_12) );
BUF_X2 newInst_1184 ( .a(newNet_1183), .o(newNet_1184) );
BUF_X2 newInst_294 ( .a(newNet_3), .o(newNet_294) );
NOR2_Z1 g15147 ( .a(n_444), .b(n_268), .o(n_465) );
NAND2_Z01 cordic_AddY_Add_g688 ( .a(cordic_AddY_Add_n_44), .b(cordic_AddY_Add_n_7), .o(cordic_AddY_Add_n_46) );
BUF_X2 newInst_527 ( .a(newNet_526), .o(newNet_527) );
NAND2_Z01 g15509 ( .a(n_116), .b(CBE_par_0_), .o(n_152) );
NAND2_Z01 cordic_SH1_srl_35_26_g1171 ( .a(cordic_SH1_srl_35_26_n_46), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_81) );
BUF_X2 newInst_827 ( .a(newNet_826), .o(newNet_827) );
NAND2_Z01 g15242 ( .a(n_274), .b(Access_Address_1_28_), .o(n_418) );
BUF_X2 newInst_156 ( .a(newNet_155), .o(newNet_156) );
NAND2_Z01 g15425 ( .a(n_186), .b(System_Busy), .o(n_276) );
fflopd Check_Data_Parity_reg ( .CK(newNet_1057), .D(n_372), .Q(Check_Data_Parity) );
NAND2_Z01 cordic_SH1_srl_35_26_g1173 ( .a(cordic_SH1_srl_35_26_n_57), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_79) );
NAND2_Z01 cordic_SH2_srl_35_26_g1201 ( .a(cordic_SH2_srl_35_26_n_16), .b(cordic_SH2_srl_35_26_n_28), .o(cordic_SH2_srl_35_26_n_51) );
BUF_X2 newInst_737 ( .a(newNet_736), .o(newNet_737) );
BUF_X2 newInst_399 ( .a(newNet_398), .o(newNet_399) );
NOR2_Z1 g15533 ( .a(n_87), .b(n_44), .o(n_123) );
NAND3_Z1 g15142 ( .a(n_362), .b(n_359), .c(n_10), .o(n_469) );
BUF_X2 newInst_1191 ( .a(newNet_933), .o(newNet_1191) );
NAND2_Z01 cordic_g434 ( .a(cordic_SumAngle_11_), .b(cordic_n_7), .o(cordic_n_73) );
BUF_X2 newInst_1200 ( .a(newNet_1199), .o(newNet_1200) );
XOR2_X1 cordic_AddY_Add_g715 ( .a(cordic_AddY_Btemp1_12_), .b(cordic_AddY_Atemp_12_), .o(cordic_AddY_Add_n_19) );
NOR2_Z1 cordic_SH1_srl_35_26_g1144 ( .a(cordic_SH1_srl_35_26_n_94), .b(cordic_SH1_srl_35_26_n_19), .o(cordic_BS1_12_) );
INV_X2 newInst_563 ( .a(newNet_123), .o(newNet_563) );
NAND2_Z01 cordic_g392 ( .a(cordic_n_76), .b(cordic_n_97), .o(cordic_n_115) );
BUF_X2 newInst_1173 ( .a(newNet_1172), .o(newNet_1173) );
NAND2_Z01 cordic_AddY_MUX_0_g295 ( .a(cordic_BS2_8_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_26) );
AND2_X1 g15544 ( .a(n_92), .b(Trdy_Wait_Cnt_0_), .o(n_127) );
NAND4_Z1 g14821 ( .a(n_212), .b(n_429), .c(n_687), .d(n_216), .o(n_698) );
XOR2_X1 g15596 ( .a(PI_AD_29), .b(PI_AD_3), .o(n_69) );
BUF_X2 newInst_748 ( .a(newNet_747), .o(newNet_748) );
BUF_X2 newInst_1091 ( .a(newNet_1090), .o(newNet_1091) );
NAND2_Z01 g15055 ( .a(n_473), .b(PI_AD_1), .o(n_553) );
NAND2_Z01 cordic_SH1_srl_35_26_g1126 ( .a(cordic_SH1_srl_35_26_n_119), .b(cordic_SH1_srl_35_26_n_60), .o(cordic_SH1_srl_35_26_n_126) );
BUF_X2 newInst_150 ( .a(newNet_149), .o(newNet_150) );
BUF_X2 newInst_142 ( .a(newNet_141), .o(newNet_142) );
NAND2_Z01 g15237 ( .a(n_274), .b(Access_Address_1_24_), .o(n_423) );
fflopd CoreOutputReg_reg_28_ ( .CK(newNet_621), .D(n_393), .Q(CoreOutputReg_28_) );
NAND2_Z01 cordic_Add0_MUX_1_g262 ( .a(cordic_Add0_MUX_1_n_8), .b(cordic_Add0_MUX_1_n_26), .o(cordic_Add0_Btemp_6_) );
BUF_X2 newInst_868 ( .a(newNet_867), .o(newNet_868) );
NAND2_Z01 g15257 ( .a(n_297), .b(n_298), .o(n_403) );
BUF_X2 newInst_134 ( .a(newNet_39), .o(newNet_134) );
BUF_X2 newInst_287 ( .a(newNet_56), .o(newNet_287) );
fflopd Access_Address_1_reg_18_ ( .CK(newNet_1186), .D(n_457), .Q(Access_Address_1_18_) );
NOR2_Z1 cordic_pla_g306 ( .a(cordic_iteration_3_), .b(cordic_iteration_2_), .o(cordic_pla_n_6) );
INV_X2 cordic_AddX_drc_bufs ( .a(cordic_AddX_n_0), .o(cordic_AddX_Y_2) );
BUF_X2 newInst_149 ( .a(newNet_148), .o(newNet_149) );
BUF_X2 newInst_231 ( .a(newNet_230), .o(newNet_231) );
BUF_X2 newInst_513 ( .a(newNet_512), .o(newNet_513) );
BUF_X2 newInst_181 ( .a(newNet_180), .o(newNet_181) );
NAND2_Z01 cordic_AddX_MUX_0_g305 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_3_), .o(cordic_AddX_MUX_0_n_16) );
NAND2_Z01 cordic_SH2_srl_35_26_g1203 ( .a(cordic_SH2_srl_35_26_n_22), .b(cordic_SH2_srl_35_26_n_31), .o(cordic_SH2_srl_35_26_n_50) );
BUF_X2 newInst_605 ( .a(newNet_604), .o(newNet_605) );
BUF_X2 newInst_300 ( .a(newNet_299), .o(newNet_300) );
NAND2_Z01 g13560 ( .a(n_712), .b(CoreOutputReg_14_), .o(n_727) );
BUF_X2 newInst_361 ( .a(newNet_360), .o(newNet_361) );
BUF_X2 newInst_80 ( .a(newNet_79), .o(newNet_80) );
NAND2_Z01 cordic_SH2_srl_35_26_g1233 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_8_), .o(cordic_SH2_srl_35_26_n_16) );
BUF_X2 newInst_1049 ( .a(newNet_1048), .o(newNet_1049) );
INV_Z1 cordic_Add0_g47 ( .a(cordic_Add0_Btemp_14_), .o(cordic_Add0_n_15) );
NAND2_Z01 cordic_Add0_MUX_1_g269 ( .a(cordic_AngleCin), .b(cordic_Angle_11_), .o(cordic_Add0_MUX_1_n_32) );
NAND2_Z01 cordic_AddY_MUX_0_g317 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_5_), .o(cordic_AddY_MUX_0_n_4) );
NAND2_Z01 cordic_AddY_Add_g724 ( .a(cordic_AddY_Btemp1_14_), .b(cordic_AddY_Atemp_14_), .o(cordic_AddY_Add_n_10) );
XOR2_X1 g13390 ( .a(n_889), .b(PO_AD_10), .o(n_890) );
AND2_X1 g353 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_41) );
NAND2_Z01 g15302 ( .a(n_281), .b(n_222), .o(n_353) );
XOR2_X1 cordic_AddX_Compl_g344 ( .a(cordic_AddX_Compl_n_35), .b(cordic_AddX_Compl_n_3), .o(CoreOutput_28_) );
fflopd Config_Reg_reg_2_ ( .CK(newNet_904), .D(n_666), .Q(Config_Reg_2_) );
NAND2_Z01 cordic_Add0_MUX_0_g299 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_9_), .o(cordic_Add0_MUX_0_n_4) );
BUF_X2 newInst_463 ( .a(newNet_462), .o(newNet_463) );
AND2_X1 cordic_AddY_g64 ( .a(cordic_AddY_Y_3), .b(cordic_AddY_n_1), .o(cordic_AddY_n_3) );
AND2_X1 cordic_AddX_Compl_g341 ( .a(cordic_AddX_Compl_n_39), .b(cordic_AddX_Compl_n_8), .o(cordic_AddX_Compl_n_41) );
AND2_X1 cordic_pla_g291 ( .a(cordic_pla_n_4), .b(cordic_iteration_3_), .o(cordic_pla_n_23) );
NAND2_Z01 cordic_SH1_srl_35_26_g1240 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_0_), .o(cordic_SH1_srl_35_26_n_9) );
BUF_X2 newInst_545 ( .a(newNet_544), .o(newNet_545) );
fflopd Access_Address_1_reg_26_ ( .CK(newNet_1143), .D(n_477), .Q(Access_Address_1_26_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1114 ( .a(cordic_SH1_srl_35_26_n_127), .b(cordic_iteration_3_), .o(cordic_BS1_11_) );
AND2_X1 g336 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_58) );
BUF_X2 newInst_225 ( .a(newNet_224), .o(newNet_225) );
fflopd CoreOutputReg_reg_14_ ( .CK(newNet_704), .D(n_409), .Q(CoreOutputReg_14_) );
NAND2_Z01 g15014 ( .a(n_505), .b(n_537), .o(n_568) );
NAND2_Z01 g13514 ( .a(Idsel), .b(Config_Reg_18_), .o(n_772) );
NAND2_Z01 cordic_Add0_Add_g704 ( .a(cordic_Add0_n_3), .b(cordic_Add0_Atemp_2_), .o(cordic_Add0_Add_n_3) );
fflopd State_reg_1_ ( .CK(newNet_380), .D(n_709), .Q(State_1_) );
NOR2_Z1 cordic_g472 ( .a(Issue_Rst), .b(cordic_iteration_0_), .o(cordic_n_35) );
NAND2_Z01 cordic_Add0_MUX_0_g261 ( .a(cordic_Add0_MUX_0_n_28), .b(cordic_Add0_MUX_0_n_14), .o(cordic_Add0_Atemp_0_) );
NOR2_Z1 g15310 ( .a(n_221), .b(n_154), .o(n_384) );
NAND2_Z01 g15284 ( .a(n_274), .b(Access_Address_1_16_), .o(n_371) );
NAND2_Z01 g14958 ( .a(n_572), .b(Config_Reg_24_), .o(n_619) );
NAND2_Z01 g13564 ( .a(n_712), .b(CoreOutputReg_10_), .o(n_723) );
NAND2_Z01 cordic_AddY_MUX_1_g319 ( .a(cordic_BS2_4_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_2) );
NAND2_Z01 cordic_g405 ( .a(cordic_n_58), .b(cordic_n_81), .o(cordic_n_102) );
AND2_X1 g344 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_50) );
NAND2_Z01 cordic_Add0_MUX_0_g266 ( .a(cordic_Add0_MUX_0_n_21), .b(cordic_Add0_MUX_0_n_4), .o(cordic_Add0_Atemp_9_) );
BUF_X2 newInst_886 ( .a(newNet_252), .o(newNet_886) );
NAND2_Z01 cordic_SH2_srl_35_26_g1208 ( .a(cordic_SH2_srl_35_26_n_4), .b(cordic_SH2_srl_35_26_n_24), .o(cordic_SH2_srl_35_26_n_46) );
NAND2_Z01 cordic_Add0_MUX_0_g280 ( .a(cordic_tanangle_12_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_23) );
BUF_X2 newInst_666 ( .a(newNet_78), .o(newNet_666) );
NAND2_Z01 cordic_Add0_MUX_1_g273 ( .a(cordic_AngleCin), .b(cordic_Angle_0_), .o(cordic_Add0_MUX_1_n_28) );
INV_X2 newInst_1080 ( .a(newNet_1079), .o(newNet_1080) );
AND2_X1 g13426 ( .a(n_855), .b(TAR_TRI_A), .o(n_856) );
XOR2_X1 cordic_AddY_g201 ( .a(cordic_AddY_Btemp_0_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_0_) );
XOR2_X1 cordic_AddX_Compl_g352 ( .a(cordic_AddX_Compl_n_27), .b(cordic_AddX_Compl_n_6), .o(CoreOutput_24_) );
BUF_X2 newInst_1060 ( .a(newNet_1059), .o(newNet_1060) );
BUF_X2 newInst_129 ( .a(newNet_128), .o(newNet_129) );
BUF_X2 newInst_343 ( .a(newNet_342), .o(newNet_343) );
NAND2_Z01 cordic_SH2_srl_35_26_g1154 ( .a(cordic_SH2_srl_35_26_n_87), .b(cordic_SH2_srl_35_26_n_75), .o(cordic_SH2_srl_35_26_n_99) );
BUF_X2 newInst_28 ( .a(newNet_27), .o(newNet_28) );
AND2_X1 g40 ( .a(n_826), .b(n_856), .o(PO_AD_24) );
XOR2_X1 g15599 ( .a(PI_AD_60), .b(PI_AD_39), .o(n_66) );
BUF_X2 newInst_665 ( .a(newNet_664), .o(newNet_665) );
BUF_X2 newInst_805 ( .a(newNet_361), .o(newNet_805) );
NAND2_Z01 cordic_SH2_srl_35_26_g1190 ( .a(cordic_SH2_srl_35_26_n_52), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_62) );
fflopd Config_Reg_reg_10_ ( .CK(newNet_1047), .D(n_637), .Q(Config_Reg_10_) );
NAND2_Z01 cordic_g441 ( .a(cordic_SumAngle_3_), .b(cordic_n_7), .o(cordic_n_66) );
NAND2_Z01 cordic_SH2_srl_35_26_g1215 ( .a(cordic_iteration_0_), .b(cordic_X_10_), .o(cordic_SH2_srl_35_26_n_37) );
NAND2_Z01 cordic_AddX_Compl_g365 ( .a(cordic_AddX_Compl_n_11), .b(cordic_AddX_Compl_n_1), .o(cordic_AddX_Compl_n_17) );
NAND2_Z01 cordic_SH2_srl_35_26_g1221 ( .a(cordic_iteration_0_), .b(cordic_X_14_), .o(cordic_SH2_srl_35_26_n_31) );
AND2_X1 g347 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_47) );
BUF_X2 newInst_53 ( .a(newNet_52), .o(newNet_53) );
AND2_X1 cordic_pla_g274 ( .a(cordic_pla_n_31), .b(cordic_pla_n_25), .o(cordic_tanangle_4_) );
BUF_X2 newInst_114 ( .a(newNet_113), .o(newNet_114) );
NAND2_Z01 cordic_AddY_MUX_1_g301 ( .a(cordic_AddY_Y_1), .b(cordic_Y_13_), .o(cordic_AddY_MUX_1_n_20) );
NAND3_Z1 g15572 ( .a(n_25), .b(n_49), .c(DevSel_Wait_Cnt_0_), .o(n_93) );
BUF_X2 newInst_282 ( .a(newNet_281), .o(newNet_282) );
BUF_X2 newInst_680 ( .a(newNet_679), .o(newNet_680) );
NAND2_Z01 cordic_AddY_MUX_1_g285 ( .a(cordic_AddY_MUX_1_n_1), .b(cordic_AddY_MUX_1_n_19), .o(cordic_AddY_Btemp_10_) );
NAND2_Z01 g14951 ( .a(n_572), .b(Config_Reg_17_), .o(n_626) );
fflopd CoreOutputReg_reg_9_ ( .CK(newNet_553), .D(n_373), .Q(CoreOutputReg_9_) );
NAND2_Z01 cordic_AddX_MUX_0_g276 ( .a(cordic_AddX_MUX_0_n_29), .b(cordic_AddX_MUX_0_n_14), .o(cordic_AddX_Atemp_2_) );
XOR2_X1 g15586 ( .a(PI_AD_20), .b(PI_AD_19), .o(n_79) );
XOR2_X1 cordic_Add0_Compl_g338 ( .a(cordic_Add0_Compl_n_41), .b(cordic_Add0_Compl_n_13), .o(cordic_SumAngle_14_) );
NOR2_Z1 cordic_g333 ( .a(cordic_n_119), .b(Issue_Rst), .o(cordic_n_122) );
BUF_X2 newInst_674 ( .a(newNet_673), .o(newNet_674) );
XOR2_X1 cordic_AddY_Compl_g356 ( .a(cordic_AddY_Compl_n_23), .b(cordic_AddY_Compl_n_5), .o(CoreOutput_5_) );
BUF_X2 newInst_478 ( .a(newNet_477), .o(newNet_478) );
fflopd Core_Cnt_reg_1_ ( .CK(newNet_543), .D(n_123), .Q(Core_Cnt_1_) );
NOR2_Z1 cordic_SH1_srl_35_26_g1150 ( .a(cordic_SH1_srl_35_26_n_89), .b(cordic_iteration_3_), .o(cordic_BS1_14_) );
NAND2_Z04 g15007 ( .a(n_563), .b(n_488), .o(n_572) );
NAND4_Z1 cordic_SH2_srl_35_26_g1106 ( .a(cordic_SH2_srl_35_26_n_70), .b(cordic_SH2_srl_35_26_n_116), .c(cordic_SH2_srl_35_26_n_143), .d(cordic_SH2_srl_35_26_n_72), .o(cordic_BS2_0_) );
BUF_X2 newInst_551 ( .a(newNet_550), .o(newNet_551) );
NOR2_X3 g15477 ( .a(n_140), .b(RESET), .o(n_188) );
XOR2_X1 cordic_Add0_Add_g652 ( .a(cordic_Add0_Add_n_53), .b(cordic_Add0_Add_n_17), .o(cordic_Add0_Stemp_8_) );
BUF_X2 newInst_1125 ( .a(newNet_1124), .o(newNet_1125) );
BUF_X2 newInst_1192 ( .a(newNet_1191), .o(newNet_1192) );
NAND2_Z01 cordic_AddX_Add_g699 ( .a(cordic_AddX_Add_n_34), .b(cordic_AddX_Add_n_18), .o(cordic_AddX_Add_n_35) );
BUF_X2 newInst_176 ( .a(newNet_175), .o(newNet_176) );
BUF_X2 newInst_1146 ( .a(newNet_1145), .o(newNet_1146) );
NAND2_Z01 cordic_AddY_MUX_1_g310 ( .a(cordic_BS2_12_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_11) );
fflopd DevSel_Wait_Cnt_reg_2_ ( .CK(newNet_492), .D(n_493), .Q(DevSel_Wait_Cnt_2_) );
XOR2_X1 cordic_AddX_Compl_g371 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_1_), .o(cordic_AddX_Compl_n_11) );
NAND3_Z1 g15130 ( .a(n_329), .b(n_424), .c(n_10), .o(n_480) );
BUF_X2 newInst_318 ( .a(newNet_317), .o(newNet_318) );
NOR2_Z1 g13439 ( .a(n_807), .b(n_710), .o(n_843) );
BUF_X2 newInst_1137 ( .a(newNet_1136), .o(newNet_1137) );
NAND2_Z01 cordic_AddY_MUX_0_g307 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_2_), .o(cordic_AddY_MUX_0_n_14) );
NAND2_Z01 g14909 ( .a(n_612), .b(n_540), .o(n_665) );
INV_Z1 g8019 ( .a(CoreOutputReg_32_), .o(n_899) );
NAND2_Z01 cordic_SH2_srl_35_26_g1122 ( .a(cordic_SH2_srl_35_26_n_113), .b(cordic_SH2_srl_35_26_n_88), .o(cordic_SH2_srl_35_26_n_130) );
NAND2_Z01 g15616 ( .a(Core_Cnt_0_), .b(Core_Cnt_1_), .o(n_52) );
NAND2_Z01 g15308 ( .a(n_267), .b(n_109), .o(n_385) );
NOR2_Z1 cordic_SH2_srl_35_26_g1194 ( .a(cordic_SH2_srl_35_26_n_41), .b(cordic_SH2_srl_35_26_n_19), .o(cordic_BS2_15_) );
NOR2_Z1 g15555 ( .a(n_45), .b(RESET), .o(n_118) );
NAND2_Z02 g15430 ( .a(n_212), .b(n_111), .o(n_274) );
BUF_X2 newInst_811 ( .a(newNet_810), .o(newNet_811) );
NOR2_Z1 g15467 ( .a(n_121), .b(RESET), .o(n_211) );
NAND2_Z01 g15461 ( .a(n_146), .b(n_47), .o(n_197) );
NAND2_Z01 cordic_AddX_Add_g728 ( .a(cordic_AddX_Btemp1_3_), .b(cordic_AddX_Atemp_3_), .o(cordic_AddX_Add_n_6) );
BUF_X2 newInst_477 ( .a(newNet_46), .o(newNet_477) );
BUF_X2 newInst_381 ( .a(newNet_243), .o(newNet_381) );
NAND2_Z01 cordic_AddY_Add_g731 ( .a(cordic_AddY_Btemp1_2_), .b(cordic_AddY_Atemp_2_), .o(cordic_AddY_Add_n_3) );
AND2_X1 g14832 ( .a(n_686), .b(n_139), .o(n_689) );
BUF_X2 newInst_457 ( .a(newNet_456), .o(newNet_457) );
NAND2_Z01 g15385 ( .a(n_214), .b(CoreOutputReg_26_), .o(n_265) );
fflopd Config_Reg_reg_1_ ( .CK(newNet_983), .D(n_677), .Q(Config_Reg_1_) );
NAND4_Z1 cordic_SH2_srl_35_26_g1103 ( .a(cordic_SH2_srl_35_26_n_78), .b(cordic_SH2_srl_35_26_n_122), .c(cordic_SH2_srl_35_26_n_139), .d(cordic_SH2_srl_35_26_n_77), .o(cordic_BS2_3_) );
BUF_X2 newInst_544 ( .a(newNet_520), .o(newNet_544) );
BUF_X2 newInst_497 ( .a(newNet_496), .o(newNet_497) );
BUF_X2 newInst_506 ( .a(newNet_505), .o(newNet_506) );
NAND2_Z01 cordic_AddY_MUX_1_g292 ( .a(cordic_AddY_Y_1), .b(cordic_Y_2_), .o(cordic_AddY_MUX_1_n_29) );
BUF_X2 newInst_18 ( .a(newNet_17), .o(newNet_18) );
fflopd cordic_X_reg_7_ ( .CK(newNet_24), .D(cordic_n_31), .Q(cordic_X_7_) );
BUF_X2 newInst_645 ( .a(newNet_158), .o(newNet_645) );
AND2_X1 g39 ( .a(n_828), .b(n_856), .o(PO_AD_25) );
BUF_X2 newInst_789 ( .a(newNet_788), .o(newNet_789) );
NOR2_Z1 g15566 ( .a(n_51), .b(State_1_), .o(n_110) );
NAND2_Z01 cordic_SH1_srl_35_26_g1202 ( .a(cordic_SH1_srl_35_26_n_9), .b(cordic_SH1_srl_35_26_n_34), .o(cordic_SH1_srl_35_26_n_49) );
BUF_X2 newInst_556 ( .a(newNet_389), .o(newNet_556) );
fflopd cordic_X_reg_13_ ( .CK(newNet_162), .D(cordic_n_56), .Q(cordic_X_13_) );
BUF_X2 newInst_587 ( .a(newNet_586), .o(newNet_587) );
NAND2_Z01 cordic_g417 ( .a(Issue_Rst), .b(CoreInput_2_), .o(cordic_n_90) );
BUF_X2 newInst_63 ( .a(newNet_17), .o(newNet_63) );
NAND2_Z01 g15423 ( .a(n_201), .b(n_142), .o(n_230) );
AND2_X1 g15132 ( .a(n_436), .b(n_138), .o(n_495) );
AND2_X1 g45 ( .a(n_834), .b(n_856), .o(PO_AD_19) );
NAND2_Z01 cordic_AddX_Add_g734 ( .a(cordic_AddX_Btemp1_6_), .b(cordic_AddX_Atemp_6_), .o(cordic_AddX_Add_n_0) );
BUF_X2 newInst_929 ( .a(newNet_928), .o(newNet_929) );
NAND2_Z01 cordic_AddY_Add_g657 ( .a(cordic_AddY_Add_n_76), .b(cordic_AddY_Add_n_25), .o(cordic_AddY_Add_n_77) );
BUF_X2 newInst_922 ( .a(newNet_921), .o(newNet_922) );
BUF_X2 newInst_297 ( .a(newNet_296), .o(newNet_297) );
NAND2_Z01 g13545 ( .a(n_712), .b(CoreOutputReg_7_), .o(n_741) );
AND2_X1 cordic_AddX_Compl_g361 ( .a(cordic_AddX_Compl_n_19), .b(cordic_AddX_Compl_n_16), .o(cordic_AddX_Compl_n_21) );
NAND2_Z01 g15050 ( .a(n_486), .b(TAR_TRI_A), .o(n_558) );
BUF_X2 newInst_167 ( .a(newNet_166), .o(newNet_167) );
NAND2_Z01 g15553 ( .a(n_28), .b(DevSel_Wait_Cnt_2_), .o(n_103) );
BUF_X2 newInst_1148 ( .a(newNet_1147), .o(newNet_1148) );
BUF_X2 newInst_992 ( .a(newNet_991), .o(newNet_992) );
NAND2_Z01 g15357 ( .a(CoreOutput_16_), .b(n_188), .o(n_304) );
BUF_X2 newInst_962 ( .a(newNet_961), .o(newNet_962) );
BUF_X2 newInst_401 ( .a(newNet_400), .o(newNet_401) );
fflopd Access_Address_1_reg_23_ ( .CK(newNet_1160), .D(n_480), .Q(Access_Address_1_23_) );
fflopd cordic_iteration_reg_1_ ( .CK(newNet_290), .D(cordic_n_120), .Q(cordic_iteration_1_) );
BUF_X2 newInst_717 ( .a(newNet_716), .o(newNet_717) );
NAND2_Z01 g15457 ( .a(n_129), .b(Trdy_Wait_Cnt_1_), .o(n_201) );
NAND2_Z01 g15361 ( .a(n_214), .b(CoreOutputReg_18_), .o(n_300) );
NAND2_Z01 g15059 ( .a(n_473), .b(PI_AD_23), .o(n_549) );
NAND4_Z1 g15110 ( .a(n_279), .b(n_220), .c(n_448), .d(n_139), .o(n_498) );
NAND2_Z01 g13488 ( .a(n_731), .b(n_764), .o(n_796) );
NAND2_Z01 cordic_AddX_MUX_1_g275 ( .a(cordic_AddX_MUX_1_n_15), .b(cordic_AddX_MUX_1_n_30), .o(cordic_AddX_Btemp_9_) );
NAND2_Z01 g15330 ( .a(n_3), .b(PI_AD_22), .o(n_331) );
NOR2_Z2 g15483 ( .a(n_134), .b(PI_FRAME_L), .o(n_184) );
XNOR2_X1 cordic_AddX_Compl_g368 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_2_), .o(cordic_AddX_Compl_n_14) );
BUF_X2 newInst_611 ( .a(newNet_610), .o(newNet_611) );
AND2_X1 cordic_AddX_Compl_g353 ( .a(cordic_AddX_Compl_n_27), .b(cordic_AddX_Compl_n_6), .o(cordic_AddX_Compl_n_29) );
BUF_X2 newInst_576 ( .a(newNet_575), .o(newNet_576) );
BUF_X2 newInst_423 ( .a(newNet_422), .o(newNet_423) );
BUF_X2 newInst_257 ( .a(newNet_256), .o(newNet_257) );
BUF_X2 newInst_202 ( .a(newNet_201), .o(newNet_202) );
NAND2_Z01 cordic_SH1_srl_35_26_g1236 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_10_), .o(cordic_SH1_srl_35_26_n_13) );
BUF_X2 newInst_635 ( .a(newNet_634), .o(newNet_635) );
fflopd CoreOutputReg_reg_29_ ( .CK(newNet_619), .D(n_392), .Q(CoreOutputReg_29_) );
NAND2_Z01 g14926 ( .a(n_595), .b(n_525), .o(n_648) );
BUF_X2 newInst_30 ( .a(newNet_29), .o(newNet_30) );
NAND2_Z01 g13538 ( .a(n_712), .b(CoreOutputReg_22_), .o(n_748) );
NAND2_Z01 cordic_Add0_MUX_0_g276 ( .a(cordic_tanangle_6_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_27) );
NAND2_Z01 cordic_SH2_srl_35_26_g1143 ( .a(cordic_SH2_srl_35_26_n_92), .b(cordic_SH2_srl_35_26_n_18), .o(cordic_SH2_srl_35_26_n_109) );
BUF_X2 newInst_1040 ( .a(newNet_1039), .o(newNet_1040) );
fflopd Config_Reg_reg_9_ ( .CK(newNet_848), .D(n_657), .Q(Config_Reg_9_) );
NAND2_Z01 g15262 ( .a(n_286), .b(n_287), .o(n_398) );
BUF_X2 newInst_846 ( .a(newNet_845), .o(newNet_846) );
NAND2_Z01 g15281 ( .a(n_239), .b(n_240), .o(n_374) );
NAND2_Z01 g15291 ( .a(n_275), .b(Access_Type_1_1_), .o(n_364) );
BUF_X2 newInst_1023 ( .a(newNet_1022), .o(newNet_1023) );
NAND2_Z01 cordic_Add0_MUX_1_g283 ( .a(cordic_AngleCin), .b(cordic_Angle_13_), .o(cordic_Add0_MUX_1_n_18) );
BUF_X2 newInst_720 ( .a(newNet_638), .o(newNet_720) );
AND2_X1 cordic_AddY_Compl_g339 ( .a(cordic_AddY_Compl_n_41), .b(cordic_AddY_Compl_n_13), .o(cordic_AddY_Compl_n_43) );
XOR2_X1 cordic_AddY_Add_g659 ( .a(cordic_AddY_Add_n_73), .b(cordic_AddY_Add_n_22), .o(cordic_AddY_Stemp_14_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1134 ( .a(cordic_SH2_srl_35_26_n_98), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_118) );
BUF_X2 newInst_1051 ( .a(newNet_1050), .o(newNet_1051) );
XOR2_X1 cordic_AddY_Add_g671 ( .a(cordic_AddY_Add_n_61), .b(cordic_AddY_Add_n_27), .o(cordic_AddY_Stemp_10_) );
BUF_X2 newInst_439 ( .a(newNet_438), .o(newNet_439) );
fflopd Access_Address_1_reg_17_ ( .CK(newNet_1187), .D(n_458), .Q(Access_Address_1_17_) );
INV_X1 cordic_SH2_srl_35_26_g1250 ( .a(cordic_iteration_2_), .o(cordic_SH2_srl_35_26_n_2) );
XOR2_X1 cordic_AddY_Add_g698 ( .a(cordic_AddY_Add_n_34), .b(cordic_AddY_Add_n_18), .o(cordic_AddY_Stemp_1_) );
BUF_X2 newInst_209 ( .a(newNet_208), .o(newNet_209) );
NAND2_Z01 cordic_AddY_MUX_1_g288 ( .a(cordic_AddY_MUX_1_n_16), .b(cordic_AddY_MUX_1_n_17), .o(cordic_AddY_Btemp_3_) );
NAND2_Z01 g15093 ( .a(n_473), .b(PI_AD_0), .o(n_515) );
AND2_X1 g34 ( .a(n_845), .b(n_856), .o(PO_AD_30) );
XOR2_X1 cordic_AddX_Add_g692 ( .a(cordic_AddX_Add_n_40), .b(cordic_AddX_Add_n_24), .o(cordic_AddX_Stemp_3_) );
BUF_X2 newInst_101 ( .a(newNet_100), .o(newNet_101) );
NAND2_Z01 cordic_g420 ( .a(Issue_Rst), .b(CoreInput_5_), .o(cordic_n_87) );
NAND2_Z01 g14982 ( .a(n_571), .b(CoreInput_1_), .o(n_595) );
BUF_X2 newInst_106 ( .a(newNet_105), .o(newNet_106) );
INV_X1 cordic_SH2_srl_35_26_g1151 ( .a(cordic_SH2_srl_35_26_n_101), .o(cordic_SH2_srl_35_26_n_100) );
INV_Z1 cordic_Add0_g52 ( .a(cordic_Add0_Btemp_9_), .o(cordic_Add0_n_10) );
NAND2_Z01 cordic_Add0_Add_g671 ( .a(cordic_Add0_Add_n_35), .b(cordic_Add0_Add_n_20), .o(cordic_Add0_Add_n_36) );
fflopd CoreOutputReg_reg_4_ ( .CK(newNet_579), .D(n_378), .Q(CoreOutputReg_4_) );
fflopd CoreInput_reg_2_ ( .CK(newNet_774), .D(n_647), .Q(CoreInput_2_) );
NOR3_Z1 g15225 ( .a(n_191), .b(n_226), .c(n_110), .o(n_429) );
NAND2_Z01 g13481 ( .a(n_744), .b(n_765), .o(n_803) );
BUF_X2 newInst_273 ( .a(newNet_272), .o(newNet_273) );
NAND2_Z01 cordic_SH2_srl_35_26_g1167 ( .a(cordic_SH2_srl_35_26_n_50), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_85) );
INV_X1 g15626 ( .a(n_37), .o(n_38) );
INV_X1 drc_bufs15658 ( .a(n_7), .o(n_4) );
INV_Z1 cordic_Add0_g60 ( .a(cordic_Add0_Btemp_1_), .o(cordic_Add0_n_2) );
INV_X2 newInst_234 ( .a(newNet_163), .o(newNet_234) );
NAND3_Z1 cordic_pla_g272 ( .a(cordic_pla_n_17), .b(cordic_pla_n_18), .c(cordic_pla_n_23), .o(cordic_tanangle_8_) );
XOR2_X1 cordic_AddX_Add_g665 ( .a(cordic_AddX_Add_n_67), .b(cordic_AddX_Add_n_19), .o(cordic_AddX_Stemp_12_) );
BUF_X2 newInst_522 ( .a(newNet_429), .o(newNet_522) );
XOR2_X1 g15605 ( .a(PI_AD_42), .b(PI_AD_34), .o(n_60) );
BUF_X2 newInst_786 ( .a(newNet_785), .o(newNet_786) );
NAND2_Z01 cordic_AddX_MUX_1_g319 ( .a(cordic_BS1_4_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_2) );
NAND2_Z01 cordic_Add0_MUX_1_g296 ( .a(cordic_tanangle_4_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_5) );
BUF_X2 newInst_729 ( .a(newNet_247), .o(newNet_729) );
fflopd PAR_Int_reg ( .CK(newNet_446), .D(n_683), .Q(PAR_Int) );
BUF_X2 newInst_51 ( .a(newNet_16), .o(newNet_51) );
BUF_X2 newInst_329 ( .a(newNet_328), .o(newNet_329) );
BUF_X2 newInst_188 ( .a(newNet_187), .o(newNet_188) );
NAND3_Z1 g15145 ( .a(n_361), .b(n_356), .c(n_10), .o(n_466) );
NAND2_Z01 cordic_AddX_MUX_1_g307 ( .a(cordic_BS1_2_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_14) );
fflopd PO_PERR_L_reg ( .CK(newNet_1198), .D(n_859), .Q(PO_PERR_L) );
XOR2_X1 g15162 ( .a(n_340), .b(n_341), .o(n_450) );
NAND2_Z01 cordic_SH2_srl_35_26_g1173 ( .a(cordic_SH2_srl_35_26_n_57), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_79) );
XOR2_X1 g13419 ( .a(n_860), .b(CBE_par_3_), .o(n_861) );
XNOR2_X1 cordic_AddX_Compl_g374 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_13_), .o(cordic_AddX_Compl_n_8) );
NAND2_Z01 cordic_SH2_srl_35_26_g1222 ( .a(cordic_iteration_0_), .b(cordic_X_5_), .o(cordic_SH2_srl_35_26_n_30) );
BUF_X2 newInst_107 ( .a(newNet_106), .o(newNet_107) );
XOR2_X1 g15320 ( .a(n_161), .b(n_162), .o(n_340) );
INV_X1 g15642 ( .a(Access_Address_1_18_), .o(n_23) );
XOR2_X1 cordic_AddY_Add_g704 ( .a(cordic_AddY_Btemp1_7_), .b(cordic_AddY_Atemp_7_), .o(cordic_AddY_Add_n_30) );
NAND2_Z01 cordic_SH2_srl_35_26_g1138 ( .a(cordic_SH2_srl_35_26_n_96), .b(cordic_SH2_srl_35_26_n_18), .o(cordic_SH2_srl_35_26_n_114) );
BUF_X2 newInst_741 ( .a(newNet_740), .o(newNet_741) );
XOR2_X1 cordic_AddY_Compl_g340 ( .a(cordic_AddY_Compl_n_39), .b(cordic_AddY_Compl_n_8), .o(CoreOutput_13_) );
NAND2_Z01 g15377 ( .a(CoreOutput_24_), .b(n_2), .o(n_284) );
BUF_X2 newInst_655 ( .a(newNet_654), .o(newNet_655) );
BUF_X2 newInst_368 ( .a(newNet_367), .o(newNet_368) );
BUF_X2 newInst_139 ( .a(newNet_138), .o(newNet_139) );
BUF_X2 newInst_1071 ( .a(newNet_425), .o(newNet_1071) );
INV_X1 cordic_SH2_srl_35_26_g1119 ( .a(cordic_SH2_srl_35_26_n_132), .o(cordic_SH2_srl_35_26_n_133) );
BUF_X2 newInst_636 ( .a(newNet_592), .o(newNet_636) );
NAND3_Z1 g15154 ( .a(n_234), .b(n_370), .c(n_10), .o(n_458) );
BUF_X2 newInst_703 ( .a(newNet_702), .o(newNet_703) );
fflopd Set_Data_Parity_reg ( .CK(newNet_397), .D(n_574), .Q(Set_Data_Parity) );
BUF_X2 newInst_812 ( .a(newNet_811), .o(newNet_812) );
NAND2_Z01 cordic_AddX_Add_g670 ( .a(cordic_AddX_Add_n_62), .b(cordic_AddX_Add_n_13), .o(cordic_AddX_Add_n_64) );
NAND2_Z01 cordic_SH1_srl_35_26_g1153 ( .a(cordic_SH1_srl_35_26_n_67), .b(cordic_SH1_srl_35_26_n_38), .o(cordic_SH1_srl_35_26_n_101) );
XOR2_X1 g13414 ( .a(n_865), .b(PO_AD_27), .o(n_866) );
XNOR2_X1 cordic_AddX_Compl_g380 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_11_), .o(cordic_AddX_Compl_n_3) );
BUF_X2 newInst_144 ( .a(newNet_143), .o(newNet_144) );
NAND2_Z01 g15071 ( .a(n_495), .b(PO_STOP_L), .o(n_537) );
BUF_X2 newInst_911 ( .a(newNet_910), .o(newNet_911) );
fflopd cordic_Y_reg_9_ ( .CK(newNet_202), .D(cordic_n_78), .Q(cordic_Y_9_) );
NAND2_Z01 g14898 ( .a(n_623), .b(n_552), .o(n_676) );
XOR2_X1 cordic_AddX_g204 ( .a(cordic_AddX_Btemp_6_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_6_) );
BUF_X2 newInst_671 ( .a(newNet_101), .o(newNet_671) );
NAND3_Z1 g15139 ( .a(n_238), .b(n_419), .c(n_10), .o(n_472) );
NAND3_Z1 cordic_SH2_srl_35_26_g1212 ( .a(cordic_iteration_1_), .b(cordic_SH2_srl_35_26_n_0), .c(cordic_X_15_), .o(cordic_SH2_srl_35_26_n_38) );
NAND2_Z01 cordic_SH1_srl_35_26_g1145 ( .a(cordic_SH1_srl_35_26_n_95), .b(cordic_SH1_srl_35_26_n_20), .o(cordic_SH1_srl_35_26_n_107) );
BUF_X2 newInst_987 ( .a(newNet_176), .o(newNet_987) );
BUF_X2 newInst_379 ( .a(newNet_378), .o(newNet_379) );
XNOR2_X1 cordic_Add0_Compl_g366 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_3_), .o(cordic_Add0_Compl_n_16) );
NOR2_Z1 g13448 ( .a(n_801), .b(n_710), .o(n_834) );
AND2_X1 cordic_pla_g279 ( .a(cordic_pla_n_31), .b(cordic_pla_n_19), .o(cordic_tanangle_5_) );
NAND2_Z01 cordic_AddY_Add_g661 ( .a(cordic_AddY_Add_n_71), .b(cordic_AddY_Add_n_12), .o(cordic_AddY_Add_n_73) );
NAND2_Z01 cordic_AddY_MUX_0_g282 ( .a(cordic_AddY_MUX_0_n_22), .b(cordic_AddY_MUX_0_n_5), .o(cordic_AddY_Atemp_6_) );
NAND2_Z01 g15419 ( .a(n_183), .b(n_156), .o(n_280) );
NAND2_Z01 g14966 ( .a(n_572), .b(Config_Reg_31_), .o(n_611) );
BUF_X2 newInst_198 ( .a(newNet_197), .o(newNet_198) );
NAND2_Z01 g13500 ( .a(n_745), .b(n_780), .o(n_784) );
BUF_X2 newInst_200 ( .a(newNet_199), .o(newNet_200) );
NAND2_Z01 g15238 ( .a(n_274), .b(Access_Address_1_26_), .o(n_422) );
NAND2_Z01 cordic_AddX_Add_g720 ( .a(cordic_AddX_Btemp1_11_), .b(cordic_AddX_Atemp_11_), .o(cordic_AddX_Add_n_14) );
NAND2_Z01 cordic_AddX_MUX_0_g314 ( .a(cordic_AddX_MUX_0_n_0), .b(cordic_X_15_), .o(cordic_AddX_MUX_0_n_7) );
NOR2_Z1 cordic_g458 ( .a(cordic_n_3), .b(Issue_Rst), .o(cordic_n_49) );
NAND2_Z01 g15232 ( .a(n_274), .b(Access_Address_1_19_), .o(n_428) );
INV_X1 g15657 ( .a(PI_FRAME_L), .o(n_8) );
NAND2_Z01 cordic_AddY_MUX_0_g304 ( .a(cordic_BS2_3_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_17) );
NAND2_Z01 cordic_Add0_MUX_1_g258 ( .a(cordic_Add0_MUX_1_n_14), .b(cordic_Add0_MUX_1_n_30), .o(cordic_Add0_Btemp_1_) );
AND2_X1 cordic_AddY_Compl_g345 ( .a(cordic_AddY_Compl_n_35), .b(cordic_AddY_Compl_n_3), .o(cordic_AddY_Compl_n_37) );
NAND2_Z01 cordic_AddX_MUX_0_g295 ( .a(cordic_BS1_8_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_26) );
NOR2_Z1 g15438 ( .a(n_6), .b(PI_REQ64_L), .o(n_221) );
NAND2_Z01 g15370 ( .a(CoreOutput_21_), .b(n_188), .o(n_291) );
NAND2_Z01 cordic_Add0_MUX_0_g281 ( .a(cordic_tanangle_4_), .b(cordic_AngleCin), .o(cordic_Add0_MUX_0_n_22) );
NAND2_Z01 cordic_AddX_Add_g700 ( .a(cordic_AddX_Add_n_32), .b(cordic_AddX_Add_n_9), .o(cordic_AddX_Add_n_34) );
BUF_X2 newInst_249 ( .a(newNet_248), .o(newNet_249) );
BUF_X2 newInst_1032 ( .a(newNet_1031), .o(newNet_1032) );
XOR2_X1 cordic_AddX_g201 ( .a(cordic_AddX_Btemp_0_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_0_) );
BUF_X2 newInst_492 ( .a(newNet_491), .o(newNet_492) );
NAND2_Z01 g14945 ( .a(n_499), .b(n_575), .o(n_629) );
BUF_X2 newInst_1103 ( .a(newNet_1102), .o(newNet_1103) );
NAND2_Z01 cordic_SH1_srl_35_26_g1215 ( .a(cordic_iteration_0_), .b(cordic_Y_10_), .o(cordic_SH1_srl_35_26_n_37) );
BUF_X2 newInst_1014 ( .a(newNet_557), .o(newNet_1014) );
BUF_X2 newInst_430 ( .a(newNet_429), .o(newNet_430) );
BUF_X2 newInst_1056 ( .a(newNet_1055), .o(newNet_1056) );
BUF_X2 newInst_834 ( .a(newNet_829), .o(newNet_834) );
NAND2_Z01 cordic_SH2_srl_35_26_g1170 ( .a(cordic_SH2_srl_35_26_n_48), .b(cordic_iteration_1_), .o(cordic_SH2_srl_35_26_n_82) );
fflopd CoreInput_reg_4_ ( .CK(newNet_763), .D(n_645), .Q(CoreInput_4_) );
INV_X1 cordic_g488 ( .a(CoreOutput_23_), .o(cordic_n_19) );
BUF_X2 newInst_261 ( .a(newNet_260), .o(newNet_261) );
NAND2_Z01 g13496 ( .a(n_732), .b(n_755), .o(n_788) );
BUF_X2 newInst_334 ( .a(newNet_319), .o(newNet_334) );
NAND2_Z01 cordic_AddY_MUX_0_g310 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_12_), .o(cordic_AddY_MUX_0_n_11) );
XOR2_X1 cordic_AddX_Add_g713 ( .a(cordic_AddX_Btemp1_9_), .b(cordic_AddX_Atemp_9_), .o(cordic_AddX_Add_n_21) );
NOR2_Z1 g13453 ( .a(n_796), .b(n_710), .o(n_829) );
BUF_X2 newInst_1114 ( .a(newNet_1113), .o(newNet_1114) );
XNOR2_X1 cordic_AddX_Compl_g378 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_15_), .o(cordic_AddX_Compl_n_2) );
INV_X2 newInst_657 ( .a(newNet_656), .o(newNet_657) );
NAND2_Z01 cordic_SH2_srl_35_26_g1162 ( .a(cordic_SH2_srl_35_26_n_80), .b(cordic_SH2_srl_35_26_n_62), .o(cordic_SH2_srl_35_26_n_90) );
NAND2_Z01 cordic_AddX_MUX_0_g288 ( .a(cordic_AddX_MUX_0_n_17), .b(cordic_AddX_MUX_0_n_16), .o(cordic_AddX_Atemp_3_) );
BUF_X2 newInst_595 ( .a(newNet_594), .o(newNet_595) );
XOR2_X1 cordic_AddX_g209 ( .a(cordic_AddX_Btemp_3_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_3_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1244 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_6_), .o(cordic_SH1_srl_35_26_n_5) );
BUF_X2 newInst_873 ( .a(newNet_872), .o(newNet_873) );
BUF_X2 newInst_1065 ( .a(newNet_1064), .o(newNet_1065) );
BUF_X2 newInst_767 ( .a(newNet_766), .o(newNet_767) );
NAND2_Z01 cordic_AddY_Compl_g365 ( .a(cordic_AddY_Compl_n_11), .b(cordic_AddY_Compl_n_1), .o(cordic_AddY_Compl_n_17) );
INV_Z2 g13575 ( .a(Idsel), .o(n_712) );
NOR2_Z1 g13434 ( .a(n_814), .b(n_710), .o(n_848) );
AND3_X1 g15485 ( .a(n_44), .b(n_107), .c(OutputAvail), .o(n_178) );
XOR2_X1 g15322 ( .a(n_177), .b(n_168), .o(n_338) );
BUF_X2 newInst_900 ( .a(newNet_899), .o(newNet_900) );
NAND2_Z01 g14996 ( .a(n_572), .b(Config_Reg_14_), .o(n_581) );
BUF_X2 newInst_907 ( .a(newNet_906), .o(newNet_907) );
INV_X1 g15653 ( .a(Trdy_Wait_Cnt_2_), .o(n_12) );
BUF_X2 newInst_590 ( .a(newNet_249), .o(newNet_590) );
NAND2_Z01 cordic_SH2_srl_35_26_g1181 ( .a(cordic_SH2_srl_35_26_n_57), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_71) );
BUF_X2 newInst_774 ( .a(newNet_773), .o(newNet_774) );
NAND2_Z01 g14906 ( .a(n_615), .b(n_543), .o(n_668) );
fflopd OutputAvail_reg ( .CK(newNet_459), .D(n_578), .Q(OutputAvail) );
XOR2_X1 cordic_Add0_Compl_g340 ( .a(cordic_Add0_Compl_n_39), .b(cordic_Add0_Compl_n_8), .o(cordic_SumAngle_13_) );
INV_X1 drc_bufs15678 ( .a(n_188), .o(n_1) );
NAND2_Z01 cordic_Add0_Add_g672 ( .a(cordic_Add0_Add_n_33), .b(cordic_Add0_Add_n_2), .o(cordic_Add0_Add_n_35) );
BUF_X2 newInst_794 ( .a(newNet_793), .o(newNet_794) );
BUF_X2 newInst_396 ( .a(newNet_395), .o(newNet_396) );
fflopd Access_Type_1_reg_1_ ( .CK(newNet_1104), .D(n_468), .Q(Access_Type_1_1_) );
INV_X1 cordic_AddY_Compl_g382 ( .a(cordic_AddY_Y_4), .o(cordic_AddY_Compl_n_0) );
BUF_X2 newInst_1138 ( .a(newNet_1037), .o(newNet_1138) );
BUF_X2 newInst_246 ( .a(newNet_245), .o(newNet_246) );
NAND2_Z01 cordic_SH1_srl_35_26_g1169 ( .a(cordic_SH1_srl_35_26_n_44), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_83) );
NAND2_Z01 cordic_SH2_srl_35_26_g1241 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_3_), .o(cordic_SH2_srl_35_26_n_8) );
NAND2_Z01 g15623 ( .a(CoreCnt_En), .b(n_10), .o(n_44) );
BUF_X2 newInst_863 ( .a(newNet_862), .o(newNet_863) );
BUF_X2 newInst_337 ( .a(newNet_336), .o(newNet_337) );
XOR2_X1 cordic_AddX_Add_g709 ( .a(cordic_AddX_Btemp1_15_), .b(cordic_AddX_Atemp_15_), .o(cordic_AddX_Add_n_25) );
BUF_X2 newInst_678 ( .a(newNet_677), .o(newNet_678) );
BUF_X2 newInst_138 ( .a(newNet_137), .o(newNet_138) );
fflopd CoreOutputReg_reg_5_ ( .CK(newNet_5), .D(n_377), .Q(CoreOutputReg_5_) );
NAND2_Z01 g14967 ( .a(n_572), .b(Config_Reg_3_), .o(n_610) );
NAND2_Z01 cordic_Add0_MUX_1_g282 ( .a(cordic_AngleCin), .b(cordic_Angle_3_), .o(cordic_Add0_MUX_1_n_19) );
NAND2_Z01 cordic_AddY_Add_g700 ( .a(cordic_AddY_Add_n_32), .b(cordic_AddY_Add_n_9), .o(cordic_AddY_Add_n_34) );
BUF_X2 newInst_468 ( .a(newNet_64), .o(newNet_468) );
AND2_X1 g57 ( .a(n_823), .b(n_856), .o(PO_AD_7) );
NAND2_Z01 cordic_pla_g270 ( .a(cordic_pla_n_36), .b(cordic_pla_n_9), .o(cordic_tanangle_2_) );
BUF_X2 newInst_474 ( .a(newNet_473), .o(newNet_474) );
NOR2_Z1 cordic_SH2_srl_35_26_g1111 ( .a(cordic_SH2_srl_35_26_n_133), .b(cordic_iteration_3_), .o(cordic_BS2_8_) );
NAND2_Z01 g15373 ( .a(CoreOutput_22_), .b(n_188), .o(n_288) );
BUF_X2 newInst_802 ( .a(newNet_801), .o(newNet_802) );
BUF_X2 newInst_637 ( .a(newNet_636), .o(newNet_637) );
BUF_X2 newInst_365 ( .a(newNet_317), .o(newNet_365) );
NAND3_Z1 cordic_SH2_srl_35_26_g1115 ( .a(cordic_SH2_srl_35_26_n_115), .b(cordic_SH2_srl_35_26_n_118), .c(cordic_SH2_srl_35_26_n_59), .o(cordic_BS2_7_) );
NAND2_Z01 cordic_AddY_Add_g691 ( .a(cordic_AddY_Add_n_41), .b(cordic_AddY_Add_n_6), .o(cordic_AddY_Add_n_43) );
BUF_X2 newInst_245 ( .a(newNet_34), .o(newNet_245) );
NAND2_Z01 cordic_AddX_MUX_1_g291 ( .a(cordic_AddX_Y_1), .b(cordic_X_9_), .o(cordic_AddX_MUX_1_n_30) );
BUF_X2 newInst_661 ( .a(newNet_660), .o(newNet_661) );
NAND2_Z01 cordic_g412 ( .a(Issue_Rst), .b(CoreInput_12_), .o(cordic_n_95) );
BUF_X2 newInst_356 ( .a(newNet_355), .o(newNet_356) );
NAND2_Z01 cordic_g397 ( .a(cordic_n_68), .b(cordic_n_90), .o(cordic_n_110) );
BUF_X2 newInst_855 ( .a(newNet_854), .o(newNet_855) );
BUF_X2 newInst_541 ( .a(newNet_540), .o(newNet_541) );
BUF_X2 newInst_869 ( .a(newNet_868), .o(newNet_869) );
NAND2_Z01 cordic_g431 ( .a(cordic_Add0_Stemp_0_), .b(cordic_n_7), .o(cordic_n_76) );
BUF_X2 newInst_1205 ( .a(newNet_1139), .o(newNet_1205) );
NAND2_Z01 cordic_AddX_MUX_0_g273 ( .a(cordic_AddX_MUX_0_n_32), .b(cordic_AddX_MUX_0_n_7), .o(cordic_AddX_Atemp_15_) );
NAND2_Z01 cordic_AddX_MUX_1_g320 ( .a(cordic_BS1_10_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_1) );
NOR2_Z1 cordic_pla_g286 ( .a(cordic_pla_n_8), .b(cordic_iteration_1_), .o(cordic_pla_n_25) );
NAND2_Z01 cordic_g389 ( .a(cordic_n_74), .b(cordic_n_96), .o(cordic_n_118) );
XOR2_X1 cordic_AddX_Compl_g348 ( .a(cordic_AddX_Compl_n_31), .b(cordic_AddX_Compl_n_15), .o(CoreOutput_26_) );
INV_X1 g15639 ( .a(State_0_), .o(n_26) );
XOR2_X1 cordic_AddY_g197 ( .a(cordic_AddY_Btemp_15_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_15_) );
XOR2_X1 g15582 ( .a(PI_AD_14), .b(PI_AD_13), .o(n_83) );
BUF_X2 newInst_952 ( .a(newNet_951), .o(newNet_952) );
BUF_X2 newInst_103 ( .a(newNet_102), .o(newNet_103) );
INV_X1 g15473 ( .a(n_186), .o(n_185) );
fflopd TAR_TRI_S_reg ( .CK(newNet_340), .D(n_434), .Q(TAR_TRI_S) );
XOR2_X1 cordic_AddX_Add_g686 ( .a(cordic_AddX_Add_n_46), .b(cordic_AddX_Add_n_31), .o(cordic_AddX_Stemp_5_) );
NAND2_Z01 g14935 ( .a(n_586), .b(n_515), .o(n_639) );
NOR2_Z1 cordic_g455 ( .a(cordic_n_11), .b(Issue_Rst), .o(cordic_n_52) );
NAND2_Z01 g14954 ( .a(n_572), .b(Config_Reg_20_), .o(n_623) );
INV_X1 cordic_AddX_g36 ( .a(cordic_Xsign), .o(cordic_AddX_n_5) );
NAND2_Z01 cordic_Add0_Add_g694 ( .a(cordic_Add0_n_6), .b(cordic_Add0_Atemp_5_), .o(cordic_Add0_Add_n_13) );
BUF_X2 newInst_731 ( .a(newNet_730), .o(newNet_731) );
BUF_X2 newInst_159 ( .a(newNet_158), .o(newNet_159) );
NOR2_Z1 g13463 ( .a(n_784), .b(n_710), .o(n_819) );
NAND2_Z01 cordic_SH2_srl_35_26_g1126 ( .a(cordic_SH2_srl_35_26_n_119), .b(cordic_SH2_srl_35_26_n_60), .o(cordic_SH2_srl_35_26_n_126) );
fflopd State_reg_0_ ( .CK(newNet_387), .D(n_498), .Q(State_0_) );
NAND2_Z01 cordic_AddX_Add_g678 ( .a(cordic_AddX_Add_n_55), .b(cordic_AddX_Add_n_17), .o(cordic_AddX_Add_n_56) );
NAND2_Z01 cordic_AddX_MUX_0_g300 ( .a(cordic_BS1_5_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_21) );
BUF_X2 newInst_58 ( .a(newNet_34), .o(newNet_58) );
BUF_X2 newInst_43 ( .a(newNet_42), .o(newNet_43) );
BUF_X2 newInst_1159 ( .a(newNet_1158), .o(newNet_1159) );
BUF_X2 newInst_579 ( .a(newNet_578), .o(newNet_579) );
NAND2_Z01 cordic_AddY_Add_g720 ( .a(cordic_AddY_Btemp1_11_), .b(cordic_AddY_Atemp_11_), .o(cordic_AddY_Add_n_14) );
BUF_X2 newInst_622 ( .a(newNet_506), .o(newNet_622) );
INV_X1 cordic_g499 ( .a(CoreOutput_13_), .o(cordic_n_8) );
XOR2_X1 g15022 ( .a(n_452), .b(n_451), .o(n_560) );
XOR2_X1 cordic_AddY_Add_g662 ( .a(cordic_AddY_Add_n_70), .b(cordic_AddY_Add_n_23), .o(cordic_AddY_Stemp_13_) );
BUF_X2 newInst_854 ( .a(newNet_853), .o(newNet_854) );
BUF_X2 newInst_823 ( .a(newNet_663), .o(newNet_823) );
BUF_X2 newInst_662 ( .a(newNet_661), .o(newNet_662) );
BUF_X2 newInst_498 ( .a(newNet_497), .o(newNet_498) );
NOR2_Z1 g13458 ( .a(n_809), .b(n_710), .o(n_824) );
NAND2_Z01 cordic_AddY_Add_g679 ( .a(cordic_AddY_Add_n_53), .b(cordic_AddY_Add_n_15), .o(cordic_AddY_Add_n_55) );
BUF_X2 newInst_1015 ( .a(newNet_1014), .o(newNet_1015) );
BUF_X2 newInst_858 ( .a(newNet_857), .o(newNet_858) );
BUF_X2 newInst_221 ( .a(newNet_220), .o(newNet_221) );
XOR2_X1 g13402 ( .a(n_877), .b(PO_AD_23), .o(n_878) );
NAND2_Z01 cordic_AddY_MUX_1_g274 ( .a(cordic_AddY_MUX_1_n_11), .b(cordic_AddY_MUX_1_n_28), .o(cordic_AddY_Btemp_12_) );
AND2_X1 g358 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_36) );
BUF_X2 newInst_13 ( .a(newNet_12), .o(newNet_13) );
NOR2_Z1 cordic_g352 ( .a(cordic_n_100), .b(Issue_Rst), .o(cordic_n_120) );
INV_X1 cordic_g485 ( .a(CoreOutput_31_), .o(cordic_n_22) );
NOR2_Z1 g15434 ( .a(n_165), .b(n_44), .o(n_224) );
NAND2_Z01 g14916 ( .a(n_605), .b(n_534), .o(n_658) );
BUF_X2 newInst_642 ( .a(newNet_641), .o(newNet_642) );
NAND2_Z01 g13522 ( .a(Idsel), .b(Config_Reg_13_), .o(n_764) );
BUF_X2 newInst_296 ( .a(newNet_295), .o(newNet_296) );
NAND2_Z01 g15094 ( .a(n_464), .b(Issue_Rst), .o(n_514) );
NOR2_Z1 g13443 ( .a(n_804), .b(n_710), .o(n_839) );
NOR2_Z1 cordic_g462 ( .a(cordic_n_2), .b(Issue_Rst), .o(cordic_n_45) );
BUF_X2 newInst_889 ( .a(newNet_888), .o(newNet_889) );
BUF_X2 newInst_466 ( .a(newNet_465), .o(newNet_466) );
fflopd Config_Reg_reg_7_ ( .CK(newNet_859), .D(n_659), .Q(Config_Reg_7_) );
XOR2_X1 cordic_AddX_Add_g674 ( .a(cordic_AddX_Add_n_58), .b(cordic_AddX_Add_n_21), .o(cordic_AddX_Stemp_9_) );
XOR2_X1 cordic_AddY_Add_g665 ( .a(cordic_AddY_Add_n_67), .b(cordic_AddY_Add_n_19), .o(cordic_AddY_Stemp_12_) );
AND2_X1 cordic_Add0_Compl_g349 ( .a(cordic_Add0_Compl_n_31), .b(cordic_Add0_Compl_n_15), .o(cordic_Add0_Compl_n_33) );
INV_X1 g15644 ( .a(Access_Address_1_26_), .o(n_21) );
fflopd Config_Reg_reg_8_ ( .CK(newNet_856), .D(n_658), .Q(Config_Reg_8_) );
AND2_X1 cordic_AddY_Compl_g357 ( .a(cordic_AddY_Compl_n_23), .b(cordic_AddY_Compl_n_5), .o(cordic_AddY_Compl_n_25) );
XOR2_X1 cordic_AddY_Add_g686 ( .a(cordic_AddY_Add_n_46), .b(cordic_AddY_Add_n_31), .o(cordic_AddY_Stemp_5_) );
NAND2_Z01 g15261 ( .a(n_288), .b(n_289), .o(n_399) );
fflopd TAR_TRI_T_reg ( .CK(newNet_333), .D(n_453), .Q(TAR_TRI_T) );
NAND2_Z01 cordic_AddX_MUX_1_g278 ( .a(cordic_AddX_MUX_1_n_13), .b(cordic_AddX_MUX_1_n_27), .o(cordic_AddX_Btemp_1_) );
BUF_X2 newInst_413 ( .a(newNet_412), .o(newNet_413) );
NAND2_Z01 g13531 ( .a(Idsel), .b(Config_Reg_8_), .o(n_755) );
BUF_X2 newInst_283 ( .a(newNet_282), .o(newNet_283) );
NAND2_Z01 g15084 ( .a(n_4), .b(PI_AD_2), .o(n_524) );
NAND2_Z01 g13541 ( .a(n_712), .b(CoreOutputReg_31_), .o(n_745) );
NAND2_Z01 cordic_Add0_MUX_1_g266 ( .a(cordic_Add0_MUX_1_n_15), .b(cordic_Add0_MUX_1_n_31), .o(cordic_Add0_Btemp_8_) );
BUF_X2 newInst_1003 ( .a(newNet_1002), .o(newNet_1003) );
NAND2_Z01 cordic_Add0_Add_g696 ( .a(cordic_Add0_n_7), .b(cordic_Add0_Atemp_6_), .o(cordic_Add0_Add_n_11) );
NAND4_Z1 g15217 ( .a(n_134), .b(n_206), .c(n_216), .d(n_155), .o(n_436) );
XOR2_X1 g15497 ( .a(n_90), .b(n_89), .o(n_166) );
AND2_X1 g15452 ( .a(n_149), .b(n_967), .o(n_203) );
XOR2_X1 cordic_AddY_g208 ( .a(cordic_AddY_Btemp_4_), .b(cordic_AddY_Y_2), .o(cordic_AddY_Btemp1_4_) );
AND2_X1 cordic_AddY_Compl_g361 ( .a(cordic_AddY_Compl_n_19), .b(cordic_AddY_Compl_n_16), .o(cordic_AddY_Compl_n_21) );
NAND2_Z01 g13499 ( .a(n_718), .b(n_750), .o(n_785) );
INV_X1 g15527 ( .a(n_129), .o(n_128) );
NAND3_Z1 g15539 ( .a(Access_Type_1_3_), .b(n_36), .c(Access_Type_1_0_), .o(n_132) );
NAND2_Z01 cordic_Add0_Add_g657 ( .a(cordic_Add0_Add_n_48), .b(cordic_Add0_Add_n_11), .o(cordic_Add0_Add_n_50) );
AND2_X1 g49 ( .a(n_835), .b(n_856), .o(PO_AD_15) );
fflopd Config_Reg_reg_19_ ( .CK(newNet_985), .D(n_678), .Q(Config_Reg_19_) );
BUF_X2 newInst_480 ( .a(newNet_479), .o(newNet_480) );
BUF_X2 newInst_1120 ( .a(newNet_1119), .o(newNet_1120) );
XOR2_X1 cordic_Add0_Compl_g354 ( .a(cordic_Add0_Compl_n_25), .b(cordic_Add0_Compl_n_4), .o(cordic_SumAngle_6_) );
INV_Z1 cordic_Add0_g53 ( .a(cordic_Add0_Btemp_8_), .o(cordic_Add0_n_9) );
BUF_X2 newInst_313 ( .a(newNet_312), .o(newNet_313) );
NAND2_Z01 g15277 ( .a(n_246), .b(n_247), .o(n_378) );
fflopd CoreInput_reg_7_ ( .CK(newNet_743), .D(n_642), .Q(CoreInput_7_) );
fflopd Config_Reg_reg_13_ ( .CK(newNet_1028), .D(n_635), .Q(Config_Reg_13_) );
BUF_X2 newInst_1020 ( .a(newNet_137), .o(newNet_1020) );
INV_X1 cordic_SH2_srl_35_26_g1204 ( .a(cordic_SH2_srl_35_26_n_41), .o(cordic_SH2_srl_35_26_n_40) );
NAND2_Z01 g13493 ( .a(n_725), .b(n_758), .o(n_791) );
NAND2_Z01 g15279 ( .a(n_243), .b(n_244), .o(n_376) );
BUF_X2 newInst_764 ( .a(newNet_159), .o(newNet_764) );
INV_X1 g15612 ( .a(n_52), .o(n_53) );
BUF_X2 newInst_599 ( .a(newNet_408), .o(newNet_599) );
NAND2_Z01 g15061 ( .a(n_473), .b(PI_AD_25), .o(n_547) );
fflopd Config_Reg_reg_16_ ( .CK(newNet_1003), .D(n_632), .Q(Config_Reg_16_) );
NAND2_Z01 cordic_AddX_MUX_0_g299 ( .a(cordic_BS1_6_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_22) );
fflopd cordic_Y_reg_11_ ( .CK(newNet_89), .D(cordic_n_45), .Q(cordic_Y_11_) );
BUF_X2 newInst_24 ( .a(newNet_23), .o(newNet_24) );
NAND2_Z01 cordic_SH1_srl_35_26_g1206 ( .a(cordic_SH1_srl_35_26_n_5), .b(cordic_SH1_srl_35_26_n_27), .o(cordic_SH1_srl_35_26_n_47) );
BUF_X2 newInst_1084 ( .a(newNet_1083), .o(newNet_1084) );
BUF_X1 mybuffer1 ( .a(cordic_AngleCout), .o(PO_ACK64_L) );
NAND2_Z01 cordic_SH2_srl_35_26_g1176 ( .a(cordic_SH2_srl_35_26_n_43), .b(cordic_SH2_srl_35_26_n_52), .o(cordic_SH2_srl_35_26_n_76) );
NAND2_Z01 cordic_AddY_MUX_0_g290 ( .a(cordic_BS2_14_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_31) );
NAND2_Z01 g15333 ( .a(n_184), .b(PI_AD_24), .o(n_328) );
XNOR2_X1 cordic_AddX_Compl_g369 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_14_), .o(cordic_AddX_Compl_n_13) );
NAND2_Z01 cordic_pla_g276 ( .a(cordic_pla_n_22), .b(cordic_pla_n_16), .o(cordic_tanangle_7_) );
NAND2_Z01 cordic_Add0_Add_g665 ( .a(cordic_Add0_Add_n_41), .b(cordic_Add0_Add_n_25), .o(cordic_Add0_Add_n_42) );
NAND2_Z01 g14943 ( .a(n_506), .b(n_576), .o(n_631) );
NAND2_Z01 cordic_SH2_srl_35_26_g1158 ( .a(cordic_SH2_srl_35_26_n_81), .b(cordic_SH2_srl_35_26_n_64), .o(cordic_SH2_srl_35_26_n_95) );
NAND2_Z01 g15396 ( .a(CoreOutput_30_), .b(n_2), .o(n_254) );
BUF_X2 newInst_517 ( .a(newNet_516), .o(newNet_517) );
BUF_X2 newInst_449 ( .a(newNet_448), .o(newNet_449) );
NAND2_Z01 cordic_SH1_srl_35_26_g1133 ( .a(cordic_SH1_srl_35_26_n_98), .b(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_119) );
NAND4_Z1 cordic_SH1_srl_35_26_g1106 ( .a(cordic_SH1_srl_35_26_n_70), .b(cordic_SH1_srl_35_26_n_116), .c(cordic_SH1_srl_35_26_n_143), .d(cordic_SH1_srl_35_26_n_72), .o(cordic_BS1_0_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1234 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_1_), .o(cordic_SH2_srl_35_26_n_15) );
INV_X2 newInst_1174 ( .a(newNet_1173), .o(newNet_1174) );
INV_X1 g15550 ( .a(n_108), .o(n_107) );
NAND2_Z01 cordic_AddY_MUX_1_g299 ( .a(cordic_AddY_Y_1), .b(cordic_Y_6_), .o(cordic_AddY_MUX_1_n_22) );
NAND2_Z01 cordic_AddY_MUX_0_g297 ( .a(cordic_BS2_7_), .b(cordic_AddY_Y_1), .o(cordic_AddY_MUX_0_n_24) );
NAND2_Z01 g15404 ( .a(CoreOutput_4_), .b(n_2), .o(n_246) );
NOR2_Z1 cordic_g427 ( .a(cordic_n_25), .b(Issue_Rst), .o(cordic_n_80) );
NAND2_Z01 cordic_Add0_MUX_1_g291 ( .a(cordic_tanangle_7_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_10) );
XOR2_X1 cordic_AddY_Add_g712 ( .a(cordic_AddY_Btemp1_14_), .b(cordic_AddY_Atemp_14_), .o(cordic_AddY_Add_n_22) );
NAND2_Z01 g13568 ( .a(n_712), .b(CoreOutputReg_23_), .o(n_719) );
fflopd DWord_Trans_reg ( .CK(newNet_521), .D(n_516), .Q(DWord_Trans) );
XOR2_X1 cordic_AddY_Add_g711 ( .a(cordic_AddY_Btemp1_13_), .b(cordic_AddY_Atemp_13_), .o(cordic_AddY_Add_n_23) );
BUF_X2 newInst_809 ( .a(newNet_808), .o(newNet_809) );
XOR2_X1 g13421 ( .a(n_858), .b(CBE_par_2_), .o(n_860) );
BUF_X2 newInst_1052 ( .a(newNet_1051), .o(newNet_1052) );
BUF_X2 newInst_1008 ( .a(newNet_1007), .o(newNet_1008) );
NAND2_Z01 cordic_SH1_srl_35_26_g1183 ( .a(cordic_SH1_srl_35_26_n_48), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_69) );
XOR2_X1 cordic_Add0_Compl_g352 ( .a(cordic_Add0_Compl_n_27), .b(cordic_Add0_Compl_n_6), .o(cordic_SumAngle_7_) );
NAND2_Z01 g13553 ( .a(n_897), .b(Access_Type_1_1_), .o(n_973) );
fflopd Trdy_Wait_Cnt_reg_1_ ( .CK(newNet_313), .D(n_230), .Q(Trdy_Wait_Cnt_1_) );
BUF_X2 newInst_96 ( .a(newNet_95), .o(newNet_96) );
XOR2_X1 cordic_AddX_g198 ( .a(cordic_AddX_Btemp_14_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_14_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1185 ( .a(cordic_SH2_srl_35_26_n_50), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_67) );
BUF_X2 newInst_915 ( .a(newNet_914), .o(newNet_915) );
NOR2_Z1 cordic_Add0_Compl_g381 ( .a(cordic_Add0_Compl_n_0), .b(cordic_Add0_Stemp_0_), .o(cordic_Add0_Compl_n_1) );
NAND2_Z01 cordic_AddX_Add_g696 ( .a(cordic_AddX_Add_n_37), .b(cordic_AddX_Add_n_20), .o(cordic_AddX_Add_n_38) );
BUF_X2 newInst_648 ( .a(newNet_647), .o(newNet_648) );
NAND2_Z01 cordic_SH2_srl_35_26_g1140 ( .a(cordic_SH2_srl_35_26_n_93), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_112) );
NAND2_Z01 cordic_AddY_MUX_1_g289 ( .a(cordic_AddY_Y_1), .b(cordic_Y_15_), .o(cordic_AddY_MUX_1_n_32) );
BUF_X2 newInst_132 ( .a(newNet_131), .o(newNet_132) );
BUF_X2 newInst_1163 ( .a(newNet_1162), .o(newNet_1163) );
XOR2_X1 g15601 ( .a(PI_CBE_L_6), .b(PI_CBE_L_5), .o(n_64) );
NAND2_Z01 cordic_AddX_Add_g723 ( .a(cordic_AddX_Btemp1_5_), .b(cordic_AddX_Atemp_5_), .o(cordic_AddX_Add_n_11) );
XOR2_X1 g13388 ( .a(n_891), .b(PO_AD_13), .o(n_892) );
AND2_X1 cordic_AddY_Compl_g341 ( .a(cordic_AddY_Compl_n_39), .b(cordic_AddY_Compl_n_8), .o(cordic_AddY_Compl_n_41) );
INV_X1 cordic_SH1_srl_35_26_g1121 ( .a(cordic_SH1_srl_35_26_n_130), .o(cordic_SH1_srl_35_26_n_131) );
BUF_X2 newInst_722 ( .a(newNet_721), .o(newNet_722) );
XOR2_X1 cordic_AddY_Compl_g338 ( .a(cordic_AddY_Compl_n_41), .b(cordic_AddY_Compl_n_13), .o(CoreOutput_14_) );
NAND2_Z01 cordic_AddX_MUX_1_g285 ( .a(cordic_AddX_MUX_1_n_1), .b(cordic_AddX_MUX_1_n_19), .o(cordic_AddX_Btemp_10_) );
NAND2_Z01 g15066 ( .a(n_473), .b(PI_AD_29), .o(n_542) );
NAND2_Z01 cordic_Add0_MUX_1_g277 ( .a(cordic_AngleCin), .b(cordic_Angle_5_), .o(cordic_Add0_MUX_1_n_24) );
BUF_X2 newInst_1011 ( .a(newNet_1010), .o(newNet_1011) );
BUF_X2 newInst_880 ( .a(newNet_879), .o(newNet_880) );
fflopd cordic_Angle_reg_15_ ( .CK(newNet_244), .D(cordic_n_111), .Q(cordic_Angle_15_) );
INV_Z1 cordic_Add0_g50 ( .a(cordic_Add0_Btemp_11_), .o(cordic_Add0_n_12) );
NAND2_Z01 g14826 ( .a(n_692), .b(n_10), .o(n_694) );
BUF_X2 newInst_25 ( .a(newNet_0), .o(newNet_25) );
BUF_X2 newInst_444 ( .a(newNet_443), .o(newNet_444) );
NAND3_Z1 g14815 ( .a(n_6), .b(n_696), .c(n_187), .o(n_704) );
NAND2_Z01 cordic_SH1_srl_35_26_g1187 ( .a(cordic_SH1_srl_35_26_n_54), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_65) );
fflopd cordic_X_reg_6_ ( .CK(newNet_117), .D(cordic_n_48), .Q(cordic_X_6_) );
NAND2_Z01 cordic_Add0_Add_g701 ( .a(cordic_Add0_n_4), .b(cordic_Add0_Atemp_3_), .o(cordic_Add0_Add_n_6) );
NAND2_Z01 cordic_AddY_MUX_1_g320 ( .a(cordic_BS2_10_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_1) );
NAND2_Z01 g15391 ( .a(n_214), .b(CoreOutputReg_29_), .o(n_259) );
BUF_X2 newInst_618 ( .a(newNet_617), .o(newNet_618) );
BUF_X2 newInst_980 ( .a(newNet_979), .o(newNet_980) );
NOR2_Z1 cordic_pla_g282 ( .a(cordic_pla_n_4), .b(cordic_pla_n_2), .o(cordic_pla_n_28) );
XOR2_X1 g13393 ( .a(n_886), .b(PO_AD_1), .o(n_887) );
BUF_X2 newInst_1183 ( .a(newNet_1182), .o(newNet_1183) );
BUF_X2 newInst_1135 ( .a(newNet_1134), .o(newNet_1135) );
BUF_X2 newInst_371 ( .a(newNet_370), .o(newNet_371) );
NAND2_Z01 g15625 ( .a(Set_Data_Parity), .b(n_10), .o(n_40) );
NAND2_Z01 cordic_AddX_MUX_1_g313 ( .a(cordic_BS1_7_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_8) );
NAND2_Z01 g15280 ( .a(n_241), .b(n_242), .o(n_375) );
BUF_X2 newInst_427 ( .a(newNet_426), .o(newNet_427) );
XOR2_X1 g15491 ( .a(n_74), .b(n_75), .o(n_172) );
NAND2_Z01 cordic_Add0_Add_g632 ( .a(cordic_Add0_Add_n_74), .b(cordic_Add0_Add_n_24), .o(cordic_Add0_Add_n_75) );
NAND2_Z01 cordic_Add0_MUX_1_g287 ( .a(cordic_tanangle_1_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_14) );
NAND2_Z01 cordic_SH1_srl_35_26_g1154 ( .a(cordic_SH1_srl_35_26_n_87), .b(cordic_SH1_srl_35_26_n_75), .o(cordic_SH1_srl_35_26_n_99) );
BUF_X2 newInst_1083 ( .a(newNet_1082), .o(newNet_1083) );
BUF_X2 newInst_496 ( .a(newNet_495), .o(newNet_496) );
fflopd CoreOutputReg_reg_15_ ( .CK(newNet_701), .D(n_408), .Q(CoreOutputReg_15_) );
BUF_X2 newInst_684 ( .a(newNet_487), .o(newNet_684) );
BUF_X2 newInst_87 ( .a(newNet_35), .o(newNet_87) );
NAND2_Z01 g15407 ( .a(CoreOutput_6_), .b(n_188), .o(n_243) );
XOR2_X1 g15574 ( .a(Trdy_Wait_Cnt_0_), .b(Trdy_Wait_Cnt_1_), .o(n_91) );
BUF_X2 newInst_782 ( .a(newNet_781), .o(newNet_782) );
NAND2_Z01 g14973 ( .a(n_572), .b(Config_Reg_9_), .o(n_604) );
INV_X1 cordic_g502 ( .a(CoreOutput_4_), .o(cordic_n_5) );
NAND3_Z1 g15158 ( .a(n_354), .b(n_355), .c(n_109), .o(n_454) );
NAND2_Z01 cordic_g424 ( .a(Issue_Rst), .b(CoreInput_9_), .o(cordic_n_83) );
NAND2_Z02 g15226 ( .a(n_348), .b(n_127), .o(n_445) );
NAND2_Z01 cordic_AddY_MUX_0_g277 ( .a(cordic_AddY_MUX_0_n_26), .b(cordic_AddY_MUX_0_n_10), .o(cordic_AddY_Atemp_8_) );
BUF_X2 newInst_193 ( .a(newNet_192), .o(newNet_193) );
NAND2_Z01 cordic_AddX_MUX_1_g279 ( .a(cordic_AddX_MUX_1_n_12), .b(cordic_AddX_MUX_1_n_25), .o(cordic_AddX_Btemp_0_) );
NAND2_Z01 cordic_SH2_srl_35_26_g1244 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_6_), .o(cordic_SH2_srl_35_26_n_5) );
BUF_X2 newInst_175 ( .a(newNet_174), .o(newNet_175) );
BUF_X2 newInst_238 ( .a(newNet_153), .o(newNet_238) );
BUF_X2 newInst_311 ( .a(newNet_278), .o(newNet_311) );
NOR4_Z1 g13427 ( .a(n_22), .b(n_798), .c(n_799), .d(PI_IRDY_L), .o(n_855) );
NAND2_Z01 cordic_SH1_srl_35_26_g1239 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_11_), .o(cordic_SH1_srl_35_26_n_10) );
NAND2_Z01 cordic_AddY_MUX_1_g296 ( .a(cordic_AddY_Y_1), .b(cordic_Y_0_), .o(cordic_AddY_MUX_1_n_25) );
AND2_X1 cordic_g477 ( .a(CoreOutput_25_), .b(Issue_Rst), .o(cordic_n_30) );
XNOR2_X1 cordic_AddX_g2 ( .a(cordic_n_144), .b(cordic_Xsign), .o(cordic_AddX_n_0) );
NAND2_Z01 g13550 ( .a(n_712), .b(CoreOutputReg_19_), .o(n_736) );
BUF_X2 newInst_692 ( .a(newNet_691), .o(newNet_692) );
NAND2_Z01 g15337 ( .a(CoreOutput_5_), .b(n_2), .o(n_324) );
NAND2_Z01 cordic_g440 ( .a(cordic_SumAngle_2_), .b(cordic_n_7), .o(cordic_n_67) );
BUF_X2 newInst_206 ( .a(newNet_100), .o(newNet_206) );
BUF_X2 newInst_172 ( .a(newNet_171), .o(newNet_172) );
INV_X1 g15525 ( .a(n_137), .o(n_136) );
BUF_X2 newInst_969 ( .a(newNet_968), .o(newNet_969) );
BUF_X2 newInst_626 ( .a(newNet_625), .o(newNet_626) );
NAND2_Z01 g13511 ( .a(Idsel), .b(Config_Reg_30_), .o(n_775) );
AND2_X1 g343 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_51) );
NAND2_Z01 cordic_Add0_MUX_0_g265 ( .a(cordic_Add0_MUX_0_n_25), .b(cordic_Add0_MUX_0_n_8), .o(cordic_Add0_Atemp_5_) );
BUF_X2 newInst_624 ( .a(newNet_359), .o(newNet_624) );
BUF_X2 newInst_559 ( .a(newNet_558), .o(newNet_559) );
BUF_X2 newInst_650 ( .a(newNet_649), .o(newNet_650) );
NAND2_Z01 cordic_SH1_srl_35_26_g1232 ( .a(cordic_SH1_srl_35_26_n_0), .b(cordic_Y_2_), .o(cordic_SH1_srl_35_26_n_17) );
NAND2_Z01 cordic_AddX_Add_g730 ( .a(cordic_AddX_Btemp1_12_), .b(cordic_AddX_Atemp_12_), .o(cordic_AddX_Add_n_4) );
BUF_X2 newInst_290 ( .a(newNet_289), .o(newNet_290) );
NAND2_Z01 g14980 ( .a(n_571), .b(CoreInput_15_), .o(n_597) );
BUF_X2 newInst_34 ( .a(newNet_15), .o(newNet_34) );
fflopd CoreOutputReg_reg_8_ ( .CK(newNet_555), .D(n_374), .Q(CoreOutputReg_8_) );
NAND2_Z01 g15054 ( .a(n_473), .b(PI_AD_19), .o(n_554) );
INV_X1 cordic_g496 ( .a(CoreOutput_20_), .o(cordic_n_11) );
AND2_X1 g15466 ( .a(n_134), .b(n_8), .o(n_212) );
XOR2_X1 g15589 ( .a(PI_AD_24), .b(PI_AD_17), .o(n_76) );
BUF_X2 newInst_330 ( .a(newNet_163), .o(newNet_330) );
INV_X1 g15650 ( .a(TAR_TRI_E), .o(n_15) );
AND2_X1 cordic_Add0_Compl_g339 ( .a(cordic_Add0_Compl_n_41), .b(cordic_Add0_Compl_n_13), .o(cordic_Add0_Compl_n_43) );
NOR2_Z1 g15126 ( .a(n_445), .b(n_217), .o(n_497) );
XNOR2_X1 cordic_AddX_Compl_g377 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_5_), .o(cordic_AddX_Compl_n_5) );
XOR2_X1 g13407 ( .a(n_872), .b(PO_AD_7), .o(n_873) );
fflopd Access_Address_1_reg_20_ ( .CK(newNet_1180), .D(n_482), .Q(Access_Address_1_20_) );
BUF_X2 newInst_276 ( .a(newNet_275), .o(newNet_276) );
fflopd Trdy_Cnt_En_reg ( .CK(newNet_329), .D(n_708), .Q(Trdy_Cnt_En) );
NAND2_Z01 g14912 ( .a(n_611), .b(n_539), .o(n_662) );
NAND2_Z01 cordic_SH1_srl_35_26_g1185 ( .a(cordic_SH1_srl_35_26_n_50), .b(cordic_SH1_srl_35_26_n_3), .o(cordic_SH1_srl_35_26_n_67) );
BUF_X2 newInst_1198 ( .a(newNet_1197), .o(newNet_1198) );
BUF_X2 newInst_212 ( .a(newNet_211), .o(newNet_212) );
XOR2_X1 cordic_AddX_g197 ( .a(cordic_AddX_Btemp_15_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_15_) );
NAND2_Z01 g13527 ( .a(Idsel), .b(Config_Reg_10_), .o(n_759) );
NAND2_Z01 cordic_SH1_srl_35_26_g1178 ( .a(cordic_SH1_srl_35_26_n_42), .b(cordic_SH1_srl_35_26_n_53), .o(cordic_SH1_srl_35_26_n_74) );
BUF_X2 newInst_351 ( .a(newNet_350), .o(newNet_351) );
fflopd CBE_par_reg_0_ ( .CK(newNet_1091), .D(n_352), .Q(CBE_par_0_) );
NAND2_Z01 g15080 ( .a(n_473), .b(PI_AD_5), .o(n_528) );
BUF_X2 newInst_832 ( .a(newNet_831), .o(newNet_832) );
NAND2_Z01 g15386 ( .a(CoreOutput_26_), .b(n_188), .o(n_264) );
NAND2_Z01 cordic_SH1_srl_35_26_g1196 ( .a(cordic_SH1_srl_35_26_n_12), .b(cordic_SH1_srl_35_26_n_37), .o(cordic_SH1_srl_35_26_n_56) );
NOR2_Z1 cordic_g465 ( .a(cordic_n_0), .b(Issue_Rst), .o(cordic_n_42) );
BUF_X2 newInst_957 ( .a(newNet_956), .o(newNet_957) );
BUF_X2 newInst_726 ( .a(newNet_725), .o(newNet_726) );
NAND2_Z01 g15087 ( .a(n_494), .b(PI_AD_5), .o(n_521) );
BUF_X2 newInst_1044 ( .a(newNet_1043), .o(newNet_1044) );
BUF_X2 newInst_904 ( .a(newNet_903), .o(newNet_904) );
BUF_X2 newInst_348 ( .a(newNet_347), .o(newNet_348) );
BUF_X2 newInst_184 ( .a(newNet_183), .o(newNet_184) );
NAND2_Z01 g13525 ( .a(Idsel), .b(Config_Reg_15_), .o(n_761) );
NAND3_Z1 g15127 ( .a(n_321), .b(n_421), .c(n_10), .o(n_483) );
NAND2_Z01 cordic_g445 ( .a(cordic_SumAngle_7_), .b(cordic_n_7), .o(cordic_n_62) );
BUF_X2 newInst_641 ( .a(newNet_482), .o(newNet_641) );
BUF_X2 newInst_376 ( .a(newNet_375), .o(newNet_376) );
NAND2_Z01 cordic_Add0_MUX_0_g294 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_3_), .o(cordic_Add0_MUX_0_n_9) );
XNOR2_X1 cordic_AddX_Compl_g370 ( .a(cordic_AddX_Y_4), .b(cordic_AddX_Stemp_12_), .o(cordic_AddX_Compl_n_12) );
BUF_X2 newInst_470 ( .a(newNet_469), .o(newNet_470) );
fflopd cordic_X_reg_15_ ( .CK(newNet_33), .D(cordic_n_32), .Q(cordic_X_15_) );
NAND2_Z01 g15353 ( .a(CoreOutput_14_), .b(n_188), .o(n_308) );
BUF_X2 newInst_1075 ( .a(newNet_1074), .o(newNet_1075) );
BUF_X2 newInst_502 ( .a(newNet_501), .o(newNet_502) );
INV_X1 cordic_pla_g310 ( .a(cordic_iteration_3_), .o(cordic_pla_n_1) );
BUF_X2 newInst_5 ( .a(newNet_4), .o(newNet_5) );
NAND2_Z01 cordic_AddX_Add_g667 ( .a(cordic_AddX_Add_n_65), .b(cordic_AddX_Add_n_14), .o(cordic_AddX_Add_n_67) );
fflopd DevSel_Cnt_En_reg ( .CK(newNet_517), .D(n_438), .Q(DevSel_Cnt_En) );
XOR2_X1 cordic_AddX_Add_g704 ( .a(cordic_AddX_Btemp1_7_), .b(cordic_AddX_Atemp_7_), .o(cordic_AddX_Add_n_30) );
NOR2_Z1 cordic_SH1_srl_35_26_g1111 ( .a(cordic_SH1_srl_35_26_n_133), .b(cordic_iteration_3_), .o(cordic_BS1_8_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1198 ( .a(cordic_SH1_srl_35_26_n_13), .b(cordic_SH1_srl_35_26_n_26), .o(cordic_SH1_srl_35_26_n_54) );
NAND2_Z01 cordic_AddY_MUX_0_g308 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_1_), .o(cordic_AddY_MUX_0_n_13) );
XOR2_X1 cordic_Add0_Compl_g371 ( .a(cordic_AngleCout), .b(cordic_Add0_Stemp_1_), .o(cordic_Add0_Compl_n_11) );
NAND2_Z01 g14976 ( .a(n_571), .b(CoreInput_11_), .o(n_601) );
INV_X1 cordic_pla_g303 ( .a(cordic_pla_n_8), .o(cordic_pla_n_7) );
BUF_X2 newInst_1177 ( .a(newNet_1176), .o(newNet_1177) );
BUF_X2 newInst_851 ( .a(newNet_850), .o(newNet_851) );
NAND2_Z01 g13570 ( .a(n_712), .b(CoreOutputReg_26_), .o(n_717) );
BUF_X2 newInst_1129 ( .a(newNet_1128), .o(newNet_1129) );
AND2_X1 cordic_Add0_Compl_g363 ( .a(cordic_Add0_Compl_n_17), .b(cordic_Add0_Compl_n_14), .o(cordic_Add0_Compl_n_19) );
fflopd cordic_Angle_reg_13_ ( .CK(newNet_252), .D(cordic_n_113), .Q(cordic_Angle_13_) );
AND2_X1 g13571 ( .a(PAR_Int), .b(RESET), .o(n_716) );
XOR2_X1 cordic_AddY_Compl_g352 ( .a(cordic_AddY_Compl_n_27), .b(cordic_AddY_Compl_n_6), .o(CoreOutput_7_) );
NAND2_Z01 g15150 ( .a(n_444), .b(n_277), .o(n_462) );
XOR2_X1 g13418 ( .a(n_861), .b(CBE_par_0_), .o(n_862) );
NAND2_Z01 g14904 ( .a(n_617), .b(n_545), .o(n_670) );
BUF_X2 newInst_418 ( .a(newNet_417), .o(newNet_418) );
BUF_X2 newInst_943 ( .a(newNet_942), .o(newNet_943) );
NOR2_Z1 cordic_AddY_Compl_g381 ( .a(cordic_AddY_Compl_n_0), .b(cordic_AddY_Stemp_0_), .o(cordic_AddY_Compl_n_1) );
NAND2_Z01 cordic_AddX_MUX_0_g290 ( .a(cordic_BS1_14_), .b(cordic_AddX_Y_1), .o(cordic_AddX_MUX_0_n_31) );
AND3_X1 g14810 ( .a(n_444), .b(n_698), .c(RESET), .o(n_706) );
NOR2_Z1 cordic_g471 ( .a(cordic_n_14), .b(Issue_Rst), .o(cordic_n_36) );
BUF_X2 newInst_1153 ( .a(newNet_1152), .o(newNet_1153) );
BUF_X2 newInst_326 ( .a(newNet_325), .o(newNet_326) );
NAND2_Z01 g15248 ( .a(n_315), .b(n_316), .o(n_412) );
NAND2_Z01 g15415 ( .a(CoreOutput_9_), .b(n_188), .o(n_235) );
NAND2_Z01 g13475 ( .a(n_721), .b(n_753), .o(n_809) );
NAND2_Z01 cordic_AddX_MUX_0_g284 ( .a(cordic_AddX_MUX_0_n_20), .b(cordic_AddX_MUX_0_n_3), .o(cordic_AddX_Atemp_13_) );
BUF_X2 newInst_713 ( .a(newNet_712), .o(newNet_713) );
AND2_X1 g38 ( .a(n_836), .b(n_856), .o(PO_AD_26) );
fflopd Config_Reg_reg_15_ ( .CK(newNet_1013), .D(n_633), .Q(Config_Reg_15_) );
INV_X1 g15523 ( .a(n_140), .o(n_141) );
BUF_X2 newInst_322 ( .a(newNet_102), .o(newNet_322) );
NAND2_Z01 cordic_AddX_MUX_1_g316 ( .a(cordic_BS1_6_), .b(cordic_AddX_MUX_1_n_0), .o(cordic_AddX_MUX_1_n_5) );
INV_X1 g13485 ( .a(n_799), .o(n_976) );
BUF_X2 newInst_528 ( .a(newNet_527), .o(newNet_528) );
BUF_X2 newInst_750 ( .a(newNet_440), .o(newNet_750) );
NAND2_Z01 g14992 ( .a(n_572), .b(Config_Reg_10_), .o(n_585) );
NAND2_Z01 cordic_Add0_MUX_0_g296 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_10_), .o(cordic_Add0_MUX_0_n_7) );
fflopd cordic_Angle_reg_6_ ( .CK(newNet_228), .D(cordic_n_105), .Q(cordic_Angle_6_) );
NAND2_Z01 g15252 ( .a(n_306), .b(n_307), .o(n_408) );
XOR2_X1 g13396 ( .a(n_883), .b(PO_AD_26), .o(n_884) );
NAND2_Z01 cordic_SH1_srl_35_26_g1221 ( .a(cordic_iteration_0_), .b(cordic_Y_14_), .o(cordic_SH1_srl_35_26_n_31) );
BUF_X2 newInst_1029 ( .a(newNet_217), .o(newNet_1029) );
BUF_X2 newInst_837 ( .a(newNet_836), .o(newNet_837) );
NAND2_Z01 g14987 ( .a(n_571), .b(CoreInput_6_), .o(n_590) );
BUF_X2 newInst_120 ( .a(newNet_119), .o(newNet_120) );
NAND2_Z01 g15617 ( .a(PI_FRAME_L), .b(PI_IRDY_L), .o(n_43) );
NOR2_Z1 cordic_Add0_MUX_0_g300 ( .a(cordic_Add0_MUX_0_n_1), .b(cordic_AngleCin), .o(cordic_Add0_Atemp_15_) );
BUF_X2 newInst_1027 ( .a(newNet_1026), .o(newNet_1027) );
XOR2_X1 g15489 ( .a(n_88), .b(n_79), .o(n_174) );
NOR2_Z1 g15420 ( .a(n_182), .b(n_122), .o(n_279) );
NOR3_Z1 g13504 ( .a(Idsel), .b(n_900), .c(PI_REQ64_L), .o(n_782) );
BUF_X2 newInst_554 ( .a(newNet_431), .o(newNet_554) );
XOR2_X1 cordic_Add0_Compl_g346 ( .a(cordic_Add0_Compl_n_33), .b(cordic_Add0_Compl_n_9), .o(cordic_SumAngle_10_) );
NAND2_Z01 g15005 ( .a(n_565), .b(n_557), .o(n_574) );
BUF_X2 newInst_711 ( .a(newNet_710), .o(newNet_711) );
fflopd cordic_Angle_reg_8_ ( .CK(newNet_214), .D(cordic_n_103), .Q(cordic_Angle_8_) );
XOR2_X1 cordic_AddX_g208 ( .a(cordic_AddX_Btemp_4_), .b(cordic_AddX_Y_2), .o(cordic_AddX_Btemp1_4_) );
BUF_X2 newInst_745 ( .a(newNet_744), .o(newNet_745) );
BUF_X2 newInst_1116 ( .a(newNet_1115), .o(newNet_1116) );
BUF_X2 newInst_872 ( .a(newNet_871), .o(newNet_872) );
NAND2_Z01 cordic_Add0_Add_g669 ( .a(cordic_Add0_Add_n_36), .b(cordic_Add0_Add_n_3), .o(cordic_Add0_Add_n_38) );
NAND2_Z01 cordic_SH1_srl_35_26_g1167 ( .a(cordic_SH1_srl_35_26_n_50), .b(cordic_iteration_1_), .o(cordic_SH1_srl_35_26_n_85) );
fflopd cordic_X_reg_1_ ( .CK(newNet_146), .D(cordic_n_54), .Q(cordic_X_1_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1160 ( .a(cordic_SH1_srl_35_26_n_82), .b(cordic_SH1_srl_35_26_n_63), .o(cordic_SH1_srl_35_26_n_92) );
NAND3_Z1 cordic_SH1_srl_35_26_g1118 ( .a(cordic_SH1_srl_35_26_n_105), .b(cordic_SH1_srl_35_26_n_107), .c(cordic_SH1_srl_35_26_n_104), .o(cordic_BS1_4_) );
BUF_X2 newInst_960 ( .a(newNet_959), .o(newNet_960) );
BUF_X2 newInst_935 ( .a(newNet_934), .o(newNet_935) );
NAND2_Z01 cordic_Add0_Add_g647 ( .a(cordic_Add0_Add_n_59), .b(cordic_Add0_Add_n_26), .o(cordic_Add0_Add_n_60) );
fflopd cordic_Angle_reg_1_ ( .CK(newNet_240), .D(cordic_n_110), .Q(cordic_Angle_1_) );
BUF_X2 newInst_988 ( .a(newNet_987), .o(newNet_988) );
BUF_X2 newInst_594 ( .a(newNet_593), .o(newNet_594) );
NAND2_Z01 cordic_Add0_MUX_0_g287 ( .a(cordic_Add0_MUX_0_n_2), .b(cordic_Angle_1_), .o(cordic_Add0_MUX_0_n_16) );
BUF_X2 newInst_816 ( .a(newNet_728), .o(newNet_816) );
BUF_X2 newInst_582 ( .a(newNet_581), .o(newNet_582) );
BUF_X2 newInst_38 ( .a(newNet_37), .o(newNet_38) );
NAND2_Z01 cordic_SH2_srl_35_26_g1239 ( .a(cordic_SH2_srl_35_26_n_0), .b(cordic_X_11_), .o(cordic_SH2_srl_35_26_n_10) );
NAND2_Z01 g15294 ( .a(n_275), .b(Access_Type_1_3_), .o(n_361) );
BUF_X2 newInst_971 ( .a(newNet_970), .o(newNet_971) );
NAND2_Z01 cordic_SH2_srl_35_26_g1188 ( .a(cordic_SH2_srl_35_26_n_44), .b(cordic_SH2_srl_35_26_n_3), .o(cordic_SH2_srl_35_26_n_64) );
NAND3_Z1 g15141 ( .a(n_332), .b(n_416), .c(n_10), .o(n_470) );
BUF_X2 newInst_264 ( .a(newNet_263), .o(newNet_264) );
BUF_X2 newInst_1036 ( .a(newNet_1035), .o(newNet_1036) );
NAND2_Z01 cordic_AddY_MUX_1_g314 ( .a(cordic_BS2_15_), .b(cordic_AddY_MUX_1_n_0), .o(cordic_AddY_MUX_1_n_7) );
NAND2_Z01 cordic_AddY_MUX_1_g279 ( .a(cordic_AddY_MUX_1_n_12), .b(cordic_AddY_MUX_1_n_25), .o(cordic_AddY_Btemp_0_) );
NOR2_Z1 g15559 ( .a(n_33), .b(Check_Data_Parity), .o(n_100) );
NOR2_Z1 g13438 ( .a(n_810), .b(n_710), .o(n_844) );
XOR2_X1 g15319 ( .a(n_163), .b(n_169), .o(n_341) );
NAND2_Z01 cordic_SH2_srl_35_26_g1197 ( .a(cordic_SH2_srl_35_26_n_8), .b(cordic_SH2_srl_35_26_n_35), .o(cordic_SH2_srl_35_26_n_55) );
BUF_X2 newInst_570 ( .a(newNet_569), .o(newNet_570) );
XOR2_X1 cordic_Add0_Add_g676 ( .a(cordic_Add0_n_12), .b(cordic_Add0_Atemp_11_), .o(cordic_Add0_Add_n_31) );
NAND2_Z01 cordic_SH1_srl_35_26_g1248 ( .a(cordic_SH1_srl_35_26_n_1), .b(cordic_SH1_srl_35_26_n_2), .o(cordic_SH1_srl_35_26_n_19) );
fflopd Trdy_Wait_Cnt_reg_3_ ( .CK(newNet_302), .D(n_417), .Q(Trdy_Wait_Cnt_3_) );
NAND2_Z01 g14931 ( .a(n_590), .b(n_520), .o(n_643) );
INV_X1 cordic_pla_g296 ( .a(cordic_pla_n_14), .o(cordic_pla_n_15) );
NAND2_Z01 cordic_SH1_srl_35_26_g1218 ( .a(cordic_iteration_0_), .b(cordic_Y_1_), .o(cordic_SH1_srl_35_26_n_34) );
BUF_X2 newInst_632 ( .a(newNet_631), .o(newNet_632) );
BUF_X2 newInst_769 ( .a(newNet_768), .o(newNet_769) );
NOR2_Z1 g15480 ( .a(n_131), .b(n_36), .o(n_179) );
NAND2_Z01 cordic_AddX_Add_g660 ( .a(cordic_AddX_Add_n_73), .b(cordic_AddX_Add_n_22), .o(cordic_AddX_Add_n_74) );
NAND2_Z01 g15343 ( .a(n_214), .b(CoreOutputReg_10_), .o(n_318) );
BUF_X2 newInst_309 ( .a(newNet_308), .o(newNet_309) );
BUF_X2 newInst_893 ( .a(newNet_72), .o(newNet_893) );
BUF_X2 newInst_572 ( .a(newNet_146), .o(newNet_572) );
BUF_X2 newInst_877 ( .a(newNet_876), .o(newNet_877) );
NAND2_Z01 cordic_SH2_srl_35_26_g1130 ( .a(cordic_SH2_srl_35_26_n_97), .b(cordic_SH2_srl_35_26_n_21), .o(cordic_SH2_srl_35_26_n_122) );
NAND2_Z01 cordic_AddX_MUX_1_g303 ( .a(cordic_AddX_Y_1), .b(cordic_X_4_), .o(cordic_AddX_MUX_1_n_18) );
BUF_X2 newInst_510 ( .a(newNet_509), .o(newNet_510) );
BUF_X2 newInst_228 ( .a(newNet_227), .o(newNet_228) );
BUF_X2 newInst_293 ( .a(newNet_292), .o(newNet_293) );
NAND2_Z01 cordic_SH1_srl_35_26_g1143 ( .a(cordic_SH1_srl_35_26_n_92), .b(cordic_SH1_srl_35_26_n_18), .o(cordic_SH1_srl_35_26_n_109) );
NAND2_Z01 g15268 ( .a(n_258), .b(n_259), .o(n_392) );
NAND2_Z01 g13492 ( .a(n_737), .b(n_757), .o(n_792) );
NOR2_Z1 cordic_g454 ( .a(cordic_n_24), .b(Issue_Rst), .o(cordic_n_53) );
NAND2_Z01 g15075 ( .a(n_494), .b(PI_AD_0), .o(n_533) );
BUF_X2 newInst_612 ( .a(newNet_611), .o(newNet_612) );
BUF_X2 newInst_973 ( .a(newNet_269), .o(newNet_973) );
BUF_X2 newInst_538 ( .a(newNet_537), .o(newNet_538) );
fflopd Config_Reg_reg_3_ ( .CK(newNet_892), .D(n_664), .Q(Config_Reg_3_) );
fflopd Core_Cnt_reg_2_ ( .CK(newNet_534), .D(n_181), .Q(Core_Cnt_2_) );
BUF_X2 newInst_166 ( .a(newNet_165), .o(newNet_166) );
BUF_X2 newInst_733 ( .a(newNet_732), .o(newNet_733) );
BUF_X2 newInst_47 ( .a(newNet_46), .o(newNet_47) );
NAND2_Z01 g15236 ( .a(n_274), .b(Access_Address_1_23_), .o(n_424) );
BUF_X2 newInst_391 ( .a(newNet_390), .o(newNet_391) );
NOR2_Z1 cordic_g469 ( .a(cordic_n_4), .b(Issue_Rst), .o(cordic_n_38) );
BUF_X2 newInst_191 ( .a(newNet_190), .o(newNet_191) );
NOR2_Z1 g15512 ( .a(n_116), .b(n_16), .o(n_149) );
BUF_X2 newInst_253 ( .a(newNet_147), .o(newNet_253) );
NAND2_Z01 cordic_AddY_MUX_0_g313 ( .a(cordic_AddY_MUX_0_n_0), .b(cordic_Y_7_), .o(cordic_AddY_MUX_0_n_8) );
XOR2_X1 cordic_Add0_Add_g684 ( .a(cordic_Add0_n_4), .b(cordic_Add0_Atemp_3_), .o(cordic_Add0_Add_n_23) );
BUF_X2 newInst_486 ( .a(newNet_485), .o(newNet_486) );
NAND2_Z01 g15429 ( .a(n_212), .b(n_125), .o(n_275) );
BUF_X2 newInst_925 ( .a(newNet_924), .o(newNet_925) );
fflopd Access_Address_1_reg_27_ ( .CK(newNet_1141), .D(n_476), .Q(Access_Address_1_27_) );
BUF_X2 newInst_759 ( .a(newNet_758), .o(newNet_759) );
NAND2_Z01 cordic_Add0_MUX_1_g290 ( .a(cordic_tanangle_11_), .b(cordic_Add0_MUX_1_n_2), .o(cordic_Add0_MUX_1_n_11) );
INV_X1 g15444 ( .a(n_209), .o(n_210) );
NAND2_Z01 g15458 ( .a(n_138), .b(PI_CBE_L_3), .o(n_200) );
NAND2_Z01 cordic_Add0_Add_g644 ( .a(cordic_Add0_Add_n_62), .b(cordic_Add0_Add_n_31), .o(cordic_Add0_Add_n_63) );
NAND2_Z01 cordic_AddX_MUX_0_g280 ( .a(cordic_AddX_MUX_0_n_23), .b(cordic_AddX_MUX_0_n_6), .o(cordic_AddX_Atemp_11_) );
AND2_X1 g333 ( .a(TAR_TRI_A), .b(n_856), .o(PO_AD_61) );
BUF_X2 newInst_566 ( .a(newNet_565), .o(newNet_566) );
BUF_X2 newInst_577 ( .a(newNet_576), .o(newNet_577) );
NAND2_Z01 cordic_g438 ( .a(cordic_SumAngle_15_), .b(cordic_n_7), .o(cordic_n_69) );
NAND2_Z01 g14962 ( .a(n_572), .b(Config_Reg_28_), .o(n_615) );
BUF_X2 newInst_230 ( .a(newNet_229), .o(newNet_230) );
NAND2_Z01 g15392 ( .a(CoreOutput_29_), .b(n_188), .o(n_258) );
NAND3_Z1 g15561 ( .a(Core_Cnt_1_), .b(Core_Cnt_2_), .c(Core_Cnt_3_), .o(n_99) );
NAND2_Z01 cordic_Add0_MUX_0_g260 ( .a(cordic_Add0_MUX_0_n_30), .b(cordic_Add0_MUX_0_n_16), .o(cordic_Add0_Atemp_1_) );
NAND2_Z01 cordic_SH1_srl_35_26_g1158 ( .a(cordic_SH1_srl_35_26_n_81), .b(cordic_SH1_srl_35_26_n_64), .o(cordic_SH1_srl_35_26_n_95) );

endmodule
