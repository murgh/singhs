module cordic_ispd ;

// Start PIs
input beta_11;
input beta_24;
input beta_8;
input beta_5;
input beta_25;
input beta_22;
input beta_30;
input beta_6;
input beta_27;
input beta_3;
input beta_13;
input beta_29;
input beta_12;
input beta_15;
input tau_clk;
input beta_20;
input beta_21;
input beta_28;
input beta_1;
input beta_2;
input beta_9;
input beta_7;
input rst;
input beta_16;
input beta_18;
input beta_0;
input beta_19;
input beta_14;
input beta_10;
input beta_31;
input beta_17;
input beta_23;
input beta_4;
input beta_26;

// Start POs
output cos_out_2;
output cos_out_13;
output sin_out_2;
output sin_out_17;
output sin_out_21;
output sin_out_8;
output sin_out_19;
output cos_out_30;
output cos_out_28;
output sin_out_20;
output cos_out_10;
output cos_out_17;
output cos_out_18;
output sin_out_16;
output cos_out_7;
output cos_out_11;
output sin_out_29;
output sin_out_9;
output sin_out_3;
output cos_out_4;
output sin_out_27;
output cos_out_12;
output cos_out_15;
output cos_out_19;
output sin_out_22;
output sin_out_7;
output cos_out_23;
output sin_out_31;
output sin_out_14;
output cos_out_26;
output cos_out_14;
output sin_out_23;
output sin_out_5;
output cos_out_25;
output sin_out_1;
output cos_out_1;
output cos_out_9;
output sin_out_24;
output cos_out_20;
output sin_out_30;
output sin_out_26;
output cos_out_0;
output sin_out_15;
output sin_out_28;
output sin_out_10;
output sin_out_13;
output cos_out_31;
output sin_out_0;
output cos_out_29;
output cos_out_3;
output cos_out_21;
output cos_out_6;
output cos_out_16;
output sin_out_11;
output cos_out_24;
output sin_out_4;
output sin_out_25;
output sin_out_18;
output sin_out_12;
output cos_out_27;
output cos_out_5;
output cos_out_8;
output cos_out_22;
output sin_out_6;

// Start wires
wire n_8095;
wire n_43417;
wire n_29500;
wire FE_RN_1356_0;
wire FE_RN_304_0;
wire n_6891;
wire n_25465;
wire n_4132;
wire n_6068;
wire n_9472;
wire n_40843;
wire n_685;
wire n_2907;
wire n_6543;
wire n_9953;
wire n_37946;
wire n_38956;
wire n_17324;
wire n_1266;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_24_;
wire n_33903;
wire FE_RN_539_0;
wire newNet_3271;
wire n_23457;
wire n_25827;
wire n_41200;
wire n_41443;
wire n_26528;
wire n_98;
wire n_37097;
wire FE_OCP_RBN1184_n_14638;
wire n_20476;
wire n_5731;
wire n_30165;
wire n_43681;
wire n_2794;
wire n_39657;
wire n_19568;
wire n_32806;
wire FE_RN_1438_0;
wire n_3935;
wire n_36591;
wire n_28388;
wire n_43023;
wire n_15533;
wire n_17259;
wire FE_OCPUNCON3145_n_21058;
wire newNet_562;
wire n_36923;
wire n_14094;
wire n_12555;
wire n_14554;
wire n_18925;
wire n_14012;
wire n_9864;
wire n_26910;
wire n_13478;
wire n_23017;
wire n_24923;
wire n_7231;
wire n_16645;
wire n_25006;
wire n_43803;
wire n_9162;
wire n_6175;
wire n_44814;
wire n_38770;
wire n_38484;
wire n_35972;
wire delay_xor_ln22_unr3_stage2_stallmux_q_12_;
wire n_3167;
wire n_24893;
wire n_24140;
wire FE_OFN812_n_2405;
wire n_7945;
wire n_23074;
wire n_8079;
wire n_36120;
wire n_35714;
wire n_35738;
wire n_9916;
wire FE_OCP_RBN2485_n_38601;
wire n_36236;
wire n_4042;
wire n_10014;
wire n_2158;
wire n_18406;
wire newNet_1202;
wire n_18590;
wire n_6945;
wire n_17214;
wire n_27463;
wire n_10992;
wire n_43000;
wire n_20268;
wire n_37211;
wire FE_OCP_RBN2484_n_38601;
wire newNet_1237;
wire n_20024;
wire n_28536;
wire n_11017;
wire n_6587;
wire n_25607;
wire FE_OCP_RBN2996_n_11004;
wire n_27565;
wire n_31477;
wire n_15518;
wire n_3845;
wire n_7122;
wire n_37780;
wire n_39559;
wire n_2148;
wire n_34222;
wire FE_OCP_RBN3424_n_37794;
wire n_29172;
wire n_35483;
wire n_32551;
wire n_35427;
wire n_39958;
wire n_1233;
wire n_27777;
wire n_12510;
wire n_17680;
wire newNet_1446;
wire n_6737;
wire n_11898;
wire n_26549;
wire FE_OCP_RBN2928_n_39614;
wire FE_OCPN1741_n_19138;
wire n_38636;
wire n_3472;
wire n_10785;
wire newNet_1895;
wire n_24874;
wire n_11569;
wire n_30427;
wire n_5684;
wire n_26506;
wire FE_OCP_RBN3294_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire n_27670;
wire FE_RN_1374_0;
wire n_21921;
wire n_9386;
wire n_12875;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_27_;
wire n_39907;
wire n_31424;
wire n_25185;
wire n_35095;
wire n_11885;
wire n_39424;
wire n_15398;
wire n_33081;
wire n_36919;
wire n_38281;
wire n_4110;
wire n_15878;
wire n_13900;
wire n_36406;
wire n_40765;
wire n_15595;
wire delay_add_ln22_unr20_stage8_stallmux_q_21_;
wire n_11622;
wire newNet_721;
wire n_43317;
wire n_41313;
wire FE_RN_1519_0;
wire n_22728;
wire newNet_967;
wire n_28034;
wire newNet_1704;
wire n_23509;
wire n_42290;
wire newNet_867;
wire n_1500;
wire n_5845;
wire n_14568;
wire newNet_882;
wire n_3467;
wire n_21885;
wire n_13173;
wire n_41438;
wire n_20316;
wire n_27168;
wire n_38131;
wire n_3500;
wire FE_OCP_RBN1129_n_24179;
wire n_34632;
wire n_10996;
wire n_43334;
wire n_44881;
wire n_4386;
wire n_24568;
wire n_13851;
wire n_13211;
wire n_7250;
wire n_10536;
wire n_6206;
wire FE_OCP_RBN3646_n_44490;
wire n_2065;
wire n_12861;
wire n_6098;
wire n_19231;
wire n_24632;
wire n_37661;
wire n_6618;
wire n_1988;
wire FE_RN_1440_0;
wire n_9701;
wire n_34526;
wire delay_xor_ln22_unr12_stage5_stallmux_q_18_;
wire n_3950;
wire newNet_3132;
wire n_6825;
wire FE_RN_1714_0;
wire newNet_2433;
wire n_14805;
wire n_477;
wire n_13620;
wire n_8721;
wire n_29332;
wire n_24067;
wire n_23053;
wire n_6507;
wire n_5868;
wire FE_RN_1752_0;
wire n_3236;
wire n_10038;
wire n_8048;
wire newNet_1175;
wire newNet_1949;
wire n_27504;
wire n_19507;
wire n_38350;
wire n_12049;
wire n_13084;
wire n_11433;
wire n_46182;
wire newNet_3396;
wire n_41254;
wire n_39785;
wire n_28803;
wire cos_out_19;
wire n_17636;
wire n_26223;
wire n_16106;
wire n_20693;
wire n_5656;
wire n_27546;
wire n_18900;
wire n_2833;
wire n_17371;
wire n_26821;
wire n_27355;
wire n_6984;
wire n_31075;
wire newNet_748;
wire n_19654;
wire n_30958;
wire n_35391;
wire n_5378;
wire n_24313;
wire n_2415;
wire n_38725;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_24_;
wire n_11173;
wire newNet_1315;
wire n_42592;
wire n_24457;
wire newNet_35;
wire n_6708;
wire n_4561;
wire n_30582;
wire n_12478;
wire newNet_2271;
wire n_33053;
wire n_27744;
wire n_8690;
wire n_41890;
wire n_17357;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_27_;
wire n_8966;
wire n_38240;
wire n_29246;
wire n_5067;
wire n_21537;
wire n_32024;
wire n_22660;
wire n_23618;
wire n_30690;
wire n_6634;
wire n_2023;
wire n_20064;
wire FE_RN_577_0;
wire n_2615;
wire n_5823;
wire n_24036;
wire n_3885;
wire n_38440;
wire n_19210;
wire n_3391;
wire n_10208;
wire FE_OCP_RBN2390_n_19434;
wire n_36504;
wire FE_OCP_RBN2511_n_19884;
wire n_31409;
wire n_3086;
wire n_21377;
wire n_499;
wire n_19055;
wire n_46975;
wire n_245;
wire n_20116;
wire n_29063;
wire n_14695;
wire n_39104;
wire n_40942;
wire newNet_2330;
wire n_40842;
wire n_21358;
wire FE_RN_988_0;
wire n_2851;
wire n_11662;
wire n_41499;
wire n_28276;
wire n_7400;
wire n_6742;
wire n_15983;
wire n_40292;
wire FE_RN_961_0;
wire n_967;
wire n_31171;
wire n_26594;
wire n_13052;
wire n_7865;
wire n_44101;
wire n_833;
wire newNet_87;
wire n_666;
wire n_19926;
wire n_16249;
wire n_22684;
wire n_36619;
wire n_28378;
wire n_12964;
wire n_15813;
wire n_12682;
wire n_30066;
wire n_13507;
wire newNet_259;
wire newNet_2643;
wire n_33702;
wire n_14215;
wire n_131;
wire n_37674;
wire n_33924;
wire n_7475;
wire n_31721;
wire n_24320;
wire n_15022;
wire newNet_2310;
wire n_18728;
wire n_38266;
wire n_1074;
wire n_30103;
wire newNet_526;
wire n_20168;
wire n_7501;
wire n_31971;
wire newNet_2147;
wire n_31699;
wire FE_RN_1692_0;
wire FE_RN_1117_0;
wire n_23012;
wire FE_OCP_RBN2345_FE_OCPN870_n_2737;
wire FE_OCP_RBN1174_n_18981;
wire newNet_281;
wire n_46245;
wire n_16665;
wire n_35482;
wire n_36800;
wire n_16996;
wire n_41383;
wire FE_OCP_RBN2052_delay_xor_ln22_unr15_stage6_stallmux_q_2_;
wire n_9855;
wire n_754;
wire n_2378;
wire newNet_2958;
wire n_25020;
wire n_14607;
wire n_40011;
wire n_33624;
wire n_30461;
wire n_31834;
wire n_43826;
wire n_14613;
wire n_5409;
wire n_15915;
wire n_31008;
wire n_12005;
wire newNet_766;
wire n_3457;
wire n_39829;
wire n_34743;
wire n_5710;
wire FE_OCP_RBN2407_n_8242;
wire n_28581;
wire n_9399;
wire newNet_1610;
wire n_32999;
wire n_29813;
wire n_23562;
wire n_35866;
wire n_14846;
wire FE_OCP_RBN3466_n_7886;
wire n_27656;
wire FE_OCPN1030_n_28423;
wire n_29051;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_12_;
wire n_30199;
wire n_27434;
wire n_21824;
wire n_23400;
wire n_38538;
wire n_40658;
wire n_5892;
wire n_40615;
wire n_18664;
wire n_35958;
wire newNet_2267;
wire n_7871;
wire n_25224;
wire n_19030;
wire n_16836;
wire n_41041;
wire n_9041;
wire n_26365;
wire n_36023;
wire n_6356;
wire newNet_476;
wire n_37948;
wire n_15308;
wire n_11122;
wire n_22457;
wire n_40439;
wire n_17505;
wire n_33327;
wire n_34003;
wire FE_RN_479_0;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_10_;
wire n_7839;
wire newNet_2399;
wire n_4231;
wire n_29252;
wire n_23635;
wire n_26479;
wire FE_OCPN1861_n_30319;
wire n_9670;
wire n_20830;
wire n_36495;
wire n_24384;
wire n_34786;
wire n_47263;
wire n_3727;
wire newNet_1323;
wire FE_OCP_RBN2466_n_8393;
wire n_1805;
wire n_29576;
wire n_9641;
wire n_28010;
wire newNet_15;
wire n_26744;
wire n_1184;
wire n_18175;
wire n_22129;
wire n_25572;
wire newNet_2061;
wire n_9647;
wire n_17594;
wire newNet_2630;
wire n_28071;
wire n_40305;
wire n_30551;
wire n_43068;
wire n_40387;
wire FE_OCP_RBN1156_n_18375;
wire n_9291;
wire n_41926;
wire n_13206;
wire n_4061;
wire n_5259;
wire newNet_1835;
wire n_5807;
wire n_10640;
wire n_25746;
wire FE_OCP_RBN3619_n_15135;
wire n_19147;
wire n_20615;
wire n_1567;
wire n_3860;
wire n_40247;
wire n_8127;
wire n_25807;
wire n_37287;
wire n_37929;
wire n_14116;
wire n_15276;
wire n_17687;
wire n_41561;
wire n_40479;
wire n_27493;
wire FE_RN_1305_0;
wire n_30259;
wire n_43009;
wire n_28707;
wire n_33220;
wire n_24822;
wire n_2987;
wire n_33735;
wire n_4498;
wire n_27270;
wire n_43700;
wire n_13495;
wire n_6597;
wire n_20514;
wire n_23687;
wire n_36369;
wire n_47246;
wire FE_RN_1803_0;
wire n_23117;
wire FE_RN_932_0;
wire n_39173;
wire FE_OCPN3172_n_34222;
wire n_27037;
wire n_10047;
wire FE_RN_1023_0;
wire n_4217;
wire n_10739;
wire n_1917;
wire n_36846;
wire newNet_1090;
wire n_11243;
wire n_42731;
wire n_23411;
wire newNet_217;
wire newNet_696;
wire n_1114;
wire newNet_2686;
wire n_28715;
wire n_27046;
wire n_23588;
wire n_19105;
wire n_19722;
wire n_29892;
wire n_21904;
wire n_15674;
wire n_41958;
wire n_26521;
wire n_23741;
wire n_20505;
wire n_5785;
wire n_5984;
wire n_34591;
wire n_41795;
wire n_1161;
wire n_37236;
wire n_44621;
wire n_34343;
wire FE_OCP_RBN2898_n_45484;
wire n_33952;
wire n_26853;
wire n_38653;
wire n_39843;
wire newNet_1552;
wire n_47185;
wire n_25998;
wire FE_RN_190_0;
wire n_12592;
wire newNet_1101;
wire n_23862;
wire n_25507;
wire n_35401;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_21_;
wire n_44053;
wire n_432;
wire n_25141;
wire n_35921;
wire n_44042;
wire FE_OCPN1014_n_32820;
wire n_36473;
wire n_23336;
wire n_6053;
wire n_876;
wire n_16534;
wire n_21864;
wire n_43624;
wire FE_OCP_RBN1217_n_20595;
wire n_32035;
wire n_40921;
wire newNet_2842;
wire n_337;
wire newNet_2392;
wire n_30963;
wire newNet_2200;
wire n_22591;
wire n_7413;
wire n_29597;
wire n_38417;
wire n_7530;
wire n_38765;
wire FE_OCP_RBN1142_n_25816;
wire n_24995;
wire n_14963;
wire n_22488;
wire n_36162;
wire sin_out_26;
wire FE_RN_1166_0;
wire n_18576;
wire n_22783;
wire n_41049;
wire delay_add_ln22_unr27_stage10_stallmux_q_10_;
wire n_28342;
wire n_14062;
wire n_7695;
wire n_11214;
wire n_26401;
wire n_13879;
wire n_4190;
wire n_24238;
wire n_12056;
wire n_37478;
wire n_3109;
wire n_16736;
wire n_41851;
wire n_42645;
wire n_31400;
wire n_8517;
wire n_33110;
wire n_7928;
wire n_6212;
wire delay_add_ln22_unr23_stage9_stallmux_q_4_;
wire n_43568;
wire n_36844;
wire n_37872;
wire n_23136;
wire n_28189;
wire n_18321;
wire n_8529;
wire n_28002;
wire n_5598;
wire n_13371;
wire n_46236;
wire n_22743;
wire n_18987;
wire sin_out_14;
wire n_43634;
wire FE_OCP_RBN3502_n_38592;
wire newNet_1283;
wire newNet_2893;
wire n_442;
wire n_9267;
wire n_17532;
wire n_13704;
wire n_20495;
wire n_39205;
wire newNet_3740;
wire n_22604;
wire n_9521;
wire n_26277;
wire n_34971;
wire n_35616;
wire n_22540;
wire newNet_608;
wire n_27627;
wire n_36275;
wire n_41645;
wire n_36957;
wire n_34417;
wire FE_RN_1645_0;
wire newNet_3437;
wire n_12703;
wire n_1416;
wire n_3812;
wire n_29687;
wire n_24607;
wire n_520;
wire n_15702;
wire n_17817;
wire n_40340;
wire newNet_2110;
wire n_14593;
wire FE_RN_1630_0;
wire n_23367;
wire n_38446;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_20_;
wire newNet_1863;
wire n_30334;
wire newNet_2378;
wire n_2546;
wire FE_RN_1183_0;
wire FE_OCP_RBN2441_n_8402;
wire n_31323;
wire n_41628;
wire n_5486;
wire n_41422;
wire n_32923;
wire n_40298;
wire n_21955;
wire n_28261;
wire FE_OCP_RBN2151_n_22822;
wire n_17464;
wire FE_OCP_RBN1836_FE_RN_1542_0;
wire n_41026;
wire n_157;
wire n_31266;
wire n_6107;
wire n_41065;
wire n_22854;
wire n_13109;
wire n_2753;
wire n_23523;
wire n_20640;
wire n_25118;
wire n_19748;
wire n_36238;
wire n_26727;
wire n_43276;
wire FE_RN_1292_0;
wire n_20193;
wire n_724;
wire n_2592;
wire n_40282;
wire FE_OCP_RBN3414_n_12739;
wire n_5535;
wire n_37816;
wire n_5407;
wire n_11089;
wire n_31880;
wire FE_OCP_RBN1358_FE_RN_677_0;
wire newNet_1799;
wire n_30457;
wire n_8170;
wire n_10325;
wire n_41981;
wire n_20822;
wire n_4978;
wire n_30573;
wire n_33423;
wire n_11376;
wire n_21455;
wire n_1012;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_14_;
wire FE_RN_1225_0;
wire n_34915;
wire n_38059;
wire n_12450;
wire n_13378;
wire newNet_3188;
wire n_5463;
wire n_38741;
wire n_7085;
wire n_9114;
wire n_29505;
wire n_9712;
wire newNet_3541;
wire n_13662;
wire n_43911;
wire FE_OCP_RBN2138_n_11909;
wire FE_OCP_RBN2121_n_45224;
wire n_29359;
wire newNet_1426;
wire n_28467;
wire FE_RN_905_0;
wire n_43321;
wire n_41697;
wire n_4084;
wire n_34713;
wire n_43154;
wire newNet_343;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_13_;
wire n_18376;
wire n_14977;
wire n_15456;
wire n_30232;
wire delay_add_ln22_unr27_stage10_stallmux_q_14_;
wire FE_RN_607_0;
wire newNet_2996;
wire n_37126;
wire n_24426;
wire n_37838;
wire n_12545;
wire n_17900;
wire n_12223;
wire n_70;
wire n_12354;
wire delay_xor_ln21_unr6_stage3_stallmux_q_16_;
wire delay_add_ln22_unr23_stage9_stallmux_q_6_;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_22_;
wire n_20606;
wire n_21556;
wire newNet_2997;
wire newNet_2834;
wire n_23904;
wire n_40020;
wire n_43717;
wire FE_OCP_RBN3016_n_31117;
wire n_25039;
wire n_37283;
wire n_33553;
wire FE_RN_796_0;
wire newNet_2218;
wire n_16018;
wire delay_add_ln22_unr14_stage6_stallmux_q_30_;
wire FE_RN_1580_0;
wire n_11422;
wire n_15719;
wire n_17602;
wire delay_xor_ln22_unr3_stage2_stallmux_q_5_;
wire n_30597;
wire n_41710;
wire FE_OCP_RBN3067_n_43230;
wire n_23521;
wire beta_8;
wire n_8746;
wire n_19993;
wire n_5925;
wire n_36736;
wire FE_OCP_RBN3615_n_20249;
wire n_17778;
wire n_37071;
wire n_22688;
wire FE_OCP_RBN2620_n_44561;
wire n_19755;
wire n_14201;
wire n_28636;
wire n_35121;
wire n_41577;
wire n_18951;
wire n_32424;
wire newNet_169;
wire n_41533;
wire n_47334;
wire n_21542;
wire FE_OCPN1501_n_20723;
wire n_3453;
wire n_41630;
wire newNet_1953;
wire n_14293;
wire n_10161;
wire n_1100;
wire n_7975;
wire n_32777;
wire FE_OCP_RBN3659_n_15314;
wire n_43555;
wire n_25148;
wire n_35057;
wire n_33122;
wire n_34553;
wire n_3151;
wire n_8469;
wire n_24407;
wire FE_OCP_RBN3514_n_13960;
wire n_17438;
wire FE_RN_544_0;
wire n_36822;
wire newNet_3344;
wire n_12773;
wire n_43168;
wire FE_OCP_RBN2709_n_15135;
wire n_37346;
wire n_16463;
wire n_46996;
wire n_27183;
wire delay_xor_ln22_unr3_stage2_stallmux_q_24_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_27_;
wire n_30242;
wire FE_RN_1020_0;
wire n_13998;
wire n_29231;
wire n_8061;
wire n_25531;
wire n_21228;
wire n_13559;
wire n_4166;
wire n_7317;
wire n_12051;
wire FE_OCP_RBN3449_n_37945;
wire n_34411;
wire n_39355;
wire n_29111;
wire n_34083;
wire n_25463;
wire n_38941;
wire n_21058;
wire n_39938;
wire n_41114;
wire FE_RN_602_0;
wire n_12951;
wire n_42812;
wire n_27104;
wire FE_OCP_RBN3836_n_19241;
wire n_32522;
wire n_22833;
wire n_40220;
wire n_29217;
wire n_36174;
wire n_26864;
wire n_607;
wire n_2307;
wire n_14354;
wire n_1147;
wire n_21775;
wire n_27838;
wire n_1527;
wire n_40934;
wire FE_OCP_RBN2882_n_26318;
wire n_16570;
wire n_13294;
wire newNet_1675;
wire n_29784;
wire n_41407;
wire FE_OCPN1048_n_24819;
wire n_40747;
wire n_712;
wire n_6010;
wire n_9601;
wire n_16307;
wire n_43183;
wire n_30053;
wire n_25433;
wire n_6380;
wire n_5005;
wire n_7774;
wire n_34190;
wire n_11863;
wire n_39373;
wire newNet_3515;
wire n_6915;
wire n_19334;
wire n_36641;
wire n_31185;
wire n_21609;
wire newNet_2194;
wire newNet_1041;
wire newNet_3632;
wire n_17132;
wire n_37889;
wire newNet_1266;
wire n_22239;
wire n_16481;
wire n_3211;
wire n_24076;
wire n_23703;
wire newNet_704;
wire n_31991;
wire n_19520;
wire newNet_668;
wire n_7351;
wire n_34163;
wire n_34208;
wire n_39152;
wire n_21560;
wire newNet_949;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_11_;
wire n_921;
wire n_43129;
wire n_25189;
wire n_11917;
wire n_17025;
wire FE_OCP_RBN3107_n_22590;
wire newNet_3447;
wire n_18176;
wire n_39898;
wire FE_OCP_RBN2988_n_35539;
wire n_22710;
wire n_22279;
wire delay_xor_ln22_unr18_stage7_stallmux_q_1_;
wire FE_OCP_RBN2707_n_15135;
wire FE_OCP_RBN2518_n_8762;
wire n_36390;
wire newNet_1608;
wire n_2848;
wire n_15549;
wire n_24059;
wire n_1783;
wire n_28132;
wire n_13159;
wire n_27113;
wire n_8435;
wire n_18227;
wire n_32232;
wire n_3012;
wire n_18193;
wire n_39929;
wire n_42120;
wire n_8315;
wire n_33029;
wire n_19128;
wire n_34764;
wire n_28307;
wire n_31537;
wire n_1789;
wire n_7730;
wire n_27613;
wire FE_OCPN1447_n_27463;
wire n_657;
wire n_4211;
wire n_11494;
wire n_849;
wire n_14839;
wire n_34754;
wire n_12584;
wire n_34056;
wire n_12832;
wire n_8271;
wire newNet_1481;
wire n_47003;
wire n_35262;
wire n_30539;
wire n_38856;
wire n_7518;
wire newNet_3037;
wire n_598;
wire FE_OCP_RBN2989_n_35539;
wire FE_RN_524_0;
wire FE_OCP_RBN2525_n_24902;
wire n_39742;
wire n_24492;
wire n_22479;
wire n_26304;
wire n_533;
wire n_26253;
wire FE_OCP_RBN2766_n_4376;
wire n_30273;
wire n_19487;
wire n_1099;
wire n_32946;
wire n_15754;
wire n_39962;
wire n_16902;
wire FE_OFN820_n_4333;
wire newNet_1566;
wire n_14307;
wire n_15032;
wire n_27597;
wire n_26491;
wire n_38716;
wire n_985;
wire n_1848;
wire n_16884;
wire FE_OCPN1416_FE_OCP_RBN1362_n_20504;
wire n_41340;
wire n_21107;
wire n_21408;
wire n_16852;
wire n_24162;
wire n_29036;
wire n_31205;
wire n_42084;
wire n_34645;
wire n_15160;
wire newNet_264;
wire n_4824;
wire n_11413;
wire n_9236;
wire n_17115;
wire n_27529;
wire n_39683;
wire n_27302;
wire n_29731;
wire delay_add_ln22_unr11_stage5_stallmux_q_24_;
wire FE_RN_1868_0;
wire n_23786;
wire n_25218;
wire FE_OCP_RBN2051_delay_xor_ln22_unr15_stage6_stallmux_q_2_;
wire n_15998;
wire n_12634;
wire n_12789;
wire n_38622;
wire n_7154;
wire newNet_2625;
wire n_28850;
wire n_41174;
wire n_36709;
wire n_42406;
wire n_10607;
wire n_7697;
wire n_14165;
wire n_10796;
wire n_5900;
wire newNet_2816;
wire newNet_2793;
wire n_14768;
wire n_42942;
wire newNet_2454;
wire n_37490;
wire n_3983;
wire newNet_1666;
wire FE_OCPN1466_n_13014;
wire n_37098;
wire n_41163;
wire n_42425;
wire n_26215;
wire n_34260;
wire n_40853;
wire n_42391;
wire n_11032;
wire n_21036;
wire n_26124;
wire n_40312;
wire n_29677;
wire n_771;
wire n_41213;
wire FE_RN_1564_0;
wire n_22652;
wire n_37862;
wire n_5962;
wire newNet_2546;
wire n_8189;
wire n_29130;
wire newNet_999;
wire n_15281;
wire newNet_751;
wire n_30475;
wire delay_add_ln22_unr20_stage8_stallmux_q_7_;
wire n_6083;
wire n_32116;
wire n_23917;
wire n_13320;
wire n_10217;
wire n_25294;
wire n_9185;
wire n_7547;
wire n_39297;
wire n_20674;
wire n_26005;
wire newNet_144;
wire n_4324;
wire n_8179;
wire n_10846;
wire n_5502;
wire n_15082;
wire FE_OCP_RBN3494_n_19390;
wire n_13618;
wire n_32244;
wire n_1967;
wire n_8647;
wire n_21781;
wire n_37146;
wire n_26662;
wire n_21710;
wire n_29961;
wire n_21487;
wire n_19941;
wire FE_RN_997_0;
wire FE_RN_1006_0;
wire n_3120;
wire n_28041;
wire n_40791;
wire newNet_3659;
wire n_35115;
wire n_19604;
wire n_31882;
wire n_16847;
wire newNet_953;
wire n_19060;
wire newNet_586;
wire n_8847;
wire n_14318;
wire newNet_898;
wire n_31011;
wire n_40402;
wire n_7957;
wire n_12072;
wire n_13443;
wire n_20965;
wire n_14189;
wire n_27799;
wire n_12659;
wire n_10186;
wire n_29958;
wire n_41510;
wire n_108;
wire n_36581;
wire n_31634;
wire n_37756;
wire n_21656;
wire n_27019;
wire n_34034;
wire n_43450;
wire n_22645;
wire n_39015;
wire n_41772;
wire n_36447;
wire newNet_1774;
wire n_23513;
wire n_1884;
wire n_25616;
wire n_28352;
wire n_14247;
wire n_42044;
wire n_29910;
wire n_24914;
wire n_9407;
wire n_13073;
wire n_24751;
wire n_39277;
wire n_42297;
wire n_11770;
wire n_43357;
wire n_20911;
wire n_25077;
wire n_18652;
wire n_43775;
wire n_4763;
wire FE_OCP_RBN1187_n_14823;
wire n_10320;
wire n_36862;
wire n_38513;
wire n_14457;
wire FE_OCP_DRV_N3160_n_31303;
wire n_6853;
wire n_7857;
wire FE_OCPN3768_FE_OCP_RBN2375_n_8221;
wire n_16112;
wire n_25919;
wire n_20325;
wire FE_OFN78_n_4117;
wire n_15992;
wire n_8221;
wire n_20443;
wire n_8887;
wire n_42631;
wire n_41378;
wire FE_OCP_RBN2759_n_9843;
wire n_32435;
wire n_8953;
wire n_11333;
wire n_16182;
wire n_16108;
wire n_37030;
wire FE_RN_442_0;
wire n_35500;
wire n_265;
wire n_21139;
wire n_35183;
wire n_2877;
wire n_2003;
wire n_29467;
wire n_36188;
wire n_42279;
wire n_34354;
wire n_10551;
wire n_9851;
wire n_10638;
wire n_30084;
wire n_40675;
wire FE_RN_1164_0;
wire n_23426;
wire n_21730;
wire newNet_1062;
wire n_2165;
wire n_26577;
wire n_635;
wire n_928;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_6_;
wire FE_OCP_DRV_N3150_n_12773;
wire n_10595;
wire n_16703;
wire n_17503;
wire n_24015;
wire n_15655;
wire n_16175;
wire n_22362;
wire n_19021;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_7_;
wire n_33517;
wire n_45202;
wire n_2496;
wire n_44735;
wire n_24955;
wire delay_add_ln22_unr17_stage7_stallmux_q_30_;
wire n_34933;
wire n_7041;
wire FE_OCP_RBN2974_n_5531;
wire n_34178;
wire n_34323;
wire n_39593;
wire n_42784;
wire newNet_647;
wire n_10914;
wire FE_RN_193_0;
wire n_11769;
wire n_19384;
wire delay_xor_ln21_unr6_stage3_stallmux_q_25_;
wire n_8381;
wire n_9932;
wire n_21132;
wire newNet_2086;
wire newNet_1739;
wire n_21723;
wire n_11369;
wire n_30792;
wire n_30158;
wire n_28055;
wire n_40627;
wire n_41012;
wire FE_OCP_RBN3028_n_39942;
wire n_27216;
wire n_7600;
wire n_28878;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_16_;
wire n_38121;
wire n_41887;
wire n_46156;
wire n_33676;
wire n_28688;
wire n_39385;
wire n_41587;
wire n_23350;
wire n_35965;
wire n_6782;
wire n_7024;
wire newNet_3567;
wire n_34823;
wire n_27908;
wire FE_RN_1517_0;
wire n_8988;
wire FE_RN_265_0;
wire n_5042;
wire n_13111;
wire n_44153;
wire n_21973;
wire n_14000;
wire n_6863;
wire n_2997;
wire n_19546;
wire n_6157;
wire n_24846;
wire n_40590;
wire n_19816;
wire newNet_372;
wire n_4855;
wire n_10917;
wire n_42504;
wire n_6649;
wire n_45524;
wire FE_OCP_RBN3366_n_44722;
wire n_313;
wire n_46206;
wire n_390;
wire n_8750;
wire n_3894;
wire n_47008;
wire n_6238;
wire n_5765;
wire n_7420;
wire n_30671;
wire n_31193;
wire n_26538;
wire n_6358;
wire FE_OCP_DRV_N3162_n_21419;
wire n_628;
wire n_41688;
wire n_34829;
wire n_44835;
wire FE_OCP_RBN2731_n_4219;
wire n_22987;
wire n_17709;
wire n_30602;
wire n_5141;
wire n_3189;
wire n_2258;
wire newNet_929;
wire n_40347;
wire n_8706;
wire n_29405;
wire FE_OCP_RBN2403_n_24638;
wire newNet_3364;
wire n_38022;
wire n_20150;
wire n_47004;
wire n_23499;
wire n_40523;
wire FE_RN_872_0;
wire n_7451;
wire n_40838;
wire newNet_2896;
wire n_29822;
wire newNet_536;
wire n_19959;
wire n_22235;
wire n_44776;
wire n_17126;
wire FE_RN_814_0;
wire newNet_2259;
wire n_17546;
wire n_2169;
wire newNet_2406;
wire n_17865;
wire n_8124;
wire FE_OCP_RBN2160_n_1675;
wire FE_OCP_RBN3512_n_13960;
wire n_15938;
wire newNet_2340;
wire n_28693;
wire newNet_876;
wire n_39367;
wire n_28299;
wire n_30142;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_21_;
wire n_29454;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_19_;
wire n_27480;
wire n_19471;
wire newNet_1168;
wire n_8547;
wire n_38279;
wire n_19034;
wire n_2626;
wire n_5877;
wire n_6224;
wire n_32668;
wire n_45101;
wire n_40005;
wire n_22345;
wire n_36535;
wire n_13351;
wire n_40177;
wire FE_OCP_RBN3702_n_31064;
wire n_20422;
wire newNet_1161;
wire n_12042;
wire FE_RN_47_0;
wire n_9849;
wire n_36170;
wire n_18034;
wire n_7951;
wire n_24097;
wire n_4035;
wire n_15066;
wire n_33227;
wire n_34519;
wire n_31016;
wire n_42672;
wire n_1390;
wire n_17107;
wire FE_RN_1875_0;
wire n_26308;
wire n_16611;
wire n_33933;
wire n_43125;
wire n_22068;
wire n_14531;
wire n_39584;
wire newNet_269;
wire n_30561;
wire delay_xor_ln22_unr15_stage6_stallmux_q_12_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_25_;
wire n_35592;
wire n_15048;
wire n_41158;
wire n_46944;
wire n_7860;
wire n_16674;
wire n_23072;
wire n_33827;
wire n_3352;
wire n_27867;
wire FE_RN_852_0;
wire FE_OCP_RBN3662_n_20750;
wire newNet_2248;
wire FE_RN_808_0;
wire n_37696;
wire newNet_3;
wire FE_RN_557_0;
wire n_22285;
wire n_25726;
wire n_19595;
wire n_40262;
wire n_22641;
wire n_16220;
wire n_26926;
wire n_14912;
wire n_24720;
wire n_9636;
wire n_3048;
wire n_29240;
wire FE_RN_1501_0;
wire n_35681;
wire n_41236;
wire n_8021;
wire n_14364;
wire newNet_3152;
wire n_21298;
wire n_13433;
wire n_39795;
wire n_19964;
wire n_24355;
wire n_13800;
wire n_9840;
wire n_12916;
wire n_17216;
wire n_15353;
wire n_37009;
wire n_8251;
wire n_25704;
wire FE_OCP_RBN3683_FE_RN_770_0;
wire n_14347;
wire n_5863;
wire n_22582;
wire newNet_1296;
wire n_36090;
wire n_1067;
wire n_7136;
wire n_10390;
wire newNet_964;
wire n_41434;
wire n_2142;
wire n_2059;
wire n_40251;
wire n_24271;
wire n_40995;
wire n_4568;
wire n_36287;
wire n_47260;
wire n_5134;
wire FE_RN_1650_0;
wire n_27473;
wire FE_RN_675_0;
wire n_21779;
wire n_29638;
wire n_30884;
wire n_37973;
wire n_18372;
wire n_23666;
wire n_43488;
wire n_31110;
wire n_45718;
wire n_38679;
wire n_34430;
wire n_13629;
wire FE_OCP_RBN3056_n_39913;
wire n_4507;
wire n_16890;
wire n_31638;
wire n_31681;
wire n_11723;
wire n_2953;
wire n_1402;
wire newNet_467;
wire n_36754;
wire n_22194;
wire n_4605;
wire n_21997;
wire n_14366;
wire n_20094;
wire FE_OCP_RBN1986_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_19907;
wire n_32816;
wire n_43898;
wire n_5279;
wire n_11156;
wire n_29582;
wire n_12747;
wire n_41132;
wire newNet_2732;
wire newNet_2445;
wire n_24623;
wire FE_RN_1141_0;
wire newNet_1211;
wire n_4960;
wire newNet_3528;
wire n_9564;
wire n_28941;
wire n_32866;
wire n_16345;
wire n_34011;
wire newNet_453;
wire n_514;
wire n_30933;
wire n_36314;
wire n_14431;
wire n_19286;
wire FE_RN_1837_0;
wire n_23278;
wire n_8798;
wire n_30552;
wire n_33480;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_28_;
wire n_18952;
wire n_3804;
wire n_886;
wire n_7790;
wire n_18978;
wire n_26729;
wire newNet_3121;
wire newNet_733;
wire n_39932;
wire n_8086;
wire n_36663;
wire n_23640;
wire n_2002;
wire n_21343;
wire n_11629;
wire newNet_1432;
wire n_35409;
wire FE_RN_58_0;
wire n_18734;
wire n_20197;
wire n_10549;
wire n_11229;
wire n_46235;
wire n_43644;
wire n_32519;
wire FE_OCP_RBN2271_n_13489;
wire n_32209;
wire n_39461;
wire n_15472;
wire n_42183;
wire n_3008;
wire n_2717;
wire n_29369;
wire n_42109;
wire n_19003;
wire n_30743;
wire n_21812;
wire n_17961;
wire n_22249;
wire newNet_859;
wire n_1946;
wire n_41552;
wire FE_RN_1162_0;
wire n_32712;
wire n_41826;
wire n_29102;
wire n_36466;
wire n_14025;
wire n_20811;
wire n_43771;
wire n_38102;
wire n_28948;
wire n_1040;
wire n_35365;
wire FE_OCP_RBN2172_n_32892;
wire newNet_3429;
wire n_31166;
wire n_5046;
wire delay_add_ln22_unr5_stage3_stallmux_q_1_;
wire n_18160;
wire n_38734;
wire n_25158;
wire n_26406;
wire n_22030;
wire n_7256;
wire n_23695;
wire n_29099;
wire n_33073;
wire n_36354;
wire n_7004;
wire n_13275;
wire n_21366;
wire n_30896;
wire n_329;
wire newNet_614;
wire n_12866;
wire n_20297;
wire n_21600;
wire n_10747;
wire n_2972;
wire n_27843;
wire n_7804;
wire n_22897;
wire n_39288;
wire n_12541;
wire n_2827;
wire n_7604;
wire n_37430;
wire n_26937;
wire n_40979;
wire FE_RN_55_0;
wire n_41349;
wire n_27238;
wire n_27377;
wire n_7021;
wire n_10672;
wire n_34768;
wire n_8468;
wire FE_OCP_RBN3614_n_20249;
wire FE_RN_372_0;
wire FE_RN_947_0;
wire n_35197;
wire n_7773;
wire n_32637;
wire FE_RN_101_0;
wire n_17630;
wire FE_RN_1627_0;
wire n_17336;
wire FE_OFN767_n_15670;
wire FE_OCP_RBN3525_n_29624;
wire newNet_2800;
wire n_2295;
wire FE_OCP_RBN2849_n_46982;
wire FE_OCP_DRV_N3154_n_24425;
wire n_28229;
wire n_7373;
wire n_12436;
wire n_42773;
wire FE_OCPN3169_n_23227;
wire n_11742;
wire n_26163;
wire n_10455;
wire n_16594;
wire n_19222;
wire n_41146;
wire n_32261;
wire newNet_227;
wire n_24556;
wire n_27454;
wire n_29767;
wire n_23800;
wire newNet_2960;
wire n_6653;
wire n_18441;
wire n_19564;
wire n_41365;
wire n_28348;
wire newNet_1763;
wire n_2118;
wire FE_OCP_RBN2374_n_8221;
wire n_35606;
wire n_40331;
wire n_16377;
wire n_8651;
wire n_26041;
wire n_37275;
wire n_11933;
wire n_10664;
wire n_33368;
wire n_46978;
wire n_38548;
wire FE_RN_703_0;
wire n_47340;
wire n_27094;
wire n_3264;
wire n_26955;
wire n_41281;
wire n_1499;
wire n_41671;
wire n_42024;
wire n_22850;
wire n_23769;
wire n_39570;
wire n_39217;
wire n_37020;
wire n_21518;
wire n_25677;
wire newNet_178;
wire n_24821;
wire n_29159;
wire n_36225;
wire n_34339;
wire n_9018;
wire n_3303;
wire n_22352;
wire n_40686;
wire FE_RN_1086_0;
wire n_9768;
wire n_26611;
wire n_17364;
wire n_42875;
wire n_6529;
wire n_1116;
wire n_2342;
wire n_733;
wire n_27058;
wire n_30774;
wire n_24209;
wire n_12777;
wire n_1377;
wire FE_OCP_RBN2310_n_29298;
wire n_25191;
wire FE_OCP_RBN3463_n_7886;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_14_;
wire n_15978;
wire n_31797;
wire n_30913;
wire n_10599;
wire n_30975;
wire n_26235;
wire n_33469;
wire n_40281;
wire FE_OCPN3789_n_15708;
wire n_237;
wire n_15873;
wire n_32064;
wire n_23722;
wire n_30214;
wire n_14389;
wire n_15501;
wire n_4786;
wire n_34274;
wire n_9425;
wire newNet_1233;
wire newNet_200;
wire n_42912;
wire n_9942;
wire n_27787;
wire n_26155;
wire n_36557;
wire n_8604;
wire n_42389;
wire n_785;
wire n_14303;
wire n_29079;
wire n_28659;
wire n_26682;
wire n_26584;
wire newNet_1937;
wire n_20972;
wire n_19629;
wire n_14851;
wire n_18509;
wire n_37866;
wire newNet_11;
wire n_10003;
wire n_22873;
wire n_20075;
wire n_26996;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_10_;
wire n_29663;
wire n_41052;
wire n_23607;
wire FE_OCP_RBN3830_n_19204;
wire n_16094;
wire n_20404;
wire n_7297;
wire n_31081;
wire n_1208;
wire n_17457;
wire n_18674;
wire n_12741;
wire n_31625;
wire n_13567;
wire n_32892;
wire n_34905;
wire n_14268;
wire n_44046;
wire n_23418;
wire FE_RN_832_0;
wire n_10236;
wire n_2903;
wire n_35780;
wire n_17076;
wire newNet_2941;
wire FE_RN_1621_0;
wire FE_OCP_RBN3641_n_44490;
wire n_19571;
wire n_31333;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_3_;
wire n_39416;
wire n_19681;
wire n_14146;
wire n_45214;
wire n_9909;
wire n_16401;
wire n_43265;
wire FE_RN_1773_0;
wire n_10542;
wire n_11312;
wire n_25481;
wire n_29225;
wire delay_xor_ln21_unr28_stage10_stallmux_q_2_;
wire n_7840;
wire FE_RN_556_0;
wire newNet_2166;
wire n_43444;
wire n_16600;
wire n_30283;
wire n_4121;
wire n_9608;
wire n_38493;
wire n_6407;
wire newNet_2304;
wire n_17199;
wire newNet_1945;
wire n_24735;
wire n_3910;
wire n_12462;
wire FE_RN_1844_0;
wire n_31062;
wire n_3275;
wire n_20179;
wire n_26416;
wire n_1225;
wire n_37187;
wire n_26219;
wire n_6845;
wire n_18357;
wire n_10983;
wire newNet_3412;
wire n_11455;
wire n_39164;
wire newNet_1908;
wire FE_OCP_RBN2734_n_4219;
wire n_15783;
wire n_15561;
wire n_36997;
wire newNet_27;
wire n_30847;
wire delay_add_ln22_unr17_stage7_stallmux_q_27_;
wire n_12233;
wire n_40546;
wire n_31102;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_16_;
wire n_38670;
wire n_15140;
wire n_15492;
wire n_36119;
wire n_38376;
wire n_13656;
wire n_580;
wire n_927;
wire FE_RN_1644_0;
wire n_6898;
wire n_5111;
wire n_37495;
wire n_3598;
wire n_35053;
wire n_26555;
wire FE_OCP_RBN2397_n_38586;
wire n_40238;
wire FE_OCP_DRV_N1547_n_17643;
wire n_9093;
wire n_3752;
wire n_20292;
wire n_21218;
wire n_14243;
wire FE_OFN833_n_19885;
wire n_10501;
wire n_15608;
wire FE_RN_585_0;
wire n_43618;
wire n_10828;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_27_;
wire n_20829;
wire n_10480;
wire n_34310;
wire n_7543;
wire n_12497;
wire n_35667;
wire n_45013;
wire n_25653;
wire n_23064;
wire n_203;
wire FE_OCPN3769_FE_OCP_RBN2375_n_8221;
wire FE_OFN778_n_17093;
wire n_7681;
wire n_9416;
wire n_18328;
wire n_25100;
wire n_33448;
wire n_16021;
wire n_37458;
wire n_41415;
wire n_23817;
wire n_42488;
wire n_6580;
wire n_13008;
wire n_39550;
wire n_41840;
wire n_7822;
wire n_36008;
wire n_14051;
wire n_22292;
wire newNet_782;
wire n_5070;
wire n_524;
wire n_28180;
wire n_33191;
wire n_10278;
wire n_3152;
wire newNet_816;
wire n_29042;
wire FE_OCP_RBN2315_n_41420;
wire n_24529;
wire n_10730;
wire n_30834;
wire n_38756;
wire n_26699;
wire n_3968;
wire newNet_1993;
wire n_38273;
wire n_6291;
wire n_37075;
wire n_678;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_22_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_18_;
wire n_38643;
wire n_28846;
wire FE_OCP_RBN2622_n_3601;
wire n_17995;
wire n_10834;
wire n_14737;
wire n_2360;
wire n_31354;
wire beta_23;
wire n_1362;
wire n_18863;
wire n_42333;
wire n_10841;
wire n_9011;
wire n_5417;
wire n_15841;
wire n_14614;
wire n_8319;
wire n_20463;
wire n_15339;
wire FE_OCP_RBN3675_FE_RN_1581_0;
wire n_33874;
wire n_22426;
wire n_4259;
wire FE_OCP_DRV_N1598_n_35644;
wire n_16422;
wire n_40063;
wire n_15720;
wire newNet_97;
wire n_17723;
wire n_26301;
wire newNet_650;
wire n_40886;
wire n_21152;
wire n_15773;
wire n_626;
wire n_26085;
wire n_37486;
wire FE_RN_552_0;
wire n_14069;
wire n_35253;
wire beta_10;
wire n_24142;
wire n_17859;
wire n_3428;
wire n_14780;
wire FE_OCP_RBN2131_n_32649;
wire n_7883;
wire n_33396;
wire n_26330;
wire FE_OCP_RBN2553_n_44921;
wire n_38518;
wire n_6144;
wire n_37473;
wire n_43034;
wire FE_OCPN867_n_45697;
wire n_39720;
wire newNet_831;
wire newNet_3615;
wire n_1438;
wire FE_OCP_RBN3032_n_43000;
wire n_5041;
wire newNet_2572;
wire n_365;
wire n_32877;
wire n_36779;
wire n_36894;
wire n_22670;
wire n_40743;
wire n_150;
wire n_39523;
wire FE_OCPN1473_n_24624;
wire n_30344;
wire n_26738;
wire n_15383;
wire n_24171;
wire n_25343;
wire n_2760;
wire n_14721;
wire FE_RN_1560_0;
wire newNet_278;
wire n_24019;
wire n_38238;
wire delay_xor_ln21_unr6_stage3_stallmux_q_6_;
wire n_34559;
wire n_19187;
wire n_21329;
wire n_25458;
wire n_26672;
wire n_30519;
wire n_25500;
wire n_18107;
wire n_41209;
wire n_14810;
wire n_24650;
wire n_1717;
wire n_2012;
wire n_26361;
wire FE_RN_1142_0;
wire n_10204;
wire n_25145;
wire n_17561;
wire n_41125;
wire FE_RN_1528_0;
wire n_38089;
wire n_45629;
wire n_745;
wire n_26878;
wire n_16493;
wire n_21354;
wire n_3786;
wire FE_OCPN3787_n_22156;
wire n_35948;
wire n_44222;
wire FE_RN_165_0;
wire newNet_2235;
wire n_18064;
wire n_29753;
wire n_34996;
wire n_43620;
wire n_4266;
wire FE_RN_1649_0;
wire n_32622;
wire n_41194;
wire n_26981;
wire n_34332;
wire delay_add_ln22_unr23_stage9_stallmux_q_21_;
wire n_23193;
wire n_3031;
wire n_23128;
wire newNet_3684;
wire n_18110;
wire sin_out_0;
wire n_43470;
wire FE_OCPN1858_n_22207;
wire n_10517;
wire n_41895;
wire n_42907;
wire n_16789;
wire n_20112;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_13_;
wire n_40427;
wire n_15330;
wire n_18659;
wire newNet_800;
wire n_6100;
wire n_30451;
wire newNet_1488;
wire n_39531;
wire newNet_2750;
wire n_23734;
wire n_27393;
wire newNet_3518;
wire delay_xor_ln22_unr18_stage7_stallmux_q_11_;
wire n_11385;
wire FE_RN_480_0;
wire n_38070;
wire FE_RN_1448_0;
wire FE_OCP_RBN2517_n_8762;
wire newNet_3283;
wire n_6491;
wire newNet_359;
wire n_1504;
wire n_22514;
wire n_1180;
wire n_37323;
wire n_1547;
wire n_1885;
wire n_13396;
wire n_33030;
wire newNet_3496;
wire n_3608;
wire n_3535;
wire n_13562;
wire newNet_3049;
wire FE_OCP_RBN3521_n_19663;
wire n_19608;
wire n_22370;
wire n_21593;
wire n_25394;
wire FE_RN_46_0;
wire newNet_406;
wire n_4686;
wire n_25690;
wire delay_xor_ln22_unr15_stage6_stallmux_q_9_;
wire n_15536;
wire n_9652;
wire newNet_1024;
wire n_5199;
wire n_42995;
wire n_3209;
wire n_16940;
wire n_18247;
wire n_19768;
wire n_33986;
wire n_40783;
wire n_11284;
wire n_37164;
wire n_2288;
wire FE_OCPN1243_n_44460;
wire n_41615;
wire n_12091;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_30_;
wire n_33098;
wire n_26343;
wire n_33016;
wire n_35750;
wire n_42249;
wire n_1958;
wire n_556;
wire n_18918;
wire n_11944;
wire newNet_1242;
wire n_12925;
wire FE_OCP_RBN2651_n_9030;
wire n_8399;
wire n_22859;
wire n_17498;
wire n_31940;
wire n_38262;
wire FE_RN_212_0;
wire n_1533;
wire n_19296;
wire n_27441;
wire n_1140;
wire n_16266;
wire n_26711;
wire n_39189;
wire n_20023;
wire n_36541;
wire n_26894;
wire n_519;
wire cos_out_0;
wire n_26748;
wire n_15053;
wire n_38925;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_9_;
wire n_33046;
wire n_38534;
wire n_10083;
wire n_28238;
wire n_37827;
wire n_23680;
wire n_43864;
wire newNet_1012;
wire n_31571;
wire n_22796;
wire n_23613;
wire FE_OCP_RBN2914_n_42947;
wire n_5530;
wire n_43690;
wire n_12240;
wire n_37678;
wire FE_RN_242_0;
wire FE_OFN797_n_46285;
wire n_22164;
wire n_18171;
wire n_20979;
wire n_27991;
wire n_43381;
wire n_16864;
wire n_40449;
wire FE_OCP_RBN3696_n_5284;
wire n_43343;
wire newNet_2184;
wire n_34575;
wire n_27497;
wire n_16876;
wire FE_OCP_RBN2539_n_8781;
wire n_33768;
wire n_6026;
wire n_28957;
wire FE_RN_282_0;
wire n_35321;
wire n_29441;
wire n_27001;
wire n_28987;
wire n_25070;
wire n_1356;
wire n_11809;
wire newNet_3556;
wire n_37710;
wire n_42106;
wire n_2561;
wire n_14629;
wire n_23182;
wire n_16583;
wire n_20987;
wire FE_OCP_RBN1345_n_19270;
wire n_7273;
wire FE_OCP_RBN2857_n_10399;
wire n_30368;
wire n_26769;
wire n_17488;
wire n_11973;
wire n_28934;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_16_;
wire n_26405;
wire n_37394;
wire n_36971;
wire n_15112;
wire n_33540;
wire FE_RN_525_0;
wire n_6652;
wire n_7651;
wire n_14561;
wire n_17892;
wire n_21399;
wire n_16319;
wire n_37985;
wire newNet_847;
wire n_35232;
wire n_11247;
wire n_7066;
wire n_43139;
wire n_5943;
wire FE_RN_121_0;
wire n_42861;
wire FE_OCP_RBN3592_n_8902;
wire delay_xor_ln22_unr9_stage4_stallmux_q_12_;
wire n_28974;
wire n_28712;
wire n_17479;
wire n_25282;
wire n_4548;
wire n_13863;
wire n_5606;
wire n_29900;
wire n_30805;
wire n_36399;
wire newNet_1786;
wire FE_RN_346_0;
wire n_17886;
wire n_18642;
wire n_21897;
wire n_43020;
wire FE_OCPN853_n_45450;
wire n_44311;
wire n_7146;
wire n_44265;
wire n_7508;
wire n_22032;
wire n_6112;
wire n_19096;
wire n_13381;
wire n_6681;
wire n_10890;
wire n_37310;
wire FE_OCP_RBN2247_n_13017;
wire FE_OCP_RBN2290_n_2438;
wire n_425;
wire n_17628;
wire n_18089;
wire n_11956;
wire n_46378;
wire n_36914;
wire FE_RN_1170_0;
wire newNet_1317;
wire n_13816;
wire n_1668;
wire n_45530;
wire newNet_505;
wire n_39993;
wire n_28014;
wire n_5159;
wire n_38632;
wire n_47197;
wire n_17386;
wire n_38211;
wire n_14719;
wire n_5233;
wire newNet_445;
wire FE_RN_1177_0;
wire n_10707;
wire n_906;
wire newNet_2634;
wire n_13355;
wire cos_out_22;
wire n_28826;
wire n_6690;
wire n_13491;
wire n_33684;
wire n_34739;
wire n_15181;
wire n_13324;
wire n_837;
wire n_37514;
wire n_27825;
wire n_38320;
wire n_27318;
wire n_15526;
wire n_34580;
wire FE_RN_640_0;
wire n_38683;
wire FE_RN_1038_0;
wire n_33969;
wire n_18541;
wire n_29514;
wire n_33181;
wire n_5242;
wire n_18550;
wire n_2093;
wire FE_OCP_RBN2770_n_9892;
wire n_23301;
wire n_36035;
wire n_41243;
wire n_7417;
wire n_20204;
wire n_24391;
wire sin_out_10;
wire n_42669;
wire n_14792;
wire n_8002;
wire n_20995;
wire n_1515;
wire n_162;
wire n_21186;
wire n_32914;
wire n_9836;
wire newNet_1493;
wire n_19688;
wire n_40092;
wire n_43269;
wire newNet_2160;
wire n_895;
wire n_16923;
wire n_29020;
wire n_6179;
wire n_41277;
wire delay_add_ln22_unr23_stage9_stallmux_q_29_;
wire n_5033;
wire n_16488;
wire n_12377;
wire n_27950;
wire n_5438;
wire n_36124;
wire n_34305;
wire FE_OCP_RBN2400_n_2885;
wire n_35042;
wire n_2873;
wire n_7191;
wire n_33580;
wire n_6205;
wire FE_RN_1636_0;
wire n_32313;
wire n_42287;
wire n_21742;
wire n_5441;
wire n_35272;
wire n_32429;
wire n_27813;
wire n_40925;
wire n_9379;
wire n_41831;
wire n_18234;
wire n_261;
wire n_4098;
wire newNet_960;
wire n_6067;
wire n_37979;
wire n_3941;
wire n_21688;
wire n_35130;
wire n_8211;
wire n_10909;
wire FE_OCPN1756_n_16923;
wire n_64;
wire n_39342;
wire n_5509;
wire n_12882;
wire newNet_3004;
wire n_16722;
wire n_26114;
wire n_35437;
wire n_6555;
wire newNet_3422;
wire n_40229;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_29_;
wire n_9495;
wire n_33846;
wire newNet_3148;
wire n_2243;
wire n_16641;
wire FE_RN_1135_0;
wire n_32337;
wire n_42078;
wire n_45861;
wire n_35599;
wire FE_RN_788_0;
wire delay_sub_ln23_0_unr24_stage9_stallmux_q;
wire n_10492;
wire n_30636;
wire n_4104;
wire n_25634;
wire n_24979;
wire newNet_2947;
wire n_5342;
wire n_5987;
wire n_28452;
wire n_37093;
wire n_2379;
wire n_7869;
wire n_6933;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_31_;
wire newNet_1934;
wire n_39405;
wire n_19110;
wire n_14650;
wire n_19217;
wire n_10920;
wire FE_RN_1066_0;
wire n_19308;
wire n_41952;
wire n_30697;
wire n_27083;
wire n_40817;
wire n_9560;
wire n_12036;
wire n_18892;
wire n_40437;
wire n_36693;
wire n_14581;
wire newNet_348;
wire n_24585;
wire n_29648;
wire FE_OCP_RBN2284_n_33846;
wire n_20129;
wire n_13555;
wire n_9417;
wire newNet_2054;
wire n_24169;
wire n_38566;
wire FE_RN_1283_0;
wire n_35246;
wire n_6465;
wire FE_OCPN1470_n_23818;
wire n_10292;
wire n_44652;
wire n_1009;
wire n_18348;
wire n_44763;
wire n_31276;
wire n_23226;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_1_;
wire n_5235;
wire n_22296;
wire newNet_1617;
wire n_23346;
wire n_22848;
wire n_30662;
wire n_10228;
wire n_38247;
wire n_17496;
wire n_39660;
wire n_23945;
wire n_10040;
wire newNet_2903;
wire n_19077;
wire n_25945;
wire n_41594;
wire n_4119;
wire n_6901;
wire n_41936;
wire FE_RN_243_0;
wire n_22187;
wire n_103;
wire n_9195;
wire n_3217;
wire n_30359;
wire newNet_1544;
wire n_13517;
wire n_13135;
wire n_12094;
wire n_42271;
wire n_15459;
wire newNet_1694;
wire n_6878;
wire n_29176;
wire newNet_1228;
wire n_12030;
wire newNet_2838;
wire n_23106;
wire FE_OCP_RBN3567_n_29857;
wire n_23830;
wire n_12808;
wire n_25063;
wire n_43586;
wire n_9004;
wire newNet_379;
wire n_32439;
wire n_22623;
wire n_26246;
wire n_3637;
wire n_21788;
wire FE_OCP_RBN2860_n_10399;
wire FE_OCP_RBN2116_n_45224;
wire newNet_921;
wire newNet_3490;
wire n_22646;
wire n_33381;
wire n_949;
wire n_33315;
wire n_17683;
wire n_22227;
wire n_41008;
wire n_26622;
wire n_24052;
wire n_30888;
wire n_9274;
wire n_41904;
wire n_20163;
wire n_2197;
wire n_34346;
wire n_42302;
wire n_37882;
wire n_3492;
wire n_32992;
wire FE_RN_906_0;
wire n_32764;
wire n_39857;
wire n_6990;
wire n_13464;
wire n_8368;
wire n_29382;
wire n_2512;
wire n_9984;
wire FE_RN_117_0;
wire n_9894;
wire newNet_3351;
wire n_4442;
wire n_22717;
wire n_40892;
wire n_1089;
wire newNet_2020;
wire n_13131;
wire n_19478;
wire n_40946;
wire newNet_2013;
wire n_17477;
wire n_5365;
wire FE_RN_1731_0;
wire n_35919;
wire n_38589;
wire n_37535;
wire n_40392;
wire n_35842;
wire n_9618;
wire n_20619;
wire n_12816;
wire n_21252;
wire n_39333;
wire n_18716;
wire FE_RN_1588_0;
wire FE_OCP_RBN3108_n_40586;
wire n_46210;
wire n_9452;
wire n_30030;
wire n_9079;
wire n_18946;
wire n_14126;
wire n_41481;
wire newNet_1015;
wire n_25754;
wire n_37408;
wire n_10247;
wire FE_OCPN1021_n_23195;
wire n_10557;
wire n_29937;
wire n_16767;
wire n_27639;
wire n_13578;
wire n_4731;
wire n_41223;
wire n_20848;
wire n_37587;
wire n_19070;
wire n_5394;
wire n_11058;
wire n_23759;
wire n_19491;
wire n_31232;
wire n_13080;
wire n_4579;
wire n_27542;
wire n_37233;
wire n_4046;
wire n_42525;
wire n_39330;
wire FE_RN_394_0;
wire n_5123;
wire n_36708;
wire n_33323;
wire n_1768;
wire n_31175;
wire n_13010;
wire n_13554;
wire n_7611;
wire n_11695;
wire n_19531;
wire n_37254;
wire n_11036;
wire n_24936;
wire n_24500;
wire n_26105;
wire n_21423;
wire n_8434;
wire n_32597;
wire n_22086;
wire n_25561;
wire n_14923;
wire n_6966;
wire n_32888;
wire n_12490;
wire n_28365;
wire n_27690;
wire FE_RN_858_0;
wire n_9218;
wire n_10572;
wire FE_OCP_RBN3308_n_44722;
wire n_14297;
wire n_28615;
wire n_38112;
wire n_13045;
wire n_24537;
wire n_42235;
wire n_14657;
wire n_28257;
wire n_11530;
wire n_20216;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_26_;
wire newNet_1593;
wire n_43422;
wire n_17261;
wire FE_RN_1333_0;
wire n_29223;
wire n_39589;
wire n_13262;
wire n_40694;
wire FE_RN_880_0;
wire newNet_1631;
wire n_26835;
wire n_13751;
wire FE_RN_1770_0;
wire n_17393;
wire n_30191;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_4_;
wire n_25939;
wire newNet_1158;
wire n_39630;
wire n_26758;
wire n_16168;
wire n_11082;
wire n_1085;
wire FE_RN_1786_0;
wire n_32219;
wire n_44437;
wire n_31545;
wire n_8536;
wire n_17045;
wire n_36486;
wire n_23768;
wire n_19875;
wire n_12195;
wire n_12947;
wire n_43142;
wire n_31447;
wire n_43427;
wire n_37777;
wire n_14492;
wire n_26258;
wire newNet_2727;
wire FE_OCP_RBN1144_n_29292;
wire n_26656;
wire n_9967;
wire n_35509;
wire delay_xor_ln21_unr15_stage6_stallmux_q_13_;
wire n_36886;
wire FE_RN_374_0;
wire n_28549;
wire delay_sub_ln23_0_unr27_stage10_stallmux_z;
wire FE_OCP_RBN3095_n_11413;
wire n_13078;
wire n_15838;
wire n_14704;
wire newNet_3716;
wire n_5726;
wire n_42285;
wire n_10419;
wire n_8962;
wire n_33178;
wire n_40466;
wire n_29531;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_25_;
wire delay_add_ln22_unr8_stage4_stallmux_q_11_;
wire n_17032;
wire n_14884;
wire n_23849;
wire newNet_3673;
wire newNet_1927;
wire n_2750;
wire n_22132;
wire n_13893;
wire newNet_559;
wire n_34678;
wire n_5084;
wire FE_RN_244_0;
wire n_16699;
wire newNet_2982;
wire n_13753;
wire n_608;
wire n_5617;
wire n_17346;
wire newNet_1961;
wire n_12719;
wire n_30713;
wire n_38891;
wire n_6995;
wire n_30172;
wire n_28357;
wire n_31637;
wire n_26190;
wire n_20771;
wire n_34288;
wire newNet_3584;
wire n_7596;
wire n_15376;
wire n_11866;
wire n_34434;
wire newNet_1073;
wire n_41532;
wire newNet_1381;
wire n_4787;
wire n_25554;
wire n_19081;
wire n_35926;
wire n_11704;
wire n_43794;
wire n_17595;
wire newNet_2571;
wire n_21553;
wire n_31607;
wire n_39037;
wire FE_OCP_RBN2440_n_8402;
wire n_37195;
wire n_25644;
wire n_28922;
wire n_16753;
wire n_19449;
wire n_14731;
wire n_27167;
wire n_10318;
wire n_41299;
wire n_42395;
wire FE_OCP_RBN3623_n_39097;
wire n_44825;
wire newNet_769;
wire n_601;
wire newNet_2148;
wire n_31874;
wire n_38623;
wire n_40016;
wire n_13696;
wire n_33338;
wire n_8238;
wire n_14504;
wire n_26819;
wire n_42728;
wire n_33869;
wire delay_xor_ln21_unr12_stage5_stallmux_q_18_;
wire newNet_3060;
wire n_38504;
wire FE_OCP_RBN3452_n_37945;
wire FE_RN_1763_0;
wire n_8470;
wire n_12314;
wire n_40285;
wire n_3291;
wire n_20384;
wire n_332;
wire n_9642;
wire n_33923;
wire n_42266;
wire n_16233;
wire n_1736;
wire n_12253;
wire n_31428;
wire n_23271;
wire FE_OCP_RBN2850_n_46982;
wire n_13806;
wire n_19832;
wire newNet_1110;
wire n_28434;
wire n_14748;
wire n_38717;
wire FE_RN_1579_0;
wire n_43376;
wire n_5570;
wire n_28586;
wire n_10770;
wire delay_xor_ln21_unr6_stage3_stallmux_q_4_;
wire n_24902;
wire n_15391;
wire FE_OCP_RBN2274_n_2457;
wire n_3562;
wire newNet_2796;
wire newNet_883;
wire FE_RN_550_0;
wire n_14253;
wire n_4777;
wire n_5515;
wire n_23630;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_7_;
wire n_14308;
wire newNet_261;
wire n_23250;
wire n_2914;
wire n_7084;
wire n_24310;
wire n_38268;
wire n_1834;
wire n_18838;
wire n_7575;
wire newNet_29;
wire n_24381;
wire FE_RN_1556_0;
wire n_35201;
wire n_28292;
wire n_6056;
wire n_28310;
wire n_10613;
wire n_28587;
wire n_44;
wire n_37981;
wire n_1700;
wire n_8196;
wire n_24056;
wire n_26452;
wire n_32457;
wire n_34579;
wire n_37606;
wire n_24652;
wire FE_OCP_RBN2370_n_38545;
wire n_16074;
wire n_15075;
wire n_18025;
wire n_37625;
wire FE_OCP_RBN2189_n_7346;
wire n_15378;
wire n_27382;
wire n_23825;
wire n_12708;
wire n_14466;
wire n_41927;
wire newNet_1555;
wire n_36656;
wire n_21925;
wire n_28650;
wire FE_OCP_RBN3581_n_44944;
wire FE_OCP_RBN3138_n_40568;
wire n_36686;
wire FE_RN_1009_0;
wire n_19470;
wire n_36560;
wire n_42808;
wire n_18626;
wire n_21437;
wire n_41168;
wire n_18852;
wire n_27911;
wire n_25729;
wire n_4468;
wire n_3953;
wire n_39434;
wire n_38991;
wire n_22881;
wire n_43280;
wire n_41987;
wire n_25640;
wire FE_OCP_RBN2639_n_38806;
wire n_13854;
wire FE_OCP_RBN2185_FE_RN_464_0;
wire n_34696;
wire n_11751;
wire n_33614;
wire delay_xor_ln21_unr6_stage3_stallmux_q_5_;
wire n_34757;
wire n_36766;
wire n_29196;
wire n_11630;
wire n_16368;
wire FE_OCP_RBN1372_n_35275;
wire n_334;
wire n_257;
wire FE_OCPN1235_n_32791;
wire n_35329;
wire n_37055;
wire newNet_975;
wire FE_OCP_RBN2230_n_13141;
wire n_14411;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_19_;
wire n_38687;
wire n_7236;
wire n_2215;
wire FE_RN_300_0;
wire n_36880;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_11_;
wire n_25089;
wire n_8731;
wire n_437;
wire FE_OCP_RBN2391_n_19434;
wire n_33559;
wire n_34506;
wire n_12517;
wire n_1801;
wire n_5058;
wire n_1521;
wire n_13907;
wire n_4459;
wire n_16603;
wire FE_RN_785_0;
wire n_33028;
wire FE_OCPN1857_n_22207;
wire n_12742;
wire n_11524;
wire n_35932;
wire newNet_1135;
wire n_15530;
wire n_29255;
wire FE_OCP_RBN2917_n_10644;
wire n_26957;
wire n_15361;
wire n_31096;
wire n_37047;
wire n_14190;
wire n_25301;
wire n_23809;
wire newNet_743;
wire n_30590;
wire n_38658;
wire n_2501;
wire n_8282;
wire n_9767;
wire n_39873;
wire n_45897;
wire n_36803;
wire n_658;
wire n_25993;
wire newNet_1250;
wire n_16019;
wire n_1211;
wire n_37123;
wire n_29316;
wire n_22633;
wire n_26480;
wire n_30462;
wire FE_OCPN932_n_40736;
wire n_36192;
wire FE_OCP_RBN2331_n_29353;
wire FE_OCP_RBN3821_n_44061;
wire newNet_3038;
wire n_18083;
wire n_18580;
wire n_618;
wire n_23651;
wire n_28074;
wire n_14672;
wire n_17938;
wire n_11553;
wire n_8062;
wire n_10353;
wire n_32392;
wire n_3660;
wire n_36487;
wire n_32440;
wire n_31549;
wire n_34629;
wire n_40961;
wire n_14068;
wire n_30194;
wire n_12489;
wire n_36528;
wire n_12571;
wire n_16159;
wire n_39861;
wire FE_RN_1843_0;
wire n_21711;
wire FE_OCP_RBN3694_n_26409;
wire n_40301;
wire n_13542;
wire newNet_1344;
wire n_32463;
wire n_20686;
wire n_9064;
wire n_18224;
wire n_22410;
wire delay_add_ln22_unr2_stage2_stallmux_q_22_;
wire newNet_2827;
wire n_38116;
wire n_23506;
wire n_22055;
wire FE_OCP_RBN3562_n_29857;
wire n_22555;
wire n_25460;
wire n_19610;
wire n_13549;
wire n_22594;
wire n_25110;
wire n_17846;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_23_;
wire n_43170;
wire n_6908;
wire n_4559;
wire n_46985;
wire n_16023;
wire n_15761;
wire n_35449;
wire n_5050;
wire n_21703;
wire n_7299;
wire n_19425;
wire n_31386;
wire FE_OCP_RBN2479_n_8530;
wire n_7927;
wire n_19911;
wire n_3993;
wire n_9330;
wire n_22748;
wire n_1696;
wire n_11103;
wire n_35883;
wire n_9728;
wire FE_OCP_RBN2876_n_10354;
wire n_26646;
wire n_30502;
wire n_42975;
wire n_6591;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_20_;
wire newNet_187;
wire n_15407;
wire n_35638;
wire n_12551;
wire n_39200;
wire delay_xor_ln21_unr18_stage7_stallmux_q_9_;
wire n_11316;
wire n_42211;
wire n_46172;
wire n_34414;
wire newNet_2203;
wire n_3503;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_11_;
wire newNet_3083;
wire n_18579;
wire n_31229;
wire FE_OCP_RBN1202_n_25898;
wire n_18326;
wire n_13416;
wire n_865;
wire n_23578;
wire n_37799;
wire newNet_2741;
wire n_24256;
wire n_24702;
wire n_36594;
wire FE_OCP_RBN1185_n_14823;
wire n_15467;
wire n_7663;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_6_;
wire n_31157;
wire n_25044;
wire n_5920;
wire n_10753;
wire n_21727;
wire n_31885;
wire n_17311;
wire n_14976;
wire n_41986;
wire n_1968;
wire n_26629;
wire n_38064;
wire n_1537;
wire FE_OCPN1504_n_47257;
wire newNet_1859;
wire n_16713;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_25_;
wire n_42194;
wire n_15827;
wire n_12086;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_23_;
wire n_7431;
wire newNet_895;
wire n_5621;
wire n_38191;
wire n_14221;
wire n_31720;
wire n_46950;
wire n_4006;
wire n_31852;
wire n_6187;
wire n_42448;
wire n_37437;
wire n_12558;
wire n_30738;
wire n_43533;
wire n_10065;
wire n_21766;
wire n_29410;
wire n_34230;
wire n_33695;
wire n_31585;
wire n_6666;
wire newNet_2807;
wire newNet_2423;
wire n_8069;
wire FE_OCP_RBN2739_n_20432;
wire n_11211;
wire n_1427;
wire n_16911;
wire n_32839;
wire newNet_1830;
wire n_34550;
wire n_10422;
wire n_2207;
wire n_46416;
wire newNet_1449;
wire FE_OCP_RBN3121_n_32239;
wire n_6971;
wire n_37901;
wire n_23228;
wire n_12513;
wire n_35050;
wire newNet_324;
wire n_6104;
wire newNet_222;
wire n_39304;
wire n_24188;
wire FE_OCPN1259_n_25353;
wire n_31740;
wire FE_RN_1451_0;
wire n_1439;
wire delay_add_ln22_unr17_stage7_stallmux_q_2_;
wire FE_OCPN3746_n_29439;
wire n_41807;
wire n_3041;
wire FE_OCPN1418_n_31504;
wire n_24016;
wire n_36383;
wire n_10309;
wire n_19044;
wire n_42069;
wire n_16194;
wire newNet_289;
wire n_33455;
wire n_35422;
wire n_7900;
wire n_41166;
wire n_28533;
wire FE_OCPN3770_n_8669;
wire n_23858;
wire n_36403;
wire n_1170;
wire n_12631;
wire n_18839;
wire n_31441;
wire n_12855;
wire FE_RN_21_0;
wire n_39107;
wire n_28682;
wire n_43324;
wire n_28232;
wire delay_add_ln22_unr14_stage6_stallmux_q_4_;
wire n_2297;
wire n_41764;
wire n_41875;
wire n_26118;
wire n_43572;
wire FE_OCP_RBN3583_n_9245;
wire n_13520;
wire n_32626;
wire n_28764;
wire n_33826;
wire n_5494;
wire FE_OCP_RBN3469_n_7886;
wire newNet_2935;
wire n_38141;
wire n_9572;
wire n_32988;
wire n_320;
wire n_22538;
wire n_26726;
wire n_36814;
wire n_3795;
wire n_47018;
wire newNet_3372;
wire n_34221;
wire n_33780;
wire n_30902;
wire n_14643;
wire FE_OCP_RBN2749_n_9629;
wire newNet_2866;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_26_;
wire newNet_2705;
wire newNet_655;
wire n_2895;
wire n_28460;
wire n_43653;
wire n_1001;
wire n_41780;
wire FE_OCP_RBN1379_n_20732;
wire n_10374;
wire n_8105;
wire FE_RN_792_0;
wire n_16390;
wire n_21852;
wire n_36780;
wire n_9743;
wire n_32574;
wire n_15999;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_19_;
wire n_4773;
wire n_16072;
wire n_1646;
wire n_27976;
wire n_5894;
wire FE_OCP_RBN1197_n_30619;
wire n_32802;
wire n_37279;
wire n_30168;
wire n_33722;
wire n_4246;
wire delay_add_ln22_unr8_stage4_stallmux_q_28_;
wire FE_RN_468_0;
wire n_39959;
wire FE_RN_647_0;
wire n_4016;
wire n_39468;
wire FE_OFN762_n_15670;
wire n_42428;
wire n_15714;
wire n_36869;
wire newNet_632;
wire delay_xor_ln22_unr15_stage6_stallmux_q_15_;
wire FE_OCP_RBN2641_n_34921;
wire n_24433;
wire FE_OCPN1042_n_3673;
wire n_24473;
wire n_31785;
wire n_22942;
wire n_43598;
wire n_42628;
wire FE_RN_1565_0;
wire n_22502;
wire n_43558;
wire n_33732;
wire newNet_1106;
wire n_43412;
wire n_42693;
wire newNet_2286;
wire n_34389;
wire n_9525;
wire n_17406;
wire n_42437;
wire FE_RN_1200_0;
wire delay_add_ln22_unr8_stage4_stallmux_q_25_;
wire n_36668;
wire delay_add_ln22_unr8_stage4_stallmux_q_19_;
wire n_9298;
wire n_8989;
wire n_15455;
wire newNet_866;
wire n_17617;
wire n_7601;
wire n_20181;
wire n_42687;
wire n_42340;
wire newNet_2087;
wire n_26051;
wire n_28279;
wire delay_xor_ln22_unr6_stage3_stallmux_q_19_;
wire n_22842;
wire n_2727;
wire n_4199;
wire n_19196;
wire n_28407;
wire newNet_775;
wire n_18203;
wire n_28552;
wire n_36295;
wire n_4511;
wire n_20183;
wire n_32373;
wire n_42983;
wire FE_OCP_RBN3455_FE_OCPN1240_n_7721;
wire n_41456;
wire n_5556;
wire n_26630;
wire n_3577;
wire newNet_1958;
wire n_22729;
wire n_2320;
wire FE_RN_249_0;
wire n_26812;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_8_;
wire n_1876;
wire n_27217;
wire n_29081;
wire n_34881;
wire n_22238;
wire n_36180;
wire n_36320;
wire n_32962;
wire n_4821;
wire n_14854;
wire n_47184;
wire n_31650;
wire FE_RN_983_0;
wire n_5095;
wire n_35021;
wire n_33535;
wire n_32395;
wire newNet_3247;
wire n_24306;
wire FE_RN_80_0;
wire n_29850;
wire newNet_1355;
wire n_18611;
wire n_5766;
wire n_11511;
wire n_40355;
wire delay_sub_ln21_unr24_stage9_stallmux_q_3_;
wire n_45008;
wire newNet_717;
wire n_32533;
wire newNet_2779;
wire n_30979;
wire n_40529;
wire n_11560;
wire n_34248;
wire n_37972;
wire FE_OCP_RBN3465_n_7886;
wire n_2491;
wire n_39985;
wire n_7524;
wire n_28570;
wire n_492;
wire n_13717;
wire n_29783;
wire newNet_991;
wire n_9675;
wire n_12391;
wire n_32052;
wire newNet_622;
wire n_20060;
wire n_13504;
wire n_44147;
wire n_28317;
wire n_45331;
wire newNet_3426;
wire n_3063;
wire n_24667;
wire n_6540;
wire n_21774;
wire n_33200;
wire n_25527;
wire n_32727;
wire n_7269;
wire n_23080;
wire newNet_402;
wire n_41709;
wire newNet_1736;
wire n_24747;
wire n_37690;
wire n_45865;
wire newNet_756;
wire n_26101;
wire n_28210;
wire n_30364;
wire n_33185;
wire n_9144;
wire n_11334;
wire n_23188;
wire beta_28;
wire n_1245;
wire n_1998;
wire newNet_1008;
wire n_33103;
wire n_32333;
wire n_31500;
wire newNet_2884;
wire delay_add_ln22_unr23_stage9_stallmux_q_8_;
wire n_38469;
wire n_14890;
wire FE_RN_928_0;
wire n_10977;
wire n_9554;
wire n_3392;
wire FE_OCP_RBN2358_n_13818;
wire n_24446;
wire newNet_1609;
wire newNet_1205;
wire n_26913;
wire n_18267;
wire n_6387;
wire n_13053;
wire n_40321;
wire n_20537;
wire n_20671;
wire n_13366;
wire n_1720;
wire n_40746;
wire FE_RN_271_0;
wire n_5313;
wire n_41816;
wire n_3320;
wire n_38347;
wire n_39485;
wire n_6567;
wire n_38514;
wire n_4280;
wire n_6282;
wire n_27158;
wire newNet_3477;
wire FE_RN_570_0;
wire FE_OCP_RBN3580_n_44944;
wire n_29724;
wire FE_OCP_RBN2605_FE_OCPN899_n_44593;
wire n_5529;
wire n_41341;
wire n_16328;
wire n_19797;
wire n_6321;
wire n_2180;
wire n_35654;
wire n_18128;
wire n_35337;
wire n_39864;
wire n_40893;
wire n_10863;
wire n_14588;
wire FE_RN_1723_0;
wire n_8685;
wire n_16828;
wire n_12285;
wire n_42280;
wire n_9232;
wire FE_OFN842_n_5067;
wire n_40653;
wire newNet_2379;
wire n_11955;
wire n_1193;
wire n_28969;
wire newNet_292;
wire n_11174;
wire FE_OCPN3164_n_24117;
wire n_38118;
wire n_4716;
wire n_32380;
wire n_39400;
wire FE_RN_1694_0;
wire FE_RN_1721_0;
wire n_23009;
wire n_19944;
wire n_16200;
wire n_2366;
wire newNet_3710;
wire n_9935;
wire n_19141;
wire n_33939;
wire FE_OCP_RBN1179_n_18981;
wire n_29844;
wire newNet_1515;
wire n_27505;
wire FE_OCP_RBN2638_n_38806;
wire n_37529;
wire n_9132;
wire n_23754;
wire n_41513;
wire n_1056;
wire n_14423;
wire n_29748;
wire n_21289;
wire FE_OCP_RBN2164_n_28249;
wire n_13017;
wire n_24028;
wire newNet_2486;
wire n_26641;
wire n_11816;
wire n_34490;
wire n_9830;
wire n_3932;
wire n_20720;
wire n_34954;
wire n_10587;
wire FE_OCP_RBN3470_n_7886;
wire n_13992;
wire n_14164;
wire n_8454;
wire n_9214;
wire n_25619;
wire n_40904;
wire n_1037;
wire n_25180;
wire n_6280;
wire n_16364;
wire n_4287;
wire n_26677;
wire newNet_3441;
wire n_14078;
wire n_34824;
wire n_16985;
wire FE_OFN345_n_9247;
wire FE_OCP_RBN2827_FE_RN_1573_0;
wire n_43159;
wire newNet_791;
wire FE_RN_1767_0;
wire n_19517;
wire FE_OCP_RBN1194_n_22542;
wire n_6149;
wire n_33324;
wire n_14565;
wire FE_OCP_RBN3462_n_7886;
wire n_18287;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_0_;
wire n_41382;
wire FE_OCPN1787_n_36034;
wire n_39791;
wire n_31190;
wire n_33912;
wire n_35108;
wire n_36638;
wire n_43823;
wire n_35137;
wire n_28362;
wire FE_OCPN3754_n_1451;
wire n_23565;
wire n_2255;
wire n_3172;
wire n_2530;
wire n_13607;
wire n_19819;
wire n_3322;
wire n_10479;
wire n_665;
wire n_35488;
wire n_21528;
wire n_31302;
wire n_42704;
wire n_16111;
wire newNet_1470;
wire n_3692;
wire FE_OCPUNCON1801_n_29375;
wire delay_sub_ln22_unr24_stage9_stallmux_q_3_;
wire n_27305;
wire newNet_2100;
wire n_13771;
wire FE_OCP_RBN2730_n_4219;
wire n_9243;
wire n_7673;
wire newNet_798;
wire n_10016;
wire n_11658;
wire n_19701;
wire n_45319;
wire n_22908;
wire n_23934;
wire n_8133;
wire newNet_2617;
wire n_11971;
wire n_16630;
wire n_41755;
wire n_1121;
wire n_13076;
wire newNet_1333;
wire n_27021;
wire n_46146;
wire n_12342;
wire n_42843;
wire FE_RN_1060_0;
wire n_26776;
wire n_4903;
wire n_5970;
wire n_7910;
wire n_28616;
wire n_4751;
wire n_17981;
wire n_39054;
wire FE_OCP_RBN3102_n_27571;
wire n_22762;
wire n_39079;
wire FE_RN_521_0;
wire n_16086;
wire n_30825;
wire n_5016;
wire n_2537;
wire n_15087;
wire n_325;
wire n_312;
wire n_6311;
wire n_7195;
wire FE_OCP_RBN3385_n_33108;
wire n_5255;
wire n_10591;
wire n_8520;
wire FE_RN_1826_0;
wire n_13154;
wire newNet_2541;
wire n_43738;
wire FE_RN_1403_0;
wire delay_add_ln22_unr11_stage5_stallmux_q_27_;
wire n_18678;
wire n_11187;
wire n_12373;
wire n_34219;
wire n_43605;
wire n_32862;
wire n_46362;
wire FE_OCP_RBN3211_n_44365;
wire newNet_1230;
wire n_14733;
wire n_37103;
wire n_32432;
wire n_2356;
wire n_4178;
wire n_19842;
wire n_27416;
wire n_19877;
wire n_7180;
wire n_7864;
wire n_38185;
wire newNet_542;
wire n_31912;
wire n_15420;
wire n_39627;
wire n_37525;
wire n_10916;
wire n_34899;
wire n_34326;
wire n_6644;
wire n_13087;
wire newNet_107;
wire n_17290;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_10_;
wire n_23179;
wire n_29672;
wire n_42507;
wire n_1689;
wire n_29391;
wire n_36969;
wire n_34976;
wire n_28860;
wire n_12842;
wire n_33343;
wire newNet_3594;
wire n_25870;
wire n_31376;
wire n_34117;
wire n_25347;
wire n_19543;
wire n_37702;
wire FE_OCP_RBN2858_n_10399;
wire n_51;
wire n_39452;
wire n_2891;
wire FE_OCPN989_n_28353;
wire n_20783;
wire newNet_1191;
wire FE_RN_1504_0;
wire n_9962;
wire n_40373;
wire n_20614;
wire n_23746;
wire n_33504;
wire newNet_822;
wire n_42049;
wire n_22827;
wire n_46350;
wire n_11633;
wire n_38454;
wire n_7157;
wire n_29309;
wire n_31960;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_13_;
wire newNet_2279;
wire n_34565;
wire n_31056;
wire n_4539;
wire n_35873;
wire newNet_603;
wire n_18492;
wire newNet_3574;
wire delay_xor_ln21_unr12_stage5_stallmux_q_15_;
wire n_34864;
wire n_18073;
wire FE_RN_862_0;
wire newNet_1569;
wire n_3559;
wire n_34811;
wire n_4278;
wire sin_out_13;
wire n_18869;
wire n_15652;
wire newNet_118;
wire n_32509;
wire n_632;
wire newNet_1479;
wire n_31731;
wire n_46153;
wire n_26079;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_14_;
wire n_30653;
wire n_18293;
wire n_17940;
wire n_1987;
wire n_17527;
wire n_1220;
wire n_5203;
wire n_33127;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_25_;
wire n_42938;
wire n_39580;
wire n_38509;
wire FE_OCP_RBN3410_n_45120;
wire n_915;
wire n_20806;
wire n_25109;
wire n_15751;
wire n_4935;
wire n_37650;
wire n_17927;
wire newNet_2173;
wire FE_OCP_RBN2127_n_6745;
wire newNet_3657;
wire n_17827;
wire n_21237;
wire n_21319;
wire n_25799;
wire n_29211;
wire n_41700;
wire n_41687;
wire n_21281;
wire newNet_2692;
wire n_14829;
wire n_6162;
wire n_44035;
wire n_24415;
wire FE_OCP_RBN2289_n_2314;
wire n_42453;
wire n_33955;
wire n_2302;
wire n_24268;
wire FE_OCPN914_n_7832;
wire n_27607;
wire n_6948;
wire n_17667;
wire n_28879;
wire n_548;
wire n_42401;
wire n_21013;
wire n_13446;
wire n_11748;
wire newNet_3519;
wire n_5842;
wire n_14008;
wire n_47023;
wire n_42762;
wire n_33099;
wire newNet_680;
wire n_29959;
wire n_43326;
wire n_31486;
wire n_21447;
wire n_6234;
wire n_24830;
wire n_18003;
wire n_27034;
wire n_31404;
wire n_2349;
wire n_25217;
wire n_28781;
wire n_5532;
wire n_8915;
wire n_7742;
wire newNet_1221;
wire FE_RN_1724_0;
wire n_19313;
wire n_30369;
wire n_28061;
wire n_40494;
wire newNet_1606;
wire n_43211;
wire n_24518;
wire n_15643;
wire n_41878;
wire n_12954;
wire n_45874;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_7_;
wire n_5957;
wire n_43199;
wire n_45203;
wire n_17275;
wire n_10359;
wire n_4292;
wire n_41055;
wire n_11240;
wire n_6914;
wire n_8735;
wire n_27277;
wire n_32563;
wire n_37116;
wire n_16507;
wire n_2150;
wire n_18535;
wire n_11840;
wire FE_OCP_RBN1149_n_27962;
wire n_9663;
wire n_20303;
wire n_21337;
wire n_29577;
wire n_4169;
wire newNet_427;
wire n_2565;
wire n_7045;
wire n_12563;
wire n_5770;
wire FE_RN_623_0;
wire n_5775;
wire n_28472;
wire n_7627;
wire n_4675;
wire n_16648;
wire n_29524;
wire FE_OCP_RBN2232_n_13141;
wire newNet_3747;
wire n_38740;
wire n_9105;
wire n_9518;
wire FE_OCP_RBN2729_n_4219;
wire n_32239;
wire FE_OCP_RBN2892_n_26152;
wire n_21618;
wire n_16510;
wire FE_RN_1105_0;
wire n_30945;
wire FE_RN_1028_0;
wire newNet_908;
wire newNet_968;
wire newNet_629;
wire n_22116;
wire n_42004;
wire n_13601;
wire n_17145;
wire n_2437;
wire newNet_2031;
wire n_43241;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_24_;
wire n_10751;
wire n_1187;
wire n_3106;
wire n_41777;
wire n_42615;
wire n_33637;
wire n_24870;
wire n_20355;
wire n_28799;
wire n_145;
wire n_39596;
wire n_7201;
wire newNet_1368;
wire n_5190;
wire n_4659;
wire FE_RN_888_0;
wire n_39759;
wire n_41570;
wire n_22867;
wire n_30619;
wire n_10030;
wire n_25229;
wire newNet_3229;
wire newNet_3663;
wire n_37243;
wire n_26966;
wire n_37813;
wire n_2331;
wire n_37082;
wire n_26036;
wire n_41017;
wire FE_RN_412_0;
wire n_5483;
wire n_136;
wire newNet_2008;
wire n_12539;
wire n_18793;
wire n_38325;
wire n_41694;
wire n_890;
wire n_4630;
wire n_40368;
wire newNet_3258;
wire n_25372;
wire n_15890;
wire n_27433;
wire FE_RN_342_0;
wire n_23708;
wire n_7455;
wire n_17553;
wire FE_RN_854_0;
wire n_35192;
wire n_22376;
wire n_27860;
wire n_12061;
wire n_43188;
wire FE_RN_1184_0;
wire n_21066;
wire n_37131;
wire FE_OCP_RBN2528_n_3421;
wire n_38794;
wire newNet_2739;
wire n_4979;
wire n_44867;
wire n_32732;
wire FE_RN_1814_0;
wire n_18745;
wire n_36055;
wire n_41844;
wire n_5867;
wire n_23890;
wire n_18487;
wire n_34059;
wire FE_RN_797_0;
wire n_7816;
wire newNet_1270;
wire n_37561;
wire n_43914;
wire n_18259;
wire n_22611;
wire n_17401;
wire n_21450;
wire n_5649;
wire n_40507;
wire n_23125;
wire n_31807;
wire n_3161;
wire n_16173;
wire n_41592;
wire n_8444;
wire n_43916;
wire n_27774;
wire n_21390;
wire n_45816;
wire n_10959;
wire n_45766;
wire FE_OCP_RBN1710_n_22150;
wire n_21545;
wire n_19892;
wire n_3454;
wire n_38073;
wire n_32587;
wire n_686;
wire n_36132;
wire n_16440;
wire n_37349;
wire FE_OCP_DRV_N3149_n_12773;
wire n_40447;
wire delay_add_ln22_unr2_stage2_stallmux_q_17_;
wire n_5424;
wire n_33564;
wire newNet_2210;
wire newNet_2689;
wire n_43354;
wire n_35911;
wire n_24321;
wire FE_OCPN1520_n_31403;
wire n_23481;
wire n_34936;
wire n_25506;
wire n_1366;
wire n_6201;
wire n_6228;
wire n_32425;
wire n_35899;
wire n_42722;
wire n_3543;
wire n_38853;
wire n_42920;
wire n_30153;
wire n_38004;
wire n_2467;
wire n_26188;
wire n_27923;
wire n_17706;
wire n_32935;
wire n_22603;
wire newNet_2162;
wire n_23526;
wire n_7756;
wire n_6883;
wire n_19150;
wire n_40556;
wire n_10136;
wire n_31298;
wire n_36472;
wire n_39747;
wire n_22794;
wire n_31343;
wire n_705;
wire n_39248;
wire n_2516;
wire n_5591;
wire n_27390;
wire n_2639;
wire n_13251;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_23_;
wire newNet_2345;
wire n_8164;
wire n_30478;
wire n_12107;
wire n_23491;
wire n_29881;
wire newNet_1429;
wire n_17773;
wire n_29814;
wire n_11076;
wire n_12387;
wire n_23966;
wire n_21962;
wire n_7661;
wire n_37772;
wire n_46376;
wire n_39611;
wire n_19460;
wire n_36462;
wire n_2179;
wire n_5488;
wire n_17565;
wire newNet_266;
wire n_44592;
wire n_30183;
wire newNet_980;
wire newNet_552;
wire n_20716;
wire n_5432;
wire n_19407;
wire n_26334;
wire n_22468;
wire n_23515;
wire n_43804;
wire newNet_1506;
wire n_31208;
wire n_25684;
wire n_11379;
wire n_3471;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_20_;
wire n_43777;
wire n_30230;
wire n_42135;
wire n_32192;
wire n_9754;
wire n_12220;
wire n_21970;
wire n_3285;
wire n_40636;
wire n_32181;
wire FE_OCPN3178_n_21901;
wire n_1588;
wire n_29262;
wire n_10183;
wire n_21355;
wire n_18017;
wire n_29551;
wire n_18058;
wire delay_add_ln22_unr17_stage7_stallmux_q_18_;
wire n_2791;
wire n_22208;
wire n_32654;
wire n_5967;
wire n_8876;
wire n_42828;
wire n_19693;
wire n_28815;
wire n_34818;
wire n_32271;
wire newNet_2354;
wire newNet_1581;
wire n_37572;
wire FE_RN_800_0;
wire n_16953;
wire n_7670;
wire n_7978;
wire n_35861;
wire newNet_1125;
wire newNet_809;
wire n_45630;
wire n_3023;
wire n_26372;
wire n_11230;
wire n_38978;
wire FE_RN_277_0;
wire n_21869;
wire n_25350;
wire newNet_1403;
wire n_2576;
wire newNet_1427;
wire n_17453;
wire n_30531;
wire n_22108;
wire delay_xor_ln22_unr15_stage6_stallmux_q_11_;
wire newNet_2973;
wire n_13344;
wire n_1704;
wire n_17966;
wire n_16598;
wire n_27526;
wire FE_OCP_RBN1103_n_45224;
wire n_40487;
wire FE_OCP_RBN2909_n_26173;
wire newNet_2583;
wire FE_RN_236_0;
wire delay_add_ln22_unr2_stage2_stallmux_q_15_;
wire n_17467;
wire newNet_3200;
wire FE_RN_1819_0;
wire FE_OCP_RBN1363_n_20412;
wire newNet_1814;
wire n_29464;
wire n_40936;
wire n_36368;
wire n_9328;
wire n_32592;
wire FE_RN_891_0;
wire n_13747;
wire n_45633;
wire n_4970;
wire n_42467;
wire n_3871;
wire n_6397;
wire n_21042;
wire n_28304;
wire n_17360;
wire newNet_2292;
wire n_4397;
wire n_41142;
wire FE_OCP_RBN2496_n_8641;
wire n_18415;
wire n_34387;
wire n_41098;
wire n_12766;
wire n_33761;
wire n_33881;
wire n_14763;
wire n_40510;
wire n_17678;
wire n_11868;
wire n_19932;
wire n_21271;
wire n_23319;
wire n_31031;
wire n_5990;
wire n_27994;
wire n_6041;
wire n_10660;
wire n_23384;
wire n_25932;
wire n_17014;
wire n_32695;
wire n_4664;
wire n_24944;
wire n_36086;
wire beta_24;
wire n_9509;
wire n_39253;
wire n_29545;
wire FE_OCPN1793_n_30612;
wire delay_add_ln22_unr8_stage4_stallmux_q_3_;
wire newNet_1791;
wire beta_13;
wire n_33271;
wire n_31558;
wire n_36330;
wire n_17422;
wire delay_xor_ln22_unr15_stage6_stallmux_q_16_;
wire n_8476;
wire n_20547;
wire n_22497;
wire n_35856;
wire FE_RN_819_0;
wire newNet_3052;
wire FE_OCP_RBN3093_n_11475;
wire n_38873;
wire FE_RN_1682_0;
wire newNet_651;
wire newNet_3466;
wire cos_out_1;
wire n_36264;
wire n_12670;
wire n_43103;
wire n_1462;
wire n_26111;
wire FE_OCP_DRV_N1570_n_29777;
wire n_32769;
wire newNet_2319;
wire n_16978;
wire n_23312;
wire n_28267;
wire n_34366;
wire n_28506;
wire newNet_3643;
wire n_24264;
wire n_32007;
wire n_6038;
wire n_36627;
wire FE_OFN807_n_46195;
wire n_16056;
wire n_7272;
wire FE_OCP_RBN2458_n_13765;
wire n_12024;
wire n_8107;
wire FE_RN_303_0;
wire n_27425;
wire n_6594;
wire FE_OCPN912_n_43022;
wire n_40930;
wire n_35815;
wire n_26684;
wire n_12937;
wire n_43087;
wire n_10678;
wire n_25068;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_30_;
wire n_40371;
wire n_26142;
wire n_40036;
wire n_42619;
wire n_8862;
wire n_14476;
wire n_17623;
wire n_21664;
wire n_38108;
wire n_37713;
wire n_29190;
wire newNet_3067;
wire n_15382;
wire n_8653;
wire n_42364;
wire n_34835;
wire newNet_2012;
wire n_38626;
wire n_13536;
wire newNet_2671;
wire n_12824;
wire n_15225;
wire FE_OCP_RBN1362_n_20504;
wire n_47024;
wire newNet_150;
wire n_18142;
wire n_41541;
wire n_40689;
wire n_28627;
wire FE_OCPN976_n_31594;
wire n_1201;
wire n_28161;
wire n_31316;
wire n_40397;
wire n_18843;
wire n_28427;
wire newNet_1602;
wire n_30447;
wire n_43836;
wire n_32881;
wire n_11558;
wire FE_OCP_RBN3423_n_37794;
wire newNet_1885;
wire n_42312;
wire n_4891;
wire n_141;
wire n_39464;
wire n_31456;
wire n_32610;
wire n_43619;
wire n_361;
wire n_39677;
wire n_26954;
wire n_27848;
wire n_40121;
wire n_41654;
wire n_21147;
wire n_30914;
wire n_38000;
wire n_10070;
wire newNet_51;
wire n_5228;
wire n_30687;
wire n_29792;
wire n_34662;
wire n_11777;
wire n_10027;
wire FE_OCPN857_n_45697;
wire n_27151;
wire n_34622;
wire n_34119;
wire newNet_3252;
wire n_6390;
wire n_37333;
wire n_10004;
wire n_31796;
wire n_32971;
wire n_27695;
wire n_644;
wire n_31338;
wire FE_RN_1823_0;
wire newNet_1474;
wire n_30202;
wire n_41263;
wire n_12961;
wire n_18311;
wire FE_OCPN899_n_44593;
wire FE_RN_593_0;
wire n_36834;
wire n_40810;
wire FE_RN_1112_0;
wire n_21756;
wire n_22936;
wire n_10729;
wire n_21362;
wire n_40188;
wire n_41705;
wire n_36242;
wire n_8975;
wire n_30393;
wire n_7986;
wire n_18572;
wire n_36099;
wire newNet_137;
wire n_4118;
wire n_14213;
wire n_42610;
wire n_12846;
wire n_2932;
wire n_11458;
wire n_29365;
wire n_35625;
wire n_38737;
wire n_24520;
wire n_35674;
wire n_24469;
wire n_35981;
wire n_12944;
wire n_31336;
wire n_19742;
wire n_35381;
wire n_22637;
wire n_14498;
wire n_33526;
wire n_9413;
wire n_17671;
wire n_23450;
wire n_14917;
wire n_25053;
wire n_10332;
wire n_35939;
wire n_23388;
wire n_41327;
wire n_18113;
wire n_18726;
wire n_7761;
wire n_40458;
wire n_13005;
wire n_1507;
wire n_35018;
wire n_2608;
wire n_18761;
wire newNet_197;
wire newNet_959;
wire n_31222;
wire n_3751;
wire n_6316;
wire n_4524;
wire n_14815;
wire newNet_592;
wire n_12508;
wire n_23486;
wire n_34039;
wire n_20639;
wire n_27074;
wire n_38321;
wire n_39046;
wire n_19390;
wire n_11479;
wire n_37809;
wire n_32494;
wire n_35992;
wire n_34499;
wire n_25285;
wire n_32717;
wire n_27427;
wire n_27666;
wire FE_OCP_RBN2375_n_8221;
wire n_32447;
wire n_15661;
wire FE_OCPN1769_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire n_30143;
wire n_43564;
wire n_33251;
wire n_4900;
wire n_42161;
wire n_16620;
wire n_37749;
wire n_43018;
wire n_28334;
wire n_31256;
wire n_28146;
wire FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_12616;
wire n_31825;
wire n_17990;
wire n_13551;
wire n_19859;
wire n_4956;
wire n_21945;
wire newNet_1257;
wire n_30612;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_29_;
wire newNet_1990;
wire n_4271;
wire n_28741;
wire newNet_3384;
wire n_3508;
wire n_24394;
wire n_31105;
wire n_4717;
wire n_39912;
wire n_43614;
wire FE_RN_387_0;
wire n_30839;
wire n_43549;
wire n_21262;
wire FE_OCPN1795_n_30546;
wire n_29373;
wire n_24503;
wire n_12928;
wire n_42586;
wire n_30370;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_11_;
wire n_33293;
wire n_33686;
wire n_16824;
wire n_25340;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_17_;
wire FE_RN_972_0;
wire n_26587;
wire n_29633;
wire n_2731;
wire n_41521;
wire newNet_354;
wire n_13673;
wire n_26238;
wire n_27762;
wire FE_OCPN1513_FE_OFN738_n_22641;
wire n_15302;
wire n_25801;
wire newNet_506;
wire n_45528;
wire newNet_2410;
wire n_3510;
wire cos_out_28;
wire newNet_2336;
wire n_29871;
wire n_29843;
wire n_23445;
wire n_5661;
wire FE_RN_1729_0;
wire n_10884;
wire n_23819;
wire n_19590;
wire n_2549;
wire n_37006;
wire n_37634;
wire n_460;
wire n_36677;
wire n_7844;
wire n_18937;
wire FE_RN_1111_0;
wire n_15092;
wire n_39265;
wire newNet_399;
wire n_36600;
wire FE_OCPN970_n_14716;
wire n_40687;
wire n_35524;
wire FE_OCP_RBN1911_n_20545;
wire n_41308;
wire newNet_2341;
wire n_44060;
wire n_1155;
wire n_25206;
wire n_5547;
wire n_342;
wire n_17996;
wire n_12819;
wire newNet_3361;
wire n_3963;
wire FE_OCP_RBN1373_n_35275;
wire newNet_1818;
wire n_40085;
wire newNet_570;
wire n_40336;
wire n_3807;
wire n_22763;
wire n_5299;
wire n_20724;
wire n_25402;
wire n_27489;
wire n_31526;
wire delay_add_ln22_unr2_stage2_stallmux_q_13_;
wire n_13636;
wire n_11543;
wire n_14495;
wire n_206;
wire newNet_2048;
wire n_46161;
wire n_21419;
wire n_28064;
wire newNet_3415;
wire n_2770;
wire n_3583;
wire n_11875;
wire n_39149;
wire n_28889;
wire n_30870;
wire n_43897;
wire n_43094;
wire n_14635;
wire n_31174;
wire n_26338;
wire FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_40473;
wire FE_RN_1073_0;
wire n_11170;
wire n_19353;
wire n_40608;
wire n_33007;
wire n_29788;
wire n_22346;
wire n_28281;
wire n_29810;
wire FE_RN_1253_0;
wire n_40943;
wire newNet_3493;
wire n_35613;
wire newNet_3418;
wire n_21278;
wire n_15738;
wire n_27353;
wire n_29601;
wire n_43138;
wire FE_RN_147_0;
wire n_5780;
wire n_28397;
wire n_36371;
wire n_30580;
wire n_16143;
wire n_6215;
wire n_34110;
wire n_31359;
wire n_282;
wire n_27662;
wire n_340;
wire newNet_305;
wire n_20017;
wire n_25783;
wire n_15458;
wire n_4428;
wire n_11266;
wire n_23495;
wire FE_RN_1727_0;
wire n_3361;
wire n_8781;
wire n_18418;
wire n_29150;
wire n_39882;
wire n_30177;
wire n_32188;
wire n_20464;
wire n_36011;
wire n_28593;
wire n_24671;
wire n_43121;
wire n_43501;
wire FE_RN_11_0;
wire n_28366;
wire n_698;
wire n_10304;
wire n_4606;
wire n_37764;
wire FE_RN_113_0;
wire n_32196;
wire FE_OCP_RBN1707_n_20616;
wire FE_OCP_DRV_N3153_n_24425;
wire n_32147;
wire FE_OCP_RBN3397_n_37624;
wire n_37474;
wire n_11356;
wire n_1025;
wire n_6560;
wire n_43117;
wire newNet_850;
wire n_35154;
wire n_11959;
wire delay_sub_ln23_0_unr1_stage2_stallmux_q_0_;
wire n_33243;
wire n_819;
wire n_33345;
wire n_20055;
wire n_7746;
wire n_22808;
wire n_34866;
wire n_19281;
wire n_40024;
wire n_43599;
wire n_12431;
wire newNet_2405;
wire n_35792;
wire FE_RN_1210_0;
wire n_8017;
wire n_23921;
wire n_11196;
wire n_20153;
wire n_9335;
wire n_16269;
wire n_23938;
wire n_42284;
wire n_488;
wire n_9580;
wire n_6764;
wire n_2818;
wire n_24096;
wire n_15912;
wire n_38307;
wire n_19763;
wire n_20540;
wire newNet_1056;
wire n_38648;
wire n_12108;
wire FE_OCP_RBN2965_n_26231;
wire n_38834;
wire n_14436;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_6_;
wire n_10878;
wire n_30318;
wire n_8550;
wire n_1530;
wire FE_RN_1348_0;
wire n_17719;
wire n_27964;
wire n_39805;
wire newNet_1800;
wire n_36879;
wire n_18150;
wire FE_RN_215_0;
wire n_33756;
wire n_14083;
wire n_18701;
wire n_13256;
wire n_4797;
wire n_26350;
wire FE_OCP_RBN2736_n_14985;
wire n_10495;
wire FE_RN_1207_0;
wire n_5412;
wire n_17106;
wire n_23236;
wire newNet_409;
wire n_7436;
wire n_25144;
wire n_30783;
wire n_25695;
wire n_21883;
wire n_4921;
wire n_28249;
wire n_5688;
wire n_29585;
wire newNet_2328;
wire n_15727;
wire n_35375;
wire FE_RN_896_0;
wire n_21833;
wire n_42635;
wire newNet_1453;
wire FE_OCP_RBN3710_n_46337;
wire n_30095;
wire n_11995;
wire n_15897;
wire n_28768;
wire newNet_496;
wire n_16207;
wire n_26716;
wire n_12189;
wire n_15493;
wire delay_add_ln22_unr14_stage6_stallmux_q_7_;
wire FE_OCP_RBN2475_n_8664;
wire n_11501;
wire n_7704;
wire n_13848;
wire n_38357;
wire n_27584;
wire n_20344;
wire n_37224;
wire n_32623;
wire n_3035;
wire n_34895;
wire newNet_1844;
wire n_27501;
wire n_11595;
wire newNet_1406;
wire FE_RN_1474_0;
wire n_32822;
wire n_30020;
wire n_17047;
wire n_1925;
wire n_43581;
wire n_42174;
wire n_43551;
wire n_8256;
wire n_39762;
wire n_43878;
wire n_38708;
wire n_27231;
wire n_42532;
wire n_26286;
wire n_25194;
wire n_29019;
wire n_40195;
wire newNet_32;
wire n_14120;
wire n_31109;
wire n_14344;
wire n_42103;
wire n_11734;
wire newNet_1157;
wire n_38255;
wire n_13813;
wire n_2559;
wire n_16223;
wire n_29121;
wire n_30620;
wire n_4338;
wire n_9561;
wire FE_OCP_RBN3457_n_33872;
wire n_8524;
wire n_22531;
wire FE_RN_135_0;
wire n_47235;
wire n_33959;
wire delay_xor_ln21_unr21_stage8_stallmux_q_4_;
wire n_5820;
wire n_29074;
wire n_37840;
wire n_22232;
wire n_39237;
wire n_2335;
wire n_30967;
wire n_1224;
wire n_22815;
wire n_1941;
wire n_18742;
wire n_6866;
wire newNet_2521;
wire n_25719;
wire n_9050;
wire n_43876;
wire n_39285;
wire n_7126;
wire n_14350;
wire n_28937;
wire n_3046;
wire n_16893;
wire n_14959;
wire n_28785;
wire n_6581;
wire n_501;
wire n_11270;
wire n_1189;
wire n_1821;
wire n_39945;
wire n_31684;
wire n_17194;
wire n_36906;
wire n_4622;
wire n_29451;
wire n_14361;
wire n_11072;
wire n_37088;
wire n_6524;
wire n_26975;
wire n_14549;
wire n_16444;
wire n_39977;
wire n_22299;
wire n_40531;
wire n_4045;
wire n_39972;
wire n_33833;
wire n_5363;
wire n_33404;
wire n_42596;
wire n_42182;
wire n_11059;
wire n_9593;
wire n_12445;
wire n_5194;
wire n_7392;
wire n_39413;
wire n_14679;
wire n_35368;
wire FE_RN_744_0;
wire n_33483;
wire n_4488;
wire n_27173;
wire n_18032;
wire n_3288;
wire FE_RN_565_0;
wire n_42664;
wire n_17663;
wire n_13790;
wire newNet_1279;
wire n_28711;
wire n_32366;
wire n_11221;
wire n_13858;
wire n_36306;
wire n_23155;
wire n_8110;
wire FE_OCP_RBN1703_n_19560;
wire n_20004;
wire n_43676;
wire n_35765;
wire n_26292;
wire n_32655;
wire n_22759;
wire delay_add_ln22_unr14_stage6_stallmux_q_24_;
wire newNet_224;
wire n_36366;
wire newNet_3267;
wire n_32557;
wire n_36215;
wire n_30120;
wire n_8299;
wire newNet_1820;
wire FE_OCP_RBN3558_n_8687;
wire n_42608;
wire n_21720;
wire FE_RN_1543_0;
wire n_33842;
wire n_2223;
wire n_12474;
wire n_17268;
wire n_35342;
wire n_26473;
wire n_19184;
wire n_31678;
wire FE_OCPN913_n_43022;
wire n_9791;
wire n_30324;
wire n_32345;
wire n_2154;
wire newNet_175;
wire n_12200;
wire n_7009;
wire delay_add_ln22_unr11_stage5_stallmux_q_18_;
wire newNet_3095;
wire n_7825;
wire n_467;
wire n_28127;
wire n_32663;
wire n_3680;
wire n_7289;
wire n_11589;
wire n_5289;
wire n_39418;
wire n_32304;
wire n_1138;
wire n_11197;
wire n_35545;
wire n_28829;
wire FE_OCP_RBN3549_n_44575;
wire n_35751;
wire n_15615;
wire newNet_130;
wire n_5012;
wire n_42124;
wire n_22197;
wire n_38836;
wire FE_OCP_RBN2439_n_8402;
wire n_24363;
wire newNet_117;
wire n_33513;
wire n_25834;
wire n_13409;
wire n_23798;
wire n_37433;
wire delay_add_ln22_unr2_stage2_stallmux_q_28_;
wire n_45139;
wire n_541;
wire n_37085;
wire n_12323;
wire n_5614;
wire n_28774;
wire n_37485;
wire n_451;
wire n_8899;
wire newNet_3302;
wire n_39184;
wire n_749;
wire n_29268;
wire newNet_124;
wire FE_OCPN952_n_41540;
wire n_4307;
wire n_30501;
wire n_2807;
wire newNet_730;
wire n_28297;
wire n_35779;
wire n_3761;
wire n_1453;
wire n_24113;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_4_;
wire newNet_3483;
wire n_42155;
wire n_25071;
wire newNet_1397;
wire n_6090;
wire n_25775;
wire n_6897;
wire n_18102;
wire n_37554;
wire n_30865;
wire n_36226;
wire n_43453;
wire n_28867;
wire n_15979;
wire n_16721;
wire n_37836;
wire n_38988;
wire n_17849;
wire n_18475;
wire n_7441;
wire n_30496;
wire n_36499;
wire n_17921;
wire n_5944;
wire newNet_1340;
wire n_41605;
wire n_40204;
wire n_11297;
wire n_13758;
wire n_12033;
wire n_1082;
wire n_46382;
wire n_10921;
wire n_21420;
wire n_14034;
wire n_20843;
wire n_32878;
wire newNet_891;
wire n_1729;
wire n_20256;
wire n_11408;
wire n_46357;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_20_;
wire n_9205;
wire n_23775;
wire n_21941;
wire n_17945;
wire n_23069;
wire n_13789;
wire n_25803;
wire newNet_449;
wire n_1895;
wire n_1635;
wire n_6981;
wire n_20932;
wire FE_OCP_RBN2797_n_10106;
wire n_17003;
wire newNet_464;
wire n_10061;
wire n_36064;
wire FE_OCP_RBN3374_n_6745;
wire n_37731;
wire n_7497;
wire n_39874;
wire FE_OCP_RBN1163_n_13726;
wire n_34302;
wire n_20147;
wire n_32414;
wire n_35032;
wire n_43227;
wire n_3946;
wire FE_OFN828_n_29140;
wire n_17906;
wire n_39771;
wire n_21381;
wire n_24339;
wire newNet_317;
wire n_23172;
wire n_42142;
wire n_19430;
wire n_39577;
wire n_4050;
wire FE_RN_831_0;
wire newNet_877;
wire n_7302;
wire n_7520;
wire n_43172;
wire n_2433;
wire n_32076;
wire n_32214;
wire n_17799;
wire n_32473;
wire n_39234;
wire delay_add_ln22_unr11_stage5_stallmux_q_25_;
wire n_17040;
wire n_12865;
wire n_14885;
wire n_9879;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_12_;
wire n_6993;
wire n_32223;
wire n_15634;
wire n_41228;
wire FE_OCP_RBN2790_n_4462;
wire n_28645;
wire n_44039;
wire n_40137;
wire n_21847;
wire FE_OCP_RBN3403_n_28597;
wire newNet_432;
wire n_26121;
wire n_35101;
wire FE_OCPN1509_n_44174;
wire n_7716;
wire n_32351;
wire FE_RN_1609_0;
wire n_4862;
wire n_7569;
wire n_15208;
wire FE_OCPN1453_n_18559;
wire n_27902;
wire n_34670;
wire n_34796;
wire n_40146;
wire FE_OCPN3179_FE_OCP_RBN2744_n_15319;
wire n_30995;
wire newNet_2596;
wire n_37976;
wire n_6754;
wire n_39709;
wire delay_add_ln22_unr27_stage10_stallmux_q_20_;
wire n_17543;
wire n_29738;
wire n_41907;
wire n_23107;
wire n_18630;
wire n_33571;
wire newNet_2514;
wire FE_RN_1830_0;
wire n_4543;
wire n_6873;
wire n_11636;
wire n_7638;
wire n_34531;
wire FE_OCP_RBN1170_n_13756;
wire n_2218;
wire n_43027;
wire n_18677;
wire n_38094;
wire n_30388;
wire n_2662;
wire newNet_872;
wire n_1550;
wire n_7852;
wire n_25503;
wire n_22771;
wire n_17458;
wire n_16410;
wire n_5520;
wire n_3977;
wire newNet_2071;
wire n_16265;
wire newNet_1320;
wire n_26386;
wire n_24422;
wire n_6457;
wire n_18208;
wire n_27023;
wire newNet_2772;
wire n_23283;
wire n_9760;
wire n_17474;
wire n_26414;
wire n_42621;
wire n_32254;
wire newNet_597;
wire n_19503;
wire n_24150;
wire n_3573;
wire n_6335;
wire n_29329;
wire n_36283;
wire n_7112;
wire n_17235;
wire n_37362;
wire n_37887;
wire n_17516;
wire n_6345;
wire FE_RN_816_0;
wire n_3742;
wire FE_RN_1640_0;
wire n_10889;
wire newNet_2763;
wire n_4393;
wire n_43867;
wire FE_OCP_RBN1674_n_36492;
wire n_26978;
wire FE_OCPN903_n_44581;
wire n_13338;
wire n_18803;
wire n_11714;
wire newNet_2180;
wire newNet_2105;
wire FE_RN_478_0;
wire n_40174;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_30_;
wire n_21004;
wire n_41204;
wire n_15684;
wire n_37052;
wire n_23342;
wire n_8154;
wire n_10813;
wire n_5724;
wire n_33445;
wire n_39338;
wire n_5397;
wire delay_add_ln22_unr17_stage7_stallmux_q_1_;
wire n_5188;
wire n_25845;
wire n_40461;
wire n_7580;
wire n_13160;
wire n_39366;
wire FE_OCP_RBN3638_n_44490;
wire FE_OCPN990_n_22249;
wire n_37758;
wire n_14279;
wire n_13200;
wire n_16669;
wire newNet_2846;
wire n_41589;
wire n_11177;
wire n_34728;
wire n_10665;
wire n_29644;
wire n_4346;
wire n_29657;
wire n_16814;
wire n_9393;
wire n_37169;
wire n_31029;
wire n_5305;
wire n_24564;
wire n_34846;
wire n_24085;
wire n_2798;
wire FE_OFN792_n_25938;
wire n_8203;
wire newNet_2961;
wire newNet_1386;
wire n_3206;
wire n_16554;
wire newNet_1347;
wire FE_OCP_RBN3132_n_27736;
wire n_21482;
wire n_40826;
wire FE_OCPN895_n_6521;
wire n_12135;
wire n_45180;
wire n_19961;
wire n_37852;
wire n_34459;
wire n_5997;
wire n_110;
wire n_5172;
wire n_36196;
wire n_4987;
wire n_7093;
wire n_31904;
wire n_5753;
wire sin_out_9;
wire n_29488;
wire n_5087;
wire n_35075;
wire n_25951;
wire n_17333;
wire newNet_1198;
wire FE_OCP_RBN2219_n_12698;
wire n_5261;
wire n_30078;
wire n_20855;
wire newNet_2788;
wire n_1705;
wire n_277;
wire n_17031;
wire newNet_2803;
wire n_27213;
wire n_8574;
wire newNet_2985;
wire newNet_366;
wire n_32842;
wire n_25516;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_1_;
wire n_30744;
wire newNet_2120;
wire n_32283;
wire n_3431;
wire n_42485;
wire n_38739;
wire n_15238;
wire n_2126;
wire n_36271;
wire n_42353;
wire n_11938;
wire n_1512;
wire n_5387;
wire n_9088;
wire n_38693;
wire n_11083;
wire n_13713;
wire n_42040;
wire FE_RN_384_0;
wire FE_RN_1072_0;
wire n_14701;
wire n_1237;
wire n_41517;
wire FE_OCP_RBN2471_n_34285;
wire n_8295;
wire n_677;
wire n_39505;
wire newNet_2758;
wire n_24534;
wire n_33307;
wire n_10243;
wire n_3281;
wire FE_OCP_RBN2478_n_8599;
wire n_43727;
wire n_11238;
wire n_33629;
wire n_37586;
wire n_15778;
wire n_20852;
wire newNet_1185;
wire n_23540;
wire FE_RN_1587_0;
wire newNet_238;
wire delay_xor_ln21_unr9_stage4_stallmux_q_11_;
wire newNet_3076;
wire n_21021;
wire n_27709;
wire newNet_1025;
wire n_10744;
wire newNet_1681;
wire n_13768;
wire n_3853;
wire n_20329;
wire n_27686;
wire newNet_380;
wire n_23591;
wire newNet_2912;
wire n_24590;
wire newNet_3488;
wire n_43858;
wire n_7321;
wire n_26828;
wire n_34716;
wire n_22845;
wire n_40908;
wire n_24145;
wire n_36154;
wire n_16822;
wire n_40912;
wire n_3715;
wire FE_OCP_RBN2919_n_16084;
wire n_21195;
wire n_34396;
wire n_35584;
wire n_12383;
wire n_18214;
wire newNet_2322;
wire n_25637;
wire n_37876;
wire n_12248;
wire n_7659;
wire n_26399;
wire n_15343;
wire n_23979;
wire n_32772;
wire n_18482;
wire n_10704;
wire n_15961;
wire n_38396;
wire n_2489;
wire n_22618;
wire n_41832;
wire n_31283;
wire n_30594;
wire n_29773;
wire n_18522;
wire n_23909;
wire n_25256;
wire n_11765;
wire n_14859;
wire n_6196;
wire FE_OCP_DRV_N1585_n_35594;
wire n_4352;
wire n_35235;
wire FE_OCPN1433_n_30614;
wire n_26382;
wire n_21910;
wire newNet_1036;
wire n_43577;
wire n_14147;
wire n_2172;
wire n_15116;
wire n_10951;
wire n_4837;
wire n_9401;
wire FE_OCP_RBN2696_n_14814;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_2_;
wire n_38971;
wire n_37160;
wire newNet_3211;
wire n_9482;
wire n_29606;
wire n_21785;
wire n_29516;
wire n_1420;
wire n_14972;
wire n_40390;
wire n_1498;
wire n_26888;
wire FE_OCPN966_n_47020;
wire n_25427;
wire n_15333;
wire n_8607;
wire n_42862;
wire n_1317;
wire FE_RN_665_0;
wire FE_OCP_RBN3417_n_12739;
wire n_16616;
wire n_16316;
wire n_1955;
wire n_40509;
wire n_7028;
wire n_18189;
wire n_24763;
wire newNet_1742;
wire FE_OCP_RBN3057_n_36506;
wire newNet_3732;
wire n_1910;
wire n_21692;
wire FE_OCP_RBN2768_n_9745;
wire n_16792;
wire n_42027;
wire n_7622;
wire FE_OCP_DRV_N1551_n_19010;
wire newNet_2601;
wire n_1624;
wire n_42030;
wire n_38601;
wire n_34533;
wire FE_OCP_DRV_N1566_n_28654;
wire n_19404;
wire newNet_2722;
wire n_41239;
wire n_17839;
wire n_43257;
wire n_7286;
wire n_15206;
wire n_6076;
wire n_6671;
wire n_9283;
wire n_32264;
wire n_24694;
wire n_26848;
wire n_34375;
wire newNet_419;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_5_;
wire n_6789;
wire n_7511;
wire n_29998;
wire n_42372;
wire n_9629;
wire n_18159;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_15_;
wire n_16872;
wire n_16353;
wire FE_OFN829_n_2405;
wire n_10801;
wire n_34184;
wire n_27132;
wire FE_RN_860_0;
wire newNet_2639;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_3_;
wire n_11806;
wire n_24438;
wire n_10197;
wire n_41122;
wire newNet_1628;
wire n_12871;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_8_;
wire FE_OCP_RBN2967_n_26580;
wire n_40876;
wire n_19474;
wire n_21076;
wire FE_OCP_RBN2818_n_4458;
wire newNet_3329;
wire n_34297;
wire n_27771;
wire n_24481;
wire n_34157;
wire n_38858;
wire n_31293;
wire n_13451;
wire n_957;
wire n_14107;
wire n_41081;
wire n_18055;
wire n_10389;
wire newNet_617;
wire n_34800;
wire n_34900;
wire n_1657;
wire n_42498;
wire n_32925;
wire n_31239;
wire n_34692;
wire n_29101;
wire newNet_2567;
wire newNet_1093;
wire n_5911;
wire newNet_2664;
wire n_23264;
wire n_10850;
wire n_33415;
wire delay_add_ln22_unr23_stage9_stallmux_q_19_;
wire n_6798;
wire FE_RN_1309_0;
wire delay_xor_ln21_unr18_stage7_stallmux_q_2_;
wire n_36702;
wire FE_RN_822_0;
wire n_1052;
wire n_11673;
wire n_2463;
wire n_229;
wire n_4817;
wire newNet_3377;
wire n_5469;
wire n_13395;
wire n_42511;
wire n_25925;
wire n_15795;
wire n_33151;
wire newNet_1785;
wire n_25128;
wire n_23356;
wire n_30039;
wire n_32224;
wire n_36587;
wire FE_OCP_RBN3589_n_47014;
wire n_9837;
wire n_3115;
wire newNet_1614;
wire FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire n_18546;
wire n_29713;
wire FE_RN_1610_0;
wire n_2111;
wire newNet_2366;
wire n_30633;
wire n_8646;
wire n_9322;
wire FE_RN_40_0;
wire n_29558;
wire FE_RN_982_0;
wire n_16573;
wire newNet_3264;
wire newNet_2029;
wire n_2475;
wire n_4092;
wire n_9363;
wire n_4565;
wire n_2310;
wire n_17959;
wire n_24111;
wire n_38757;
wire n_40440;
wire n_27733;
wire n_31987;
wire n_24491;
wire n_33992;
wire n_11042;
wire FE_OCP_RBN3736_n_27535;
wire n_47015;
wire n_42111;
wire newNet_1415;
wire n_14714;
wire newNet_3755;
wire newNet_3191;
wire FE_OCPN852_n_694;
wire newNet_511;
wire n_26751;
wire n_15413;
wire n_31645;
wire n_34094;
wire n_9757;
wire n_37186;
wire n_37313;
wire n_5458;
wire n_26781;
wire n_10777;
wire n_38423;
wire FE_OCPN3765_FE_OCP_RBN2222_n_13010;
wire n_18243;
wire delay_xor_ln22_unr9_stage4_stallmux_q_15_;
wire FE_OCP_RBN2595_n_25181;
wire n_43266;
wire n_31046;
wire n_38610;
wire n_25414;
wire n_31758;
wire FE_OCP_RBN3517_n_8498;
wire n_5601;
wire n_9891;
wire n_43239;
wire FE_RN_476_0;
wire n_26703;
wire n_33865;
wire n_22461;
wire n_8066;
wire n_21715;
wire n_17805;
wire n_24975;
wire n_25759;
wire FE_RN_1639_0;
wire n_22169;
wire n_79;
wire n_46979;
wire FE_OCP_RBN2677_n_9247;
wire n_29008;
wire n_33545;
wire n_1758;
wire n_3072;
wire n_17911;
wire n_25654;
wire FE_RN_1281_0;
wire n_32450;
wire n_38844;
wire n_26167;
wire n_1164;
wire newNet_2473;
wire n_21187;
wire n_33940;
wire n_3872;
wire n_21028;
wire n_19064;
wire n_43525;
wire n_4298;
wire n_12418;
wire n_28244;
wire newNet_1304;
wire n_18518;
wire n_26034;
wire n_35567;
wire n_40004;
wire newNet_3741;
wire n_9219;
wire n_37340;
wire n_21050;
wire n_5778;
wire n_12376;
wire n_23537;
wire n_30489;
wire n_41841;
wire n_12205;
wire n_1822;
wire FE_OCP_RBN2261_n_33691;
wire n_1363;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_10_;
wire n_40433;
wire n_4185;
wire n_26564;
wire n_22462;
wire n_31191;
wire n_11945;
wire n_30507;
wire FE_RN_1123_0;
wire newNet_1302;
wire n_43329;
wire n_30171;
wire n_11015;
wire n_16126;
wire n_4679;
wire n_17558;
wire FE_RN_1655_0;
wire n_11035;
wire n_17394;
wire n_28125;
wire FE_RN_909_0;
wire n_14743;
wire n_114;
wire n_35505;
wire n_6641;
wire n_13613;
wire n_32799;
wire FE_OCP_RBN2714_n_14982;
wire n_6165;
wire n_41095;
wire n_26331;
wire newNet_1178;
wire n_7190;
wire n_11655;
wire n_16373;
wire n_23870;
wire n_37601;
wire n_36389;
wire n_45462;
wire n_68;
wire n_37382;
wire n_17946;
wire n_4147;
wire FE_RN_499_0;
wire newNet_1162;
wire n_2155;
wire n_38188;
wire FE_RN_922_0;
wire n_33910;
wire n_14441;
wire n_7608;
wire n_22042;
wire n_41244;
wire n_1731;
wire n_24645;
wire newNet_1648;
wire n_10756;
wire newNet_1339;
wire n_25196;
wire n_32314;
wire n_11239;
wire n_28441;
wire n_38847;
wire FE_OCP_RBN2349_n_38515;
wire newNet_2213;
wire delay_add_ln22_unr2_stage2_stallmux_q_31_;
wire n_14003;
wire n_1856;
wire n_42775;
wire n_43728;
wire n_33930;
wire n_32121;
wire n_24651;
wire n_37023;
wire n_6791;
wire n_17459;
wire n_9781;
wire n_31483;
wire n_29886;
wire FE_OCPN1401_n_9642;
wire n_2582;
wire n_41567;
wire n_7402;
wire n_15711;
wire n_24051;
wire n_41256;
wire n_14628;
wire FE_RN_1495_0;
wire n_31340;
wire n_35357;
wire n_4394;
wire delay_xor_ln21_unr15_stage6_stallmux_q_5_;
wire n_24288;
wire newNet_3300;
wire newNet_1350;
wire n_40119;
wire n_33665;
wire n_14207;
wire n_4672;
wire FE_OCPN3795_FE_RN_1789_0;
wire n_7507;
wire n_42529;
wire n_24591;
wire n_2338;
wire FE_RN_1176_0;
wire newNet_1622;
wire n_32861;
wire FE_OCP_RBN2236_n_29055;
wire n_21442;
wire n_11795;
wire n_16576;
wire FE_OCP_RBN3707_n_16649;
wire n_3552;
wire n_7635;
wire n_28445;
wire n_37831;
wire newNet_390;
wire n_33968;
wire newNet_1487;
wire n_5055;
wire n_16511;
wire n_21793;
wire n_31647;
wire FE_OCPN1439_n_23339;
wire n_27523;
wire FE_RN_1270_0;
wire n_40342;
wire n_1053;
wire n_40881;
wire newNet_1782;
wire delay_xor_ln22_unr3_stage2_stallmux_q_2_;
wire n_35987;
wire n_21784;
wire n_4973;
wire n_42409;
wire n_9307;
wire n_18127;
wire n_28101;
wire n_38088;
wire n_29617;
wire n_4228;
wire n_12781;
wire n_37260;
wire n_29711;
wire delay_add_ln22_unr23_stage9_stallmux_q_20_;
wire newNet_2046;
wire n_14736;
wire n_33108;
wire n_33312;
wire n_37393;
wire n_11873;
wire n_35831;
wire newNet_2665;
wire n_6818;
wire n_20999;
wire n_1320;
wire n_37577;
wire n_8765;
wire FE_OCP_RBN2556_n_44576;
wire FE_OCP_RBN2621_n_44561;
wire n_22569;
wire n_200;
wire n_5171;
wire n_9204;
wire newNet_1241;
wire n_2487;
wire n_10190;
wire n_10133;
wire n_37823;
wire n_6129;
wire n_7908;
wire n_32985;
wire FE_RN_908_0;
wire n_38975;
wire n_2571;
wire n_22380;
wire n_14745;
wire n_7063;
wire n_2663;
wire n_37566;
wire delay_xor_ln22_unr21_stage8_stallmux_q_10_;
wire n_21996;
wire n_18526;
wire newNet_1400;
wire n_35229;
wire n_33567;
wire newNet_669;
wire n_27990;
wire n_26140;
wire n_23593;
wire n_36052;
wire n_6198;
wire newNet_2783;
wire n_16504;
wire n_19881;
wire newNet_983;
wire newNet_424;
wire n_12228;
wire n_32690;
wire n_42799;
wire n_6674;
wire newNet_2488;
wire FE_OCP_RBN3468_n_7886;
wire n_29030;
wire FE_OCPN1392_n_7925;
wire n_39010;
wire n_2455;
wire n_32303;
wire n_29278;
wire n_44426;
wire FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire newNet_2657;
wire n_14254;
wire n_33764;
wire n_18004;
wire n_8139;
wire n_7920;
wire n_8019;
wire n_38588;
wire delay_add_ln22_unr20_stage8_stallmux_q_31_;
wire n_26690;
wire n_16868;
wire FE_OCP_RBN2940_n_26276;
wire FE_RN_413_0;
wire FE_RN_1416_0;
wire newNet_591;
wire n_26254;
wire n_36649;
wire n_651;
wire n_4175;
wire n_15543;
wire FE_OCP_RBN2266_n_2430;
wire n_12820;
wire n_35177;
wire n_1093;
wire n_16879;
wire n_8835;
wire n_37140;
wire n_42541;
wire FE_OCP_RBN2294_n_2438;
wire n_32930;
wire n_27296;
wire n_30544;
wire n_35598;
wire newNet_3555;
wire n_34897;
wire n_34167;
wire n_14878;
wire FE_OCP_RBN2275_n_24077;
wire n_32736;
wire n_25395;
wire n_11548;
wire n_22929;
wire n_19740;
wire n_28577;
wire n_25425;
wire n_29299;
wire n_20755;
wire n_6683;
wire n_34993;
wire n_35265;
wire newNet_834;
wire n_28240;
wire n_3567;
wire n_35320;
wire newNet_3583;
wire n_10129;
wire FE_OCP_RBN3628_n_38870;
wire n_14710;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_15_;
wire n_42894;
wire n_42964;
wire n_78;
wire n_37061;
wire n_26028;
wire n_11070;
wire n_27846;
wire n_21391;
wire mux_while_ln12_psv_q_4_;
wire n_14211;
wire n_30411;
wire n_23899;
wire n_35976;
wire n_44962;
wire n_34453;
wire FE_OCP_RBN2821_n_10023;
wire n_38677;
wire n_34493;
wire n_44026;
wire n_15018;
wire n_22932;
wire n_46176;
wire n_19910;
wire sin_out_16;
wire n_23946;
wire n_1741;
wire n_22378;
wire n_23936;
wire n_8664;
wire FE_OCP_RBN2513_n_8533;
wire n_3335;
wire n_25564;
wire n_21264;
wire cos_out_15;
wire n_45513;
wire n_30300;
wire n_8389;
wire delay_xor_ln22_unr28_stage10_stallmux_q_1_;
wire n_9538;
wire n_31287;
wire n_24718;
wire n_37917;
wire FE_RN_1538_0;
wire n_23253;
wire newNet_2441;
wire n_40462;
wire n_36095;
wire n_29794;
wire n_38071;
wire n_23248;
wire n_8398;
wire n_22270;
wire n_41894;
wire n_35639;
wire n_133;
wire n_21718;
wire n_11957;
wire n_3298;
wire n_45638;
wire n_14860;
wire n_21510;
wire n_36830;
wire n_907;
wire n_2525;
wire n_43797;
wire n_26440;
wire n_14416;
wire n_40832;
wire n_43002;
wire FE_OCP_DRV_N3161_n_21419;
wire n_19719;
wire n_10584;
wire n_3506;
wire n_19949;
wire n_20915;
wire FE_RN_503_0;
wire n_28677;
wire n_23178;
wire newNet_2051;
wire n_12196;
wire FE_OCP_RBN3445_n_37945;
wire n_1906;
wire n_33261;
wire n_8494;
wire n_34562;
wire n_37081;
wire n_3419;
wire n_35538;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_8_;
wire n_22606;
wire n_23765;
wire n_23395;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_19_;
wire n_41664;
wire n_292;
wire newNet_2602;
wire n_45846;
wire n_36721;
wire n_25926;
wire n_25722;
wire n_7714;
wire n_43811;
wire n_12302;
wire n_28332;
wire n_14170;
wire n_14296;
wire n_15663;
wire n_43224;
wire n_18006;
wire n_471;
wire n_31446;
wire n_10262;
wire n_9194;
wire n_11852;
wire n_11716;
wire n_15822;
wire n_27697;
wire n_29383;
wire n_36549;
wire newNet_3173;
wire FE_RN_415_0;
wire n_5798;
wire n_30265;
wire n_12651;
wire n_19360;
wire n_28726;
wire n_45314;
wire n_34946;
wire n_33192;
wire n_376;
wire FE_RN_322_0;
wire n_13346;
wire FE_OFN779_n_17093;
wire n_25126;
wire n_16558;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_6_;
wire n_41750;
wire n_9676;
wire n_35694;
wire n_39498;
wire n_8199;
wire n_11698;
wire n_32857;
wire newNet_2240;
wire newNet_2581;
wire newNet_1805;
wire newNet_1762;
wire n_20485;
wire n_33628;
wire n_2264;
wire newNet_1880;
wire n_36125;
wire newNet_1545;
wire n_24515;
wire n_41543;
wire n_143;
wire n_29453;
wire n_4906;
wire n_8246;
wire n_17370;
wire n_3325;
wire n_36183;
wire n_2108;
wire n_32708;
wire newNet_2746;
wire n_36783;
wire n_22811;
wire n_42450;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_19_;
wire newNet_2823;
wire n_41680;
wire newNet_3592;
wire n_2633;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_5_;
wire n_7428;
wire n_21417;
wire n_28418;
wire n_34437;
wire FE_RN_389_0;
wire newNet_2343;
wire delay_xor_ln21_unr9_stage4_stallmux_q_17_;
wire newNet_1016;
wire n_3560;
wire n_5085;
wire newNet_1679;
wire n_39719;
wire n_14129;
wire n_18841;
wire n_28669;
wire n_13151;
wire n_100;
wire FE_OCP_RBN2567_n_8904;
wire n_1840;
wire n_25850;
wire n_6063;
wire n_42209;
wire n_1891;
wire n_40358;
wire n_2305;
wire n_542;
wire FE_RN_1202_0;
wire newNet_890;
wire n_4467;
wire n_17154;
wire n_21205;
wire n_29139;
wire delay_xor_ln22_unr6_stage3_stallmux_q_17_;
wire n_35490;
wire n_41224;
wire n_15944;
wire n_40250;
wire n_8682;
wire n_6324;
wire n_24084;
wire n_7744;
wire n_38749;
wire FE_OCP_RBN3120_n_27655;
wire n_28812;
wire n_37034;
wire newNet_687;
wire n_23705;
wire n_988;
wire n_31213;
wire n_5624;
wire n_38567;
wire FE_RN_1854_0;
wire FE_RN_1274_0;
wire n_32128;
wire n_7678;
wire n_2432;
wire n_34813;
wire newNet_2530;
wire n_7348;
wire n_6231;
wire n_4208;
wire n_26949;
wire n_35682;
wire newNet_3641;
wire n_6267;
wire n_30822;
wire newNet_381;
wire n_27024;
wire n_25859;
wire n_22115;
wire n_7846;
wire n_33750;
wire FE_RN_1748_0;
wire FE_OCPN889_n_7802;
wire n_15959;
wire n_28612;
wire n_43920;
wire n_10950;
wire newNet_3474;
wire n_14814;
wire FE_RN_627_0;
wire n_18620;
wire n_27926;
wire newNet_3754;
wire n_39255;
wire newNet_3339;
wire n_34446;
wire n_25889;
wire n_10657;
wire n_226;
wire n_13936;
wire n_1258;
wire n_17081;
wire n_22588;
wire n_22624;
wire n_26456;
wire n_18828;
wire delay_xor_ln22_unr6_stage3_stallmux_q_5_;
wire n_40634;
wire newNet_3050;
wire newNet_161;
wire n_12031;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_2_;
wire newNet_2619;
wire n_5115;
wire newNet_1414;
wire n_17987;
wire FE_RN_638_0;
wire n_9513;
wire newNet_2839;
wire n_19754;
wire n_29069;
wire n_27093;
wire n_15405;
wire n_19983;
wire n_27791;
wire n_6150;
wire n_36032;
wire n_32784;
wire FE_RN_1182_0;
wire n_31888;
wire n_38429;
wire n_3697;
wire n_6628;
wire n_18481;
wire n_14760;
wire newNet_2595;
wire n_40669;
wire n_18070;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_24_;
wire FE_OCP_RBN3527_n_13765;
wire n_27013;
wire n_18872;
wire n_14181;
wire n_28498;
wire n_34331;
wire n_28870;
wire FE_OCP_RBN2223_n_12902;
wire n_8709;
wire n_4518;
wire n_25309;
wire n_33342;
wire n_36887;
wire n_16962;
wire n_26866;
wire n_10365;
wire n_20450;
wire FE_OCP_RBN1909_n_20545;
wire n_37697;
wire n_29967;
wire n_33272;
wire n_11296;
wire n_28892;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_25_;
wire n_17405;
wire n_41482;
wire newNet_1731;
wire n_20818;
wire n_35292;
wire n_23831;
wire n_33544;
wire n_20244;
wire n_26069;
wire n_38408;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_31_;
wire n_37056;
wire n_14600;
wire n_22529;
wire n_27821;
wire FE_OCP_RBN3084_n_31819;
wire n_23385;
wire delay_add_ln22_unr14_stage6_stallmux_q_22_;
wire n_29853;
wire n_29267;
wire n_4536;
wire n_11328;
wire n_41966;
wire FE_OCP_RBN2288_n_2268;
wire n_26157;
wire n_5023;
wire n_41080;
wire n_3655;
wire newNet_2504;
wire n_42143;
wire n_5491;
wire FE_OCP_RBN3476_n_7886;
wire n_15366;
wire n_21251;
wire n_19029;
wire n_28179;
wire newNet_2384;
wire n_10630;
wire n_42612;
wire n_10869;
wire n_4732;
wire FE_OCPN951_n_41540;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_15_;
wire FE_RN_1861_0;
wire n_42949;
wire n_761;
wire n_14580;
wire n_41917;
wire n_6416;
wire n_16670;
wire n_7787;
wire n_30386;
wire n_34340;
wire n_44422;
wire n_4263;
wire n_24416;
wire n_5947;
wire n_41595;
wire n_36516;
wire n_32566;
wire n_29192;
wire n_24681;
wire n_4873;
wire FE_OCP_RBN3553_n_44575;
wire n_36750;
wire n_26761;
wire n_25847;
wire n_13867;
wire n_36327;
wire n_19989;
wire n_32102;
wire n_27610;
wire newNet_3685;
wire n_19920;
wire n_20348;
wire n_18221;
wire n_29647;
wire n_32973;
wire newNet_1208;
wire FE_RN_790_0;
wire n_37242;
wire n_40672;
wire newNet_920;
wire n_32272;
wire n_4742;
wire delay_add_ln22_unr5_stage3_stallmux_q_7_;
wire n_12732;
wire delay_xor_ln22_unr21_stage8_stallmux_q_6_;
wire n_1911;
wire n_24325;
wire n_15067;
wire n_4756;
wire n_31528;
wire n_34480;
wire n_8072;
wire n_6546;
wire n_32334;
wire n_32983;
wire n_29306;
wire n_2705;
wire n_3776;
wire n_28097;
wire n_35634;
wire n_11985;
wire n_13730;
wire n_4237;
wire n_41237;
wire n_1682;
wire n_42671;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_22_;
wire n_2294;
wire delay_xor_ln21_unr18_stage7_stallmux_q_3_;
wire n_37980;
wire n_13063;
wire n_9637;
wire n_17738;
wire n_21367;
wire n_3411;
wire newNet_3210;
wire n_9426;
wire n_43293;
wire n_41307;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_15_;
wire n_9922;
wire n_12100;
wire n_21626;
wire n_22156;
wire n_12576;
wire n_25132;
wire FE_OCP_RBN2396_n_24451;
wire n_29766;
wire n_2732;
wire n_39982;
wire n_10277;
wire n_2924;
wire n_31165;
wire n_38630;
wire n_12347;
wire n_5977;
wire n_9065;
wire FE_RN_267_0;
wire n_4499;
wire n_18166;
wire FE_OCP_RBN2976_n_5555;
wire n_125;
wire n_16618;
wire FE_RN_1080_0;
wire n_20942;
wire n_29842;
wire n_6748;
wire n_43400;
wire n_4793;
wire n_11934;
wire n_3263;
wire n_28701;
wire n_23094;
wire n_36904;
wire n_38139;
wire newNet_3153;
wire n_36148;
wire n_9389;
wire n_27736;
wire FE_OCP_RBN2124_n_45224;
wire n_25380;
wire n_43650;
wire FE_OCPN1408_n_672;
wire n_38035;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_14_;
wire n_10225;
wire n_18531;
wire n_28521;
wire n_28949;
wire n_2701;
wire n_36611;
wire delay_add_ln22_unr23_stage9_stallmux_q_18_;
wire newNet_286;
wire n_24622;
wire newNet_3729;
wire n_6544;
wire newNet_1363;
wire n_21615;
wire n_11249;
wire n_28525;
wire n_39284;
wire n_43678;
wire FE_RN_1340_0;
wire n_31111;
wire newNet_309;
wire newNet_226;
wire n_19563;
wire n_25459;
wire FE_RN_416_0;
wire n_4014;
wire n_8985;
wire n_12025;
wire n_28635;
wire n_27160;
wire newNet_771;
wire newNet_2115;
wire n_30380;
wire n_43530;
wire n_34253;
wire n_10933;
wire n_37667;
wire n_41761;
wire n_32636;
wire n_5917;
wire n_17117;
wire newNet_188;
wire n_23571;
wire n_24783;
wire n_31407;
wire n_40841;
wire n_3088;
wire n_16342;
wire n_20418;
wire n_39175;
wire n_40716;
wire n_32568;
wire n_37653;
wire n_4032;
wire n_30901;
wire n_3958;
wire n_28239;
wire n_12746;
wire n_37278;
wire n_9877;
wire n_40130;
wire n_1031;
wire n_16716;
wire n_5287;
wire n_13429;
wire n_867;
wire n_37477;
wire n_28105;
wire n_30737;
wire delay_add_ln22_unr5_stage3_stallmux_q_27_;
wire n_42195;
wire newNet_2731;
wire n_35408;
wire n_40584;
wire beta_22;
wire n_9577;
wire n_21630;
wire newNet_3525;
wire n_5090;
wire n_43882;
wire FE_RN_911_0;
wire n_2859;
wire n_8806;
wire FE_RN_688_0;
wire newNet_3118;
wire n_40170;
wire n_9999;
wire n_16057;
wire n_40715;
wire n_25875;
wire n_5739;
wire n_38182;
wire delay_xor_ln22_unr12_stage5_stallmux_q_15_;
wire FE_RN_1758_0;
wire n_32834;
wire FE_OCP_RBN3540_n_8784;
wire newNet_2157;
wire n_11587;
wire n_36981;
wire n_22861;
wire n_34775;
wire n_2694;
wire FE_RN_992_0;
wire n_7595;
wire n_32139;
wire n_17614;
wire n_24837;
wire n_5662;
wire n_42673;
wire n_8022;
wire n_36631;
wire delay_add_ln22_unr17_stage7_stallmux_q_29_;
wire n_11118;
wire newNet_241;
wire FE_OCPN1050_n_4459;
wire n_21299;
wire n_33828;
wire n_3677;
wire n_15005;
wire newNet_65;
wire n_16142;
wire n_11340;
wire n_24476;
wire n_33815;
wire n_40558;
wire n_27936;
wire n_5131;
wire n_16245;
wire n_28786;
wire newNet_89;
wire n_19658;
wire FE_OCP_RBN1359_FE_RN_677_0;
wire newNet_2261;
wire n_9338;
wire n_33330;
wire n_40929;
wire n_18378;
wire n_24746;
wire n_21350;
wire n_16675;
wire newNet_466;
wire n_4380;
wire FE_RN_1312_0;
wire n_13505;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_9_;
wire n_29415;
wire n_44451;
wire newNet_3111;
wire newNet_3193;
wire n_8787;
wire n_17202;
wire n_40327;
wire n_12292;
wire newNet_2407;
wire FE_RN_72_0;
wire n_15483;
wire n_3066;
wire n_11104;
wire n_25173;
wire n_16398;
wire n_21755;
wire newNet_1629;
wire n_39796;
wire n_33506;
wire n_7814;
wire n_39264;
wire n_15345;
wire n_27472;
wire newNet_636;
wire n_28959;
wire n_37788;
wire n_42887;
wire n_26846;
wire n_15980;
wire n_43043;
wire n_7320;
wire n_36372;
wire n_41366;
wire n_38358;
wire n_10092;
wire n_2408;
wire newNet_2586;
wire n_413;
wire n_10050;
wire n_18760;
wire n_4490;
wire n_32726;
wire n_39098;
wire n_4846;
wire n_41474;
wire n_42199;
wire n_31087;
wire n_35605;
wire n_2911;
wire n_32543;
wire n_36808;
wire FE_RN_1396_0;
wire n_9478;
wire n_1980;
wire n_47256;
wire n_13350;
wire FE_RN_996_0;
wire n_15628;
wire n_25028;
wire n_36176;
wire newNet_1003;
wire n_8726;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_7_;
wire FE_RN_437_0;
wire newNet_778;
wire n_4625;
wire FE_OCP_RBN2422_n_24501;
wire n_18692;
wire FE_OCP_RBN2999_n_11004;
wire newNet_2889;
wire n_497;
wire n_28942;
wire n_13058;
wire n_6974;
wire newNet_1440;
wire newNet_2305;
wire n_10962;
wire n_18206;
wire n_16271;
wire n_25001;
wire n_8337;
wire n_11267;
wire newNet_1420;
wire n_38019;
wire n_13363;
wire n_24939;
wire FE_OCPN1788_n_36034;
wire n_20534;
wire n_24183;
wire n_23308;
wire n_820;
wire n_38870;
wire n_22809;
wire n_10815;
wire n_12173;
wire n_21805;
wire n_33294;
wire n_36664;
wire n_27124;
wire n_38647;
wire n_6889;
wire n_14336;
wire n_21845;
wire n_37796;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_28_;
wire FE_OCP_RBN3630_n_25656;
wire newNet_2952;
wire n_26925;
wire n_21342;
wire newNet_713;
wire newNet_2282;
wire FE_OCP_RBN2419_n_19601;
wire n_12041;
wire n_31632;
wire n_19277;
wire n_31772;
wire n_6610;
wire n_42400;
wire n_14824;
wire delay_xor_ln21_unr12_stage5_stallmux_q_8_;
wire n_9885;
wire n_13518;
wire n_26986;
wire n_38332;
wire n_23580;
wire newNet_151;
wire n_31368;
wire n_28312;
wire n_41449;
wire n_39059;
wire n_27208;
wire delay_add_ln22_unr8_stage4_stallmux_q_14_;
wire delay_add_ln22_unr11_stage5_stallmux_q_17_;
wire n_40410;
wire n_2013;
wire n_23857;
wire n_14678;
wire newNet_671;
wire n_33180;
wire n_16799;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_21_;
wire n_18675;
wire n_5362;
wire n_21483;
wire n_43379;
wire n_6047;
wire n_3319;
wire n_3528;
wire n_15844;
wire n_37431;
wire n_23441;
wire n_29666;
wire n_17058;
wire n_12740;
wire n_21839;
wire n_11743;
wire n_24420;
wire n_5551;
wire n_26938;
wire n_26152;
wire n_5307;
wire n_43194;
wire newNet_2801;
wire FE_OCP_RBN2660_n_9292;
wire n_1336;
wire n_8346;
wire n_25346;
wire n_3042;
wire n_43900;
wire n_25741;
wire n_46226;
wire n_13729;
wire n_7666;
wire newNet_230;
wire FE_OCP_RBN3391_n_37557;
wire n_31871;
wire n_27507;
wire newNet_3532;
wire n_7108;
wire FE_RN_1829_0;
wire n_5859;
wire n_18329;
wire n_35283;
wire delay_xor_ln22_unr6_stage3_stallmux_q_7_;
wire n_39194;
wire n_5549;
wire FE_OCPN1045_n_13570;
wire n_25361;
wire n_28608;
wire n_19867;
wire FE_RN_150_0;
wire n_38377;
wire n_47341;
wire n_8428;
wire n_42972;
wire n_10454;
wire newNet_253;
wire n_13849;
wire newNet_3431;
wire FE_OCP_RBN3382_n_12365;
wire n_7576;
wire n_34037;
wire n_34131;
wire n_35172;
wire newNet_3322;
wire n_10125;
wire n_11602;
wire n_22062;
wire n_33653;
wire n_29646;
wire n_32871;
wire FE_OCPN987_n_28402;
wire n_35655;
wire FE_OCPN963_n_27287;
wire n_25893;
wire n_37459;
wire n_20683;
wire n_8009;
wire n_26976;
wire n_31363;
wire n_24309;
wire n_7283;
wire n_3068;
wire n_30176;
wire n_27152;
wire n_40866;
wire n_16808;
wire n_37021;
wire n_3019;
wire n_30487;
wire n_44336;
wire n_6033;
wire n_22415;
wire FE_RN_217_0;
wire FE_OCP_RBN2825_n_15231;
wire newNet_1881;
wire n_8521;
wire n_9299;
wire n_28766;
wire n_16559;
wire n_20149;
wire n_25152;
wire n_9959;
wire n_18076;
wire n_22028;
wire delay_xor_ln21_unr6_stage3_stallmux_q_11_;
wire n_17350;
wire n_29992;
wire n_39114;
wire n_18331;
wire n_15371;
wire n_43628;
wire n_12994;
wire n_32003;
wire n_40489;
wire n_38907;
wire n_19139;
wire newNet_2986;
wire n_23148;
wire n_21575;
wire n_27072;
wire newNet_1854;
wire FE_RN_1781_0;
wire newNet_1252;
wire n_6290;
wire n_8657;
wire newNet_600;
wire n_33339;
wire n_33067;
wire newNet_1516;
wire n_17274;
wire n_5797;
wire n_15732;
wire n_42487;
wire n_33875;
wire n_11235;
wire delay_xor_ln21_unr3_stage2_stallmux_q_18_;
wire n_42248;
wire n_42259;
wire n_15802;
wire FE_RN_1172_0;
wire n_25596;
wire n_15942;
wire n_29078;
wire n_43083;
wire n_28583;
wire n_45081;
wire n_4667;
wire FE_OCP_RBN1140_n_25816;
wire n_13817;
wire n_33164;
wire n_33595;
wire n_7831;
wire n_31093;
wire n_20764;
wire n_3572;
wire n_30817;
wire n_2531;
wire n_29043;
wire n_40545;
wire FE_OCPN928_n_26231;
wire FE_OCP_RBN2260_n_18899;
wire newNet_358;
wire n_40034;
wire n_40869;
wire n_34398;
wire n_37974;
wire n_24810;
wire n_13715;
wire n_28266;
wire n_20705;
wire n_17499;
wire n_7310;
wire n_23773;
wire FE_OCPN851_n_694;
wire FE_OCP_RBN2402_n_24638;
wire n_37487;
wire n_32234;
wire FE_RN_1671_0;
wire newNet_3668;
wire n_10026;
wire n_31976;
wire n_40240;
wire n_26950;
wire n_34258;
wire n_2324;
wire n_4010;
wire n_7797;
wire n_18864;
wire n_16609;
wire n_19158;
wire n_34196;
wire n_1119;
wire n_16080;
wire n_15124;
wire n_29709;
wire n_38908;
wire n_29740;
wire n_10379;
wire n_16361;
wire newNet_541;
wire n_15977;
wire newNet_3000;
wire n_3663;
wire n_3386;
wire n_31621;
wire n_23091;
wire n_23968;
wire n_22480;
wire FE_OCP_RBN2683_n_35213;
wire n_24884;
wire FE_OFN838_n_4632;
wire FE_RN_620_0;
wire n_35980;
wire n_13787;
wire newNet_3088;
wire n_35651;
wire n_41030;
wire newNet_1904;
wire n_13908;
wire n_24172;
wire FE_OCP_RBN2643_FE_RN_1198_0;
wire n_23419;
wire n_38115;
wire n_28924;
wire n_19991;
wire n_35446;
wire FE_OCP_RBN3380_n_1732;
wire n_13722;
wire n_2809;
wire newNet_3180;
wire newNet_2236;
wire n_25108;
wire n_5372;
wire n_12841;
wire n_7949;
wire n_13546;
wire n_24241;
wire n_4431;
wire n_42546;
wire n_44766;
wire n_4273;
wire n_31702;
wire n_41809;
wire n_30856;
wire n_42025;
wire n_17843;
wire n_16089;
wire newNet_1985;
wire n_10781;
wire delay_add_ln22_unr14_stage6_stallmux_q_13_;
wire n_3998;
wire FE_RN_1646_0;
wire n_8285;
wire n_30469;
wire n_39867;
wire n_2359;
wire n_26688;
wire n_32667;
wire newNet_2424;
wire newNet_1234;
wire n_978;
wire n_14753;
wire n_46414;
wire n_9707;
wire n_22500;
wire n_10303;
wire n_961;
wire n_7199;
wire n_3498;
wire n_13101;
wire n_29379;
wire n_16741;
wire n_23154;
wire n_2989;
wire n_42002;
wire n_2724;
wire n_43792;
wire n_22614;
wire FE_OCPN1478_n_28775;
wire FE_RN_1629_0;
wire n_16022;
wire newNet_1944;
wire newNet_3606;
wire n_17424;
wire n_15390;
wire newNet_972;
wire newNet_395;
wire n_28776;
wire n_26409;
wire n_14136;
wire n_15950;
wire n_8324;
wire n_18338;
wire n_3649;
wire n_13432;
wire n_33023;
wire n_5334;
wire n_1442;
wire n_37992;
wire n_22353;
wire n_19916;
wire n_29864;
wire newNet_723;
wire n_30497;
wire n_24774;
wire n_10857;
wire n_39458;
wire n_42157;
wire n_18738;
wire n_36769;
wire n_26062;
wire FE_RN_1365_0;
wire n_42665;
wire n_12428;
wire FE_RN_1317_0;
wire n_22876;
wire n_37042;
wire n_41915;
wire n_1814;
wire n_17365;
wire n_29348;
wire n_7301;
wire n_10000;
wire n_8060;
wire n_41075;
wire n_24850;
wire n_29624;
wire FE_OCP_RBN3519_n_8498;
wire n_32065;
wire n_42796;
wire FE_OCP_RBN2249_n_13017;
wire n_17069;
wire n_38439;
wire n_7419;
wire n_7224;
wire n_34686;
wire n_5420;
wire n_22822;
wire n_14329;
wire n_25288;
wire n_39749;
wire n_1894;
wire n_1340;
wire n_31184;
wire FE_OCP_RBN2977_n_5555;
wire n_7689;
wire n_15457;
wire n_31244;
wire n_42375;
wire n_8012;
wire n_24435;
wire n_14856;
wire n_32217;
wire n_47199;
wire n_11168;
wire n_11916;
wire n_35934;
wire n_5711;
wire n_12214;
wire n_15324;
wire n_9125;
wire n_35966;
wire n_9215;
wire n_5381;
wire n_26845;
wire n_9161;
wire newNet_2819;
wire n_10975;
wire n_21972;
wire n_28526;
wire n_9612;
wire n_13678;
wire n_40555;
wire newNet_1511;
wire n_27999;
wire n_35826;
wire n_3118;
wire n_10896;
wire n_30440;
wire FE_RN_1632_0;
wire n_20709;
wire FE_OCP_RBN2855_n_10112;
wire n_24193;
wire n_41576;
wire n_16684;
wire n_42121;
wire n_19499;
wire n_599;
wire n_37179;
wire FE_OCPN1043_n_20307;
wire n_34055;
wire n_2754;
wire n_26291;
wire n_23853;
wire n_33405;
wire n_47207;
wire n_35800;
wire n_7743;
wire n_1467;
wire n_1764;
wire newNet_1897;
wire n_19135;
wire n_8631;
wire n_404;
wire n_10604;
wire FE_OCP_RBN2625_n_3848;
wire n_27835;
wire n_12853;
wire FE_OCP_RBN2870_n_10480;
wire n_1101;
wire n_16311;
wire n_42867;
wire n_24486;
wire FE_OCP_RBN3141_n_6477;
wire n_14953;
wire FE_RN_1491_0;
wire n_13608;
wire n_19843;
wire n_3488;
wire n_30019;
wire n_13054;
wire n_5002;
wire n_11637;
wire n_8294;
wire FE_RN_1607_0;
wire n_8939;
wire n_34934;
wire n_5452;
wire n_8718;
wire n_22276;
wire n_41737;
wire n_39493;
wire n_34294;
wire n_43479;
wire n_1493;
wire n_26775;
wire n_39752;
wire n_12413;
wire n_21386;
wire n_26541;
wire n_41850;
wire n_42114;
wire n_25462;
wire n_46995;
wire n_14587;
wire n_10862;
wire n_26595;
wire n_12296;
wire n_44351;
wire n_3813;
wire n_19088;
wire FE_RN_940_0;
wire n_17818;
wire n_27009;
wire n_18661;
wire n_15579;
wire n_17232;
wire n_17390;
wire n_27626;
wire n_1350;
wire n_3673;
wire newNet_1766;
wire n_566;
wire FE_RN_1602_0;
wire n_1122;
wire newNet_2169;
wire n_40153;
wire n_16356;
wire n_30438;
wire FE_RN_1203_0;
wire n_24642;
wire n_5608;
wire n_34898;
wire newNet_1044;
wire n_12525;
wire n_42630;
wire n_36088;
wire n_2074;
wire newNet_2325;
wire n_12279;
wire n_3364;
wire n_5952;
wire n_44174;
wire n_21059;
wire newNet_3633;
wire n_17172;
wire n_21659;
wire n_9658;
wire n_5178;
wire n_29552;
wire n_9436;
wire n_41742;
wire n_14277;
wire n_41197;
wire n_22931;
wire n_25526;
wire n_27045;
wire n_19455;
wire n_31045;
wire newNet_503;
wire n_41455;
wire n_36572;
wire n_43133;
wire FE_RN_575_0;
wire n_33900;
wire n_9873;
wire n_28714;
wire n_38411;
wire FE_OCP_RBN3699_n_43015;
wire n_23317;
wire n_1541;
wire n_17378;
wire n_2355;
wire n_22887;
wire n_28466;
wire n_31288;
wire n_42830;
wire delay_xor_ln21_unr21_stage8_stallmux_q_0_;
wire n_38297;
wire FE_RN_407_0;
wire n_30504;
wire newNet_3542;
wire n_40903;
wire n_10017;
wire FE_OCPN907_n_23227;
wire n_18585;
wire n_24978;
wire FE_RN_770_0;
wire n_33918;
wire n_11817;
wire n_40442;
wire FE_RN_1213_0;
wire n_22303;
wire FE_OCP_DRV_N1569_n_29777;
wire n_7967;
wire FE_OCPN854_n_45450;
wire n_1950;
wire n_1883;
wire n_14795;
wire n_35703;
wire n_18702;
wire n_28122;
wire n_44759;
wire n_6115;
wire n_3150;
wire n_43713;
wire newNet_900;
wire FE_RN_1139_0;
wire FE_OCP_RBN2993_n_35539;
wire n_20238;
wire delay_xor_ln22_unr9_stage4_stallmux_q_4_;
wire n_14479;
wire FE_RN_245_0;
wire newNet_2101;
wire n_9115;
wire n_3706;
wire n_29642;
wire delay_add_ln22_unr27_stage10_stallmux_q_21_;
wire n_14978;
wire n_10150;
wire newNet_1464;
wire n_28420;
wire n_30617;
wire n_41558;
wire FE_OCP_RBN1329_n_18866;
wire n_38380;
wire n_17245;
wire n_42555;
wire FE_OCPN1469_n_23818;
wire n_37815;
wire n_33913;
wire n_6360;
wire n_33961;
wire n_45475;
wire FE_OCP_RBN2703_n_9411;
wire n_1176;
wire n_14433;
wire FE_OCP_RBN3612_FE_OCPN1797_n_20333;
wire newNet_1683;
wire n_2439;
wire n_17975;
wire n_20062;
wire n_28486;
wire newNet_2193;
wire n_8865;
wire n_34185;
wire newNet_344;
wire FE_RN_746_0;
wire n_33836;
wire newNet_897;
wire n_22778;
wire newNet_3296;
wire n_7244;
wire n_33168;
wire newNet_1713;
wire n_38477;
wire n_5384;
wire newNet_495;
wire n_14205;
wire n_7617;
wire delay_xor_ln21_unr6_stage3_stallmux_q_23_;
wire n_8360;
wire n_42006;
wire n_995;
wire n_26885;
wire n_41696;
wire n_38219;
wire newNet_1524;
wire n_12884;
wire n_21527;
wire delay_add_ln22_unr8_stage4_stallmux_q_8_;
wire n_8054;
wire n_4695;
wire n_30522;
wire n_37363;
wire n_36333;
wire newNet_1599;
wire n_29718;
wire n_33440;
wire n_12662;
wire FE_OCP_RBN1166_n_18437;
wire n_39614;
wire n_34845;
wire n_26078;
wire n_31554;
wire FE_RN_844_0;
wire n_34128;
wire n_12888;
wire n_22210;
wire delay_xor_ln21_unr15_stage6_stallmux_q_15_;
wire n_15703;
wire n_37996;
wire n_40221;
wire n_22536;
wire newNet_3602;
wire n_42542;
wire n_8627;
wire n_25197;
wire newNet_3507;
wire n_1329;
wire n_5538;
wire n_2982;
wire n_1652;
wire n_37301;
wire n_47010;
wire n_37330;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_27_;
wire FE_OCPN1252_n_8348;
wire n_26394;
wire n_36764;
wire newNet_2562;
wire newNet_3748;
wire n_12218;
wire n_36979;
wire n_39454;
wire n_44447;
wire n_2775;
wire n_38697;
wire FE_OCP_RBN3504_n_38592;
wire n_5191;
wire n_22337;
wire n_42698;
wire n_22504;
wire newNet_3575;
wire n_2591;
wire n_19824;
wire n_38598;
wire FE_OCP_RBN2751_n_15239;
wire n_39374;
wire n_559;
wire n_46152;
wire n_37776;
wire n_37798;
wire n_26426;
wire n_37902;
wire n_4588;
wire n_42811;
wire n_9610;
wire n_19760;
wire n_4550;
wire n_23158;
wire n_16048;
wire n_24466;
wire newNet_909;
wire n_32340;
wire n_16365;
wire n_36070;
wire n_42661;
wire n_28260;
wire n_29358;
wire newNet_1259;
wire n_38078;
wire FE_RN_196_0;
wire n_15071;
wire n_42327;
wire n_41961;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_31_;
wire n_6664;
wire n_10560;
wire n_7939;
wire n_28042;
wire n_34378;
wire n_28492;
wire n_27215;
wire n_20935;
wire n_13469;
wire newNet_3189;
wire n_345;
wire n_38339;
wire n_38122;
wire newNet_1813;
wire n_31932;
wire n_1572;
wire n_23349;
wire n_6922;
wire n_16308;
wire n_3524;
wire n_8571;
wire n_14647;
wire FE_OCPN1510_n_44174;
wire n_13235;
wire n_19817;
wire n_42691;
wire n_5051;
wire newNet_488;
wire n_6869;
wire newNet_1718;
wire delay_add_ln22_unr11_stage5_stallmux_q_2_;
wire n_39339;
wire n_23555;
wire n_268;
wire n_27630;
wire FE_OCPN968_n_19342;
wire n_36568;
wire n_41375;
wire n_9371;
wire n_9715;
wire n_10680;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_1_;
wire n_30998;
wire n_37644;
wire n_38577;
wire n_3237;
wire n_39256;
wire n_9772;
wire n_14355;
wire n_16480;
wire n_41586;
wire n_36113;
wire FE_RN_1398_0;
wire n_19705;
wire n_24366;
wire n_43261;
wire n_21425;
wire n_35106;
wire n_21240;
wire FE_OCPN3188_n_11012;
wire n_39765;
wire delay_xor_ln21_unr21_stage8_stallmux_q_3_;
wire newNet_1475;
wire n_34082;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_15_;
wire n_39776;
wire newNet_2085;
wire n_21619;
wire n_39976;
wire n_43234;
wire n_26250;
wire newNet_1639;
wire n_22078;
wire FE_RN_1855_0;
wire n_6477;
wire n_17802;
wire n_30603;
wire n_11989;
wire FE_OCPN985_n_25210;
wire n_21014;
wire n_119;
wire n_33084;
wire n_34790;
wire n_17513;
wire n_16260;
wire FE_OCP_RBN1338_n_20941;
wire n_29142;
wire n_16160;
wire n_17480;
wire n_7121;
wire n_31958;
wire n_34372;
wire n_29014;
wire n_7494;
wire n_2483;
wire n_39369;
wire FE_RN_528_0;
wire n_2969;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_0_;
wire newNet_1452;
wire n_22138;
wire n_17796;
wire n_18057;
wire newNet_3359;
wire FE_OCP_RBN2423_n_24501;
wire n_14421;
wire n_19232;
wire n_32461;
wire n_37294;
wire n_42441;
wire n_32431;
wire n_7919;
wire n_11291;
wire FE_OCP_RBN3550_n_44575;
wire n_25219;
wire n_40729;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_12_;
wire n_29392;
wire n_30651;
wire n_16546;
wire n_37107;
wire FE_OCP_RBN2540_n_8781;
wire FE_RN_732_0;
wire n_30274;
wire n_30947;
wire FE_OFN819_n_4298;
wire n_31267;
wire n_1936;
wire n_23545;
wire newNet_2346;
wire n_3920;
wire n_36210;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_0_;
wire n_8145;
wire n_19692;
wire n_19506;
wire n_11502;
wire newNet_3406;
wire FE_RN_1679_0;
wire n_5449;
wire n_46205;
wire n_24920;
wire delay_add_ln22_unr11_stage5_stallmux_q_13_;
wire n_36876;
wire FE_RN_308_0;
wire newNet_1918;
wire n_25918;
wire newNet_2026;
wire n_32383;
wire n_16973;
wire n_2805;
wire n_5913;
wire n_18238;
wire n_40313;
wire n_20200;
wire n_22015;
wire n_6633;
wire n_29003;
wire n_9926;
wire n_28631;
wire n_22661;
wire n_39668;
wire FE_OCP_RBN2826_FE_RN_1573_0;
wire FE_RN_187_0;
wire n_634;
wire n_20104;
wire n_38420;
wire n_10465;
wire n_7587;
wire n_20257;
wire n_28851;
wire n_7442;
wire n_28864;
wire n_11349;
wire newNet_3163;
wire n_43707;
wire n_9247;
wire FE_RN_1096_0;
wire newNet_933;
wire FE_OCP_RBN2562_n_34905;
wire newNet_2095;
wire n_7914;
wire n_7564;
wire newNet_415;
wire n_3548;
wire n_11395;
wire newNet_2702;
wire n_26335;
wire n_36159;
wire n_4072;
wire n_10139;
wire n_40955;
wire n_33636;
wire n_12471;
wire n_13459;
wire n_24793;
wire n_7934;
wire n_40403;
wire FE_OCP_RBN2342_FE_OCPN870_n_2737;
wire n_20881;
wire n_18105;
wire n_12372;
wire FE_OCP_RBN1215_n_20595;
wire n_4631;
wire FE_OCPN866_n_45697;
wire FE_RN_994_0;
wire n_41129;
wire newNet_2179;
wire n_21546;
wire n_30182;
wire FE_OCP_RBN2597_n_25181;
wire n_27705;
wire n_32251;
wire n_42416;
wire FE_RN_1065_0;
wire n_546;
wire n_21246;
wire n_39144;
wire n_37608;
wire n_25495;
wire n_36538;
wire n_8372;
wire n_4811;
wire n_38995;
wire n_1476;
wire n_8495;
wire n_12531;
wire n_25409;
wire FE_OCP_RBN2326_n_29378;
wire n_37025;
wire n_6185;
wire n_11676;
wire n_27986;
wire n_12691;
wire n_26750;
wire n_42381;
wire n_46364;
wire n_32079;
wire n_40139;
wire n_25511;
wire n_16827;
wire n_21764;
wire n_18607;
wire n_25139;
wire n_18192;
wire n_13643;
wire n_6453;
wire n_12697;
wire n_27144;
wire n_43110;
wire n_34675;
wire n_13163;
wire n_35993;
wire n_40008;
wire n_3570;
wire n_27267;
wire n_20853;
wire n_21879;
wire n_26539;
wire n_12990;
wire n_5540;
wire n_19175;
wire n_7163;
wire n_38828;
wire n_2813;
wire n_10635;
wire n_31133;
wire newNet_1964;
wire FE_OCPN1456_n_18860;
wire n_8358;
wire n_11137;
wire n_276;
wire n_5140;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_20_;
wire n_45067;
wire n_816;
wire n_34536;
wire FE_OCP_RBN3055_n_39913;
wire n_38852;
wire n_13748;
wire n_37894;
wire n_7483;
wire FE_OCP_RBN1712_n_21087;
wire n_5479;
wire n_38715;
wire n_2044;
wire n_29686;
wire newNet_2794;
wire n_42083;
wire newNet_1567;
wire n_2545;
wire n_27400;
wire n_22110;
wire FE_OCP_RBN2563_n_34905;
wire FE_RN_573_0;
wire newNet_950;
wire n_12243;
wire n_4304;
wire n_5756;
wire n_20575;
wire n_5759;
wire n_28509;
wire n_34568;
wire n_18689;
wire n_16853;
wire n_31529;
wire n_17022;
wire n_35764;
wire n_248;
wire n_11799;
wire n_24195;
wire n_24042;
wire n_32062;
wire newNet_2552;
wire n_12283;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_6_;
wire n_21911;
wire n_7155;
wire n_5793;
wire n_5740;
wire n_15524;
wire n_16761;
wire n_35553;
wire n_3859;
wire n_16205;
wire delay_xor_ln21_unr9_stage4_stallmux_q_20_;
wire n_18808;
wire n_25253;
wire FE_OCP_RBN1729_n_20903;
wire n_27698;
wire n_144;
wire FE_RN_1216_0;
wire n_11274;
wire n_13570;
wire n_15639;
wire n_4769;
wire n_37589;
wire n_43570;
wire n_10619;
wire n_12756;
wire FE_OCPN910_n_43022;
wire newNet_1061;
wire n_21035;
wire n_695;
wire newNet_1383;
wire n_44032;
wire n_35501;
wire n_6454;
wire n_29128;
wire n_5708;
wire n_37400;
wire n_32173;
wire n_28302;
wire n_8896;
wire n_38981;
wire n_33492;
wire n_21416;
wire n_42742;
wire n_11360;
wire n_39187;
wire n_46218;
wire n_42358;
wire n_21484;
wire FE_OFN615_n_36594;
wire n_8946;
wire n_1133;
wire newNet_2009;
wire n_33818;
wire n_27671;
wire n_5746;
wire n_12082;
wire n_21780;
wire n_30207;
wire n_5655;
wire n_25398;
wire n_29310;
wire n_13929;
wire n_8186;
wire n_24506;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_1_;
wire n_29678;
wire n_37767;
wire n_25057;
wire n_37155;
wire newNet_1457;
wire n_9741;
wire n_37066;
wire n_37527;
wire n_43873;
wire n_33419;
wire n_30406;
wire n_1272;
wire FE_RN_918_0;
wire n_39544;
wire n_25980;
wire n_19057;
wire n_14088;
wire n_39558;
wire n_23751;
wire n_2051;
wire n_3864;
wire n_18914;
wire n_8463;
wire n_27765;
wire newNet_1841;
wire n_6595;
wire n_18581;
wire n_15219;
wire n_42954;
wire n_38594;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_30_;
wire FE_OCP_RBN3609_n_14905;
wire n_42800;
wire n_8206;
wire n_40212;
wire delay_xor_ln22_unr9_stage4_stallmux_q_20_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_7_;
wire n_18266;
wire n_21854;
wire n_36241;
wire newNet_1823;
wire n_44084;
wire n_1604;
wire n_36325;
wire newNet_2875;
wire FE_OCP_RBN3844_FE_RN_1242_0;
wire n_40572;
wire n_15986;
wire n_31453;
wire n_3390;
wire n_32683;
wire n_10477;
wire n_22704;
wire newNet_3023;
wire n_29525;
wire n_37003;
wire FE_OCP_RBN3705_n_11146;
wire n_15724;
wire n_24673;
wire n_15849;
wire n_11193;
wire n_4229;
wire FE_OCP_RBN2788_n_4294;
wire FE_RN_1719_0;
wire n_14370;
wire n_43093;
wire n_5014;
wire n_24458;
wire n_44432;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_12_;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_0_;
wire n_28590;
wire n_1167;
wire FE_OCP_RBN2195_n_2103;
wire n_33953;
wire n_41100;
wire n_10535;
wire n_24068;
wire n_2066;
wire n_33129;
wire delay_xor_ln22_unr3_stage2_stallmux_q_15_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_3_;
wire n_2793;
wire n_36922;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_8_;
wire n_1396;
wire n_11075;
wire n_36988;
wire newNet_3739;
wire n_39889;
wire n_3021;
wire n_26907;
wire n_6882;
wire n_25445;
wire n_9506;
wire n_9483;
wire n_16453;
wire n_2313;
wire n_21126;
wire n_43220;
wire newNet_3596;
wire n_32109;
wire n_4494;
wire newNet_2585;
wire n_8165;
wire n_30117;
wire FE_RN_781_0;
wire n_33850;
wire n_42254;
wire n_46185;
wire n_9030;
wire n_20156;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_15_;
wire n_37952;
wire newNet_2968;
wire delay_xor_ln22_unr6_stage3_stallmux_q_25_;
wire newNet_853;
wire n_17101;
wire n_1649;
wire n_6946;
wire n_3224;
wire n_18997;
wire FE_OCP_RBN1331_n_18866;
wire n_15271;
wire n_38782;
wire n_20589;
wire n_33360;
wire n_33412;
wire n_1920;
wire n_26530;
wire n_27359;
wire newNet_3708;
wire n_38404;
wire n_1870;
wire n_32019;
wire n_42614;
wire n_16256;
wire FE_OCP_RBN3552_n_44575;
wire n_27588;
wire n_14818;
wire FE_RN_368_0;
wire n_2227;
wire n_18610;
wire delay_xor_ln22_unr9_stage4_stallmux_q_7_;
wire n_9036;
wire n_14503;
wire n_33830;
wire n_34148;
wire n_27424;
wire n_32357;
wire FE_OCP_RBN3857_FE_RN_779_0;
wire n_35795;
wire n_42622;
wire sin_out_2;
wire n_6707;
wire n_21886;
wire n_17540;
wire n_13690;
wire n_2836;
wire n_32632;
wire newNet_481;
wire n_21451;
wire n_9017;
wire n_1697;
wire n_285;
wire n_5317;
wire n_40339;
wire n_38304;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_9_;
wire newNet_221;
wire n_45;
wire n_34628;
wire n_32552;
wire n_42394;
wire n_24903;
wire n_43318;
wire n_29427;
wire n_44104;
wire newNet_435;
wire n_28213;
wire FE_RN_1125_0;
wire FE_OFN801_n_46285;
wire n_24201;
wire n_37741;
wire n_22756;
wire newNet_814;
wire n_9796;
wire n_32027;
wire n_29091;
wire FE_RN_333_0;
wire n_46190;
wire n_42188;
wire n_10507;
wire n_27460;
wire n_30025;
wire n_8714;
wire n_12201;
wire FE_OCP_RBN3109_n_43711;
wire n_13940;
wire n_10788;
wire n_28389;
wire n_40512;
wire FE_RN_314_0;
wire n_29746;
wire n_27642;
wire n_40988;
wire n_16802;
wire n_4945;
wire n_39427;
wire n_80;
wire n_16441;
wire n_30017;
wire delay_xor_ln22_unr6_stage3_stallmux_q_9_;
wire FE_RN_1392_0;
wire n_26765;
wire FE_OCP_RBN3717_n_39913;
wire newNet_2524;
wire newNet_1371;
wire n_14040;
wire n_15892;
wire delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire n_14080;
wire n_24091;
wire n_31118;
wire n_20558;
wire n_20001;
wire n_19369;
wire n_35882;
wire n_37133;
wire n_23077;
wire n_22178;
wire n_8490;
wire n_44769;
wire n_32301;
wire n_25656;
wire FE_RN_1725_0;
wire n_272;
wire n_40012;
wire n_25808;
wire n_16407;
wire newNet_1122;
wire n_3893;
wire n_8100;
wire n_32754;
wire delay_add_ln22_unr11_stage5_stallmux_q_11_;
wire n_17851;
wire n_18097;
wire n_39767;
wire n_35879;
wire FE_OCP_RBN2954_n_26231;
wire n_31828;
wire newNet_198;
wire n_34107;
wire n_3886;
wire n_27852;
wire n_11525;
wire n_29656;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_29_;
wire n_22692;
wire n_27364;
wire n_33250;
wire n_6244;
wire n_17323;
wire n_25021;
wire FE_RN_1619_0;
wire newNet_2852;
wire n_35630;
wire n_39011;
wire n_12718;
wire n_2216;
wire n_7903;
wire n_38271;
wire n_38551;
wire FE_OCP_RBN2943_n_5454;
wire FE_RN_834_0;
wire n_34982;
wire n_321;
wire n_27503;
wire n_5564;
wire n_29690;
wire n_24574;
wire FE_RN_284_0;
wire n_1174;
wire FE_RN_486_0;
wire newNet_3127;
wire n_35698;
wire n_25786;
wire n_15880;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_27_;
wire newNet_3346;
wire n_24252;
wire n_39801;
wire delay_xor_ln22_unr9_stage4_stallmux_q_14_;
wire n_22754;
wire n_35905;
wire FE_RN_432_0;
wire n_17731;
wire n_7942;
wire n_17717;
wire n_11150;
wire n_25553;
wire n_2125;
wire n_11774;
wire FE_OCP_RBN2933_n_31010;
wire n_15500;
wire n_30627;
wire n_17567;
wire FE_RN_1487_0;
wire FE_RN_1057_0;
wire n_872;
wire FE_RN_348_0;
wire n_1300;
wire n_3846;
wire FE_OCP_RBN3735_n_31819;
wire n_45814;
wire n_19731;
wire n_43755;
wire n_3244;
wire n_24897;
wire n_23237;
wire n_39246;
wire n_32611;
wire n_16751;
wire n_37559;
wire FE_RN_1223_0;
wire n_30149;
wire n_12186;
wire n_31487;
wire FE_RN_1351_0;
wire n_42869;
wire FE_OCP_RBN2381_n_3502;
wire n_18577;
wire n_30682;
wire n_38775;
wire n_41861;
wire n_19852;
wire n_34859;
wire newNet_323;
wire n_35382;
wire n_3175;
wire n_28833;
wire n_13531;
wire n_43831;
wire n_25696;
wire n_21960;
wire n_39715;
wire n_656;
wire n_30964;
wire n_1772;
wire FE_OCPN1251_n_8210;
wire rst;
wire n_47022;
wire newNet_211;
wire n_38010;
wire n_18219;
wire FE_OCP_RBN3101_n_22504;
wire n_24037;
wire n_35020;
wire n_16757;
wire n_31459;
wire n_35573;
wire n_28003;
wire n_13718;
wire n_21582;
wire n_44045;
wire n_24284;
wire n_20496;
wire newNet_1335;
wire n_29253;
wire n_40708;
wire n_43631;
wire n_34942;
wire n_35718;
wire delay_xor_ln22_unr15_stage6_stallmux_q_10_;
wire n_33273;
wire n_3645;
wire n_22392;
wire FE_RN_330_0;
wire n_670;
wire n_21176;
wire n_21268;
wire n_32977;
wire n_28129;
wire n_46981;
wire n_5217;
wire newNet_2694;
wire n_4330;
wire n_29180;
wire newNet_658;
wire n_30720;
wire n_28188;
wire n_180;
wire n_25407;
wire n_47174;
wire n_32575;
wire n_22560;
wire n_40289;
wire n_15547;
wire n_40255;
wire n_612;
wire newNet_3520;
wire n_19664;
wire n_20546;
wire n_20320;
wire newNet_3487;
wire n_12549;
wire n_3195;
wire n_34755;
wire n_32854;
wire n_34019;
wire n_4423;
wire n_29201;
wire n_6909;
wire n_13842;
wire n_17167;
wire FE_OCP_RBN2481_n_14270;
wire n_43663;
wire FE_OCP_RBN2457_n_13765;
wire n_24267;
wire n_7525;
wire n_7464;
wire n_43056;
wire newNet_1870;
wire n_17939;
wire n_1065;
wire n_15901;
wire n_2131;
wire n_13314;
wire n_27646;
wire n_17174;
wire n_40030;
wire n_1030;
wire n_3975;
wire n_29705;
wire n_41171;
wire newNet_1097;
wire n_23670;
wire n_3372;
wire n_2865;
wire n_1257;
wire FE_OCPN1013_n_41478;
wire n_35333;
wire n_42753;
wire n_33060;
wire n_44057;
wire n_7430;
wire n_1877;
wire n_19934;
wire n_22634;
wire n_28997;
wire n_32347;
wire n_22492;
wire newNet_693;
wire n_22899;
wire sin_out_31;
wire n_20333;
wire n_28807;
wire n_18336;
wire n_966;
wire newNet_3537;
wire newNet_1551;
wire n_19834;
wire newNet_514;
wire n_41185;
wire n_29759;
wire n_18821;
wire n_27570;
wire n_42839;
wire n_8406;
wire n_34803;
wire n_37373;
wire newNet_1107;
wire n_3580;
wire n_41820;
wire n_38009;
wire FE_RN_350_0;
wire newNet_3343;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_28_;
wire n_25084;
wire n_10424;
wire n_25203;
wire n_22829;
wire FE_OCPN856_n_20367;
wire newNet_3062;
wire n_17836;
wire n_26936;
wire n_14472;
wire n_32220;
wire newNet_3648;
wire newNet_948;
wire n_27601;
wire n_29050;
wire n_7639;
wire FE_RN_714_0;
wire FE_RN_1859_0;
wire newNet_14;
wire n_17598;
wire n_36626;
wire n_38615;
wire n_39356;
wire n_42095;
wire n_43779;
wire FE_OCP_RBN2921_n_31107;
wire newNet_133;
wire n_35922;
wire FE_RN_1168_0;
wire n_42463;
wire newNet_3395;
wire n_2614;
wire n_26087;
wire n_13212;
wire n_2502;
wire n_9234;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_14_;
wire n_6052;
wire n_26865;
wire n_33625;
wire n_39853;
wire FE_OCP_DRV_N1559_n_34288;
wire n_20523;
wire FE_RN_1816_0;
wire n_28083;
wire n_18560;
wire n_24868;
wire n_17084;
wire n_11752;
wire n_1973;
wire n_34209;
wire n_43499;
wire n_29812;
wire n_38652;
wire n_15076;
wire n_16462;
wire FE_OCP_RBN2583_n_3734;
wire n_18140;
wire n_35453;
wire n_31538;
wire n_22445;
wire FE_RN_907_0;
wire n_14966;
wire newNet_2787;
wire n_29341;
wire n_12675;
wire n_24546;
wire n_19051;
wire n_26484;
wire FE_OCP_RBN2812_n_15433;
wire FE_RN_41_0;
wire n_11842;
wire n_2844;
wire n_34712;
wire newNet_172;
wire n_13297;
wire n_24248;
wire newNet_3410;
wire FE_OCPN1410_n_27014;
wire newNet_2653;
wire FE_OCPN859_n_12880;
wire n_13878;
wire n_39083;
wire n_3987;
wire n_30121;
wire n_31532;
wire FE_OCP_RBN3268_n_45224;
wire newNet_820;
wire n_1150;
wire n_21697;
wire n_31026;
wire n_18512;
wire n_28705;
wire n_5221;
wire newNet_2299;
wire n_32032;
wire n_10384;
wire n_17916;
wire n_18858;
wire FE_RN_1693_0;
wire n_33781;
wire n_14727;
wire n_14682;
wire delay_xor_ln22_unr3_stage2_stallmux_q_27_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_21_;
wire n_24179;
wire n_23886;
wire n_4464;
wire n_17952;
wire n_29188;
wire n_27622;
wire newNet_55;
wire n_43567;
wire n_34406;
wire n_17449;
wire n_29424;
wire n_33001;
wire n_35204;
wire n_2747;
wire n_10485;
wire FE_OCP_RBN2280_n_24199;
wire delay_xor_ln21_unr3_stage2_stallmux_q_19_;
wire n_33534;
wire n_41289;
wire FE_OCP_RBN2619_n_44561;
wire newNet_3386;
wire n_36991;
wire n_25430;
wire n_8545;
wire newNet_1380;
wire newNet_2430;
wire newNet_1311;
wire n_19709;
wire n_19744;
wire newNet_1112;
wire n_36378;
wire n_28092;
wire n_6499;
wire n_42361;
wire n_25583;
wire n_4555;
wire n_17147;
wire n_23456;
wire n_15968;
wire n_42032;
wire n_7889;
wire n_37708;
wire newNet_2484;
wire n_4203;
wire n_5028;
wire FE_RN_898_0;
wire n_18814;
wire FE_RN_894_0;
wire n_23470;
wire n_26512;
wire delay_sub_ln23_0_unr1_stage2_stallmux_q_1_;
wire n_9464;
wire FE_OCPN1777_n_37744;
wire n_35194;
wire n_21732;
wire newNet_2057;
wire n_33241;
wire n_15602;
wire n_753;
wire newNet_3610;
wire n_4603;
wire n_9471;
wire n_43784;
wire n_30749;
wire n_8817;
wire n_18116;
wire n_18443;
wire n_11998;
wire n_28208;
wire n_1564;
wire n_42150;
wire n_30640;
wire n_32207;
wire n_40971;
wire newNet_3661;
wire n_15025;
wire n_34318;
wire n_6994;
wire n_12124;
wire n_25826;
wire n_24046;
wire n_15866;
wire n_8027;
wire n_13143;
wire n_17191;
wire n_11201;
wire n_32647;
wire n_13479;
wire n_26358;
wire n_30460;
wire n_4245;
wire n_11478;
wire n_30401;
wire newNet_1141;
wire n_18156;
wire newNet_2111;
wire n_11257;
wire newNet_78;
wire n_34699;
wire n_19737;
wire n_30701;
wire n_41547;
wire n_40952;
wire n_42642;
wire n_5856;
wire n_12917;
wire n_21571;
wire n_30002;
wire n_12446;
wire n_31476;
wire n_1195;
wire delay_xor_ln22_unr6_stage3_stallmux_q_20_;
wire n_19438;
wire n_43745;
wire FE_RN_953_0;
wire n_11886;
wire n_21144;
wire n_16234;
wire n_18257;
wire n_30585;
wire newNet_1219;
wire n_4986;
wire n_43546;
wire n_5462;
wire n_46964;
wire FE_RN_705_0;
wire n_3071;
wire n_14550;
wire n_17710;
wire n_4917;
wire n_12398;
wire n_40263;
wire n_4849;
wire newNet_1747;
wire n_42984;
wire n_43520;
wire n_12587;
wire n_37070;
wire FE_OCP_RBN2616_n_44561;
wire n_18211;
wire n_19335;
wire FE_OCPN1746_n_29420;
wire n_36001;
wire n_6305;
wire n_30832;
wire n_40183;
wire n_43001;
wire newNet_3077;
wire n_46415;
wire n_34498;
wire newNet_3589;
wire n_37534;
wire n_29953;
wire n_17197;
wire newNet_2129;
wire n_23149;
wire n_26249;
wire n_27077;
wire n_980;
wire n_22327;
wire n_37851;
wire n_26048;
wire n_3504;
wire n_36622;
wire n_42973;
wire n_4343;
wire n_4733;
wire n_24879;
wire n_37658;
wire n_29305;
wire n_35506;
wire n_20146;
wire n_41882;
wire FE_RN_1021_0;
wire n_34281;
wire n_701;
wire n_22981;
wire n_12654;
wire n_27368;
wire n_410;
wire n_3414;
wire n_35495;
wire n_7189;
wire n_40436;
wire n_41483;
wire n_9113;
wire n_23479;
wire n_25065;
wire FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire newNet_1638;
wire n_12702;
wire n_30387;
wire n_30785;
wire FE_OCP_RBN2424_n_47023;
wire n_39145;
wire newNet_2726;
wire n_36209;
wire n_40415;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_21_;
wire n_12420;
wire newNet_1199;
wire n_33254;
wire FE_OCP_RBN3393_n_37557;
wire n_24604;
wire n_29889;
wire n_26494;
wire FE_OCP_RBN3045_n_5881;
wire n_43284;
wire n_40823;
wire newNet_961;
wire delay_add_ln22_unr17_stage7_stallmux_q_22_;
wire n_2401;
wire n_15614;
wire n_27440;
wire n_25876;
wire n_34068;
wire newNet_256;
wire n_7542;
wire n_1708;
wire n_12728;
wire FE_RN_879_0;
wire n_25327;
wire FE_OCP_RBN2601_n_34388;
wire FE_OFN747_n_13889;
wire n_33086;
wire n_47273;
wire n_32280;
wire n_7362;
wire n_33066;
wire n_2382;
wire FE_OCP_RBN1148_n_27966;
wire newNet_3332;
wire n_27826;
wire n_36197;
wire n_11283;
wire n_39155;
wire n_28403;
wire n_13931;
wire n_29856;
wire n_22649;
wire n_37506;
wire n_25755;
wire n_7313;
wire n_34653;
wire n_43407;
wire n_4878;
wire FE_OCPN1781_FE_OCP_RBN1701_n_19353;
wire n_25791;
wire n_41175;
wire n_24512;
wire n_4240;
wire n_41207;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_9_;
wire n_39352;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_23_;
wire n_29966;
wire n_20134;
wire n_1553;
wire n_1139;
wire n_32596;
wire newNet_1930;
wire n_36724;
wire n_27027;
wire n_40112;
wire FE_OCP_RBN2406_n_8242;
wire n_6639;
wire n_30307;
wire n_7997;
wire n_11198;
wire n_5048;
wire newNet_1321;
wire n_17114;
wire n_43621;
wire n_28661;
wire FE_OCPN3759_n_2346;
wire n_1681;
wire n_20213;
wire n_25774;
wire n_13563;
wire n_17589;
wire n_32520;
wire n_1024;
wire n_7724;
wire n_13227;
wire n_15685;
wire n_38263;
wire n_28013;
wire FE_RN_671_0;
wire n_578;
wire n_34342;
wire n_4214;
wire n_37387;
wire n_13216;
wire n_13201;
wire n_36227;
wire FE_RN_1070_0;
wire n_16062;
wire n_4702;
wire n_34265;
wire n_23941;
wire n_13733;
wire n_34705;
wire n_9392;
wire n_23296;
wire n_35414;
wire newNet_1869;
wire n_26533;
wire n_27533;
wire n_40858;
wire newNet_1360;
wire n_17153;
wire n_7836;
wire n_43398;
wire n_31198;
wire n_38313;
wire n_17793;
wire n_11914;
wire n_36546;
wire newNet_3715;
wire n_34160;
wire n_40568;
wire newNet_2104;
wire n_29487;
wire n_3852;
wire n_29739;
wire n_37353;
wire n_13249;
wire n_9688;
wire n_26112;
wire n_35092;
wire n_32879;
wire n_28722;
wire delay_xor_ln21_unr12_stage5_stallmux_q_16_;
wire n_44036;
wire n_718;
wire n_34448;
wire n_13702;
wire n_1575;
wire n_3491;
wire n_4170;
wire n_10044;
wire newNet_2381;
wire n_40594;
wire n_6141;
wire n_6980;
wire n_12639;
wire n_24883;
wire newNet_1267;
wire n_36079;
wire n_17907;
wire n_19230;
wire n_14888;
wire newNet_3674;
wire n_17002;
wire n_7295;
wire n_16894;
wire n_33683;
wire n_22855;
wire n_30973;
wire n_29350;
wire n_10323;
wire newNet_1454;
wire n_34795;
wire n_41685;
wire n_32902;
wire FE_RN_691_0;
wire n_37208;
wire n_1786;
wire n_12775;
wire n_15357;
wire FE_OCP_RBN3002_n_10805;
wire n_34140;
wire n_41955;
wire n_10290;
wire n_40735;
wire n_29347;
wire n_28674;
wire n_6531;
wire n_19131;
wire n_27067;
wire n_1746;
wire n_19984;
wire n_22846;
wire n_6220;
wire FE_OCP_RBN2154_n_32772;
wire n_264;
wire n_35533;
wire n_37732;
wire n_1108;
wire n_15637;
wire newNet_3205;
wire n_17694;
wire FE_OCP_RBN2250_n_13017;
wire n_217;
wire newNet_3319;
wire n_21520;
wire n_29040;
wire n_11740;
wire n_9672;
wire n_29216;
wire n_26987;
wire n_41111;
wire n_14989;
wire n_30814;
wire n_34229;
wire n_36961;
wire n_9027;
wire n_2806;
wire n_3155;
wire newNet_1419;
wire FE_OCP_RBN2245_n_13017;
wire n_28566;
wire n_2657;
wire n_6488;
wire n_13242;
wire n_43309;
wire n_452;
wire n_33814;
wire FE_RN_625_0;
wire n_6860;
wire n_44944;
wire n_35463;
wire n_3379;
wire FE_RN_1801_0;
wire n_41494;
wire n_12114;
wire n_3635;
wire n_19339;
wire n_15263;
wire n_26977;
wire n_2171;
wire n_38016;
wire newNet_1542;
wire FE_OCP_RBN2490_n_3338;
wire n_5978;
wire n_21398;
wire n_26033;
wire n_28871;
wire n_2996;
wire n_2781;
wire n_40650;
wire n_39476;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_31_;
wire n_8950;
wire n_32700;
wire n_39599;
wire n_13349;
wire newNet_1040;
wire FE_OCP_RBN2302_n_7817;
wire n_2009;
wire n_44312;
wire n_16774;
wire FE_OCPN3752_n_1448;
wire n_26071;
wire n_2107;
wire n_28773;
wire n_23377;
wire n_31004;
wire n_36363;
wire n_39323;
wire n_42822;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_10_;
wire n_25948;
wire n_7182;
wire n_35518;
wire FE_RN_560_0;
wire n_42766;
wire n_34611;
wire n_1780;
wire n_32330;
wire n_20677;
wire n_27804;
wire n_22430;
wire n_34276;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_4_;
wire n_37787;
wire n_10812;
wire n_12079;
wire n_38389;
wire n_2034;
wire n_23347;
wire n_39793;
wire n_11982;
wire n_30862;
wire n_14957;
wire n_41355;
wire n_29643;
wire n_17977;
wire newNet_134;
wire n_16466;
wire n_34013;
wire n_37513;
wire delay_xor_ln22_unr3_stage2_stallmux_q_25_;
wire n_7022;
wire n_25261;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_16_;
wire n_4161;
wire n_8880;
wire n_45529;
wire n_5457;
wire n_11041;
wire newNet_1227;
wire n_16735;
wire n_19636;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_0_;
wire n_11128;
wire n_26377;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_25_;
wire n_13323;
wire n_31513;
wire FE_RN_317_0;
wire n_9510;
wire n_22029;
wire n_30056;
wire n_1018;
wire n_11497;
wire n_2096;
wire n_10119;
wire n_19403;
wire n_12457;
wire newNet_637;
wire n_4638;
wire n_3734;
wire newNet_2638;
wire n_9223;
wire n_42524;
wire n_951;
wire delay_xor_ln22_unr3_stage2_stallmux_q_6_;
wire n_26266;
wire n_676;
wire n_17779;
wire n_16309;
wire n_38789;
wire n_27929;
wire n_20009;
wire n_26780;
wire n_41889;
wire n_17044;
wire n_39904;
wire n_39395;
wire FE_OCP_RBN2190_n_7346;
wire n_5768;
wire n_36036;
wire n_37748;
wire delay_xor_ln22_unr6_stage3_stallmux_q_12_;
wire n_36468;
wire FE_RN_1194_0;
wire n_8913;
wire n_2026;
wire n_25736;
wire newNet_2909;
wire n_18515;
wire n_37877;
wire n_34320;
wire n_17536;
wire n_32004;
wire n_18373;
wire n_2876;
wire n_3551;
wire n_18861;
wire n_36978;
wire n_851;
wire n_45306;
wire n_1934;
wire n_46998;
wire n_18040;
wire n_18136;
wire n_5641;
wire n_36168;
wire n_24813;
wire n_7013;
wire FE_OCP_RBN3206_n_44365;
wire FE_RN_1095_0;
wire n_2593;
wire n_11640;
wire newNet_2081;
wire n_6514;
wire FE_OFN816_n_19885;
wire n_1506;
wire n_37145;
wire n_5207;
wire n_31292;
wire n_21472;
wire FE_RN_547_0;
wire n_17912;
wire newNet_123;
wire n_11939;
wire n_15837;
wire newNet_1594;
wire n_13864;
wire n_3168;
wire n_39208;
wire n_1098;
wire n_38934;
wire n_33034;
wire n_7394;
wire n_40345;
wire n_9323;
wire n_21188;
wire n_28028;
wire n_40145;
wire FE_OCP_RBN2136_n_11907;
wire n_65;
wire newNet_1972;
wire n_9815;
wire n_24565;
wire n_36794;
wire n_16250;
wire n_27687;
wire FE_OCP_RBN2252_n_13017;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_6_;
wire n_22207;
wire n_34207;
wire n_33150;
wire n_620;
wire n_5584;
wire n_8922;
wire n_34051;
wire n_41253;
wire n_25570;
wire n_32924;
wire n_10283;
wire n_23532;
wire n_46379;
wire FE_RN_1244_0;
wire n_2191;
wire n_28227;
wire n_10342;
wire n_6000;
wire n_14562;
wire n_3810;
wire newNet_18;
wire n_10457;
wire newNet_3622;
wire n_28747;
wire n_34596;
wire n_35959;
wire n_1079;
wire n_40003;
wire n_46249;
wire n_11900;
wire n_3477;
wire FE_RN_531_0;
wire n_10548;
wire n_16821;
wire n_36519;
wire n_43180;
wire newNet_3192;
wire n_37343;
wire FE_RN_1851_0;
wire n_3913;
wire n_10328;
wire n_41691;
wire n_40787;
wire newNet_2470;
wire delay_add_ln22_unr27_stage10_stallmux_q_15_;
wire n_8803;
wire n_20196;
wire n_19477;
wire n_24490;
wire n_18186;
wire n_8003;
wire newNet_2847;
wire n_10256;
wire n_29559;
wire n_11892;
wire n_26560;
wire n_34621;
wire n_13667;
wire n_6940;
wire n_3016;
wire n_3511;
wire newNet_2991;
wire n_38748;
wire n_45147;
wire n_3610;
wire n_28825;
wire n_4816;
wire n_15716;
wire n_5359;
wire newNet_2447;
wire newNet_3115;
wire n_13499;
wire n_37912;
wire n_13814;
wire newNet_3221;
wire n_29510;
wire n_17345;
wire n_8276;
wire n_26636;
wire n_25662;
wire n_30433;
wire n_1316;
wire FE_OCPN1005_n_13962;
wire n_43505;
wire n_37724;
wire n_11650;
wire n_40805;
wire n_33993;
wire newNet_1777;
wire n_33382;
wire n_22186;
wire n_31282;
wire n_2196;
wire n_41833;
wire n_31996;
wire n_20529;
wire n_3714;
wire n_661;
wire FE_RN_433_0;
wire n_33570;
wire FE_OCP_RBN2723_n_4219;
wire n_22200;
wire n_16434;
wire FE_RN_1730_0;
wire n_7364;
wire n_19839;
wire n_46242;
wire newNet_3733;
wire n_12809;
wire n_30855;
wire n_3600;
wire n_23581;
wire n_24714;
wire n_36948;
wire n_13628;
wire n_38989;
wire newNet_371;
wire n_33091;
wire n_9604;
wire newNet_1682;
wire n_12501;
wire n_2618;
wire n_31470;
wire n_22740;
wire n_5814;
wire n_20089;
wire FE_OCPN1444_n_45050;
wire n_19418;
wire n_38902;
wire newNet_3032;
wire n_34072;
wire n_11942;
wire n_4799;
wire n_21198;
wire n_21000;
wire n_4857;
wire n_36730;
wire n_10802;
wire n_8013;
wire n_35869;
wire newNet_1328;
wire newNet_2670;
wire n_33621;
wire n_8395;
wire n_8762;
wire n_41367;
wire n_14784;
wire n_38087;
wire n_40775;
wire n_17883;
wire n_19651;
wire n_36177;
wire FE_OCP_RBN3538_n_8597;
wire FE_OCP_DRV_N1597_n_35644;
wire n_26982;
wire n_33119;
wire n_33985;
wire n_35293;
wire n_37569;
wire n_41229;
wire n_3029;
wire n_23110;
wire n_10745;
wire n_27082;
wire newNet_1497;
wire n_26186;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_13_;
wire n_37646;
wire n_20628;
wire n_14943;
wire n_19063;
wire n_9402;
wire n_39506;
wire n_27184;
wire n_14969;
wire n_15039;
wire n_251;
wire newNet_1943;
wire n_33428;
wire FE_OCP_RBN3208_n_44365;
wire newNet_2509;
wire n_21022;
wire n_594;
wire n_20978;
wire n_16865;
wire n_19886;
wire n_4403;
wire FE_OCP_RBN2904_n_10474;
wire n_34472;
wire n_12956;
wire n_34397;
wire FE_RN_850_0;
wire n_32329;
wire n_34193;
wire n_31202;
wire FE_RN_1157_0;
wire n_10185;
wire n_29033;
wire n_2395;
wire FE_OCP_RBN2593_n_25181;
wire n_10797;
wire FE_RN_572_0;
wire n_13488;
wire FE_RN_793_0;
wire n_30556;
wire n_33189;
wire n_39919;
wire n_21566;
wire n_29919;
wire n_31673;
wire FE_OCP_RBN1198_n_30619;
wire n_24236;
wire n_28479;
wire n_25246;
wire n_31039;
wire n_15049;
wire n_40997;
wire n_37824;
wire n_4389;
wire n_38602;
wire n_6013;
wire FE_OCPN1440_n_23339;
wire n_16516;
wire n_25178;
wire n_8645;
wire n_12400;
wire n_12589;
wire n_25426;
wire n_2112;
wire n_34923;
wire n_1828;
wire n_3782;
wire n_23416;
wire n_1400;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_5_;
wire n_32517;
wire n_27352;
wire newNet_912;
wire n_23444;
wire n_40364;
wire n_35475;
wire n_1791;
wire n_26316;
wire n_29870;
wire FE_OCP_RBN2508_n_13896;
wire n_6408;
wire n_29432;
wire n_8480;
wire n_9414;
wire n_19868;
wire n_34048;
wire n_42791;
wire n_20310;
wire n_20810;
wire n_42020;
wire n_11165;
wire newNet_2413;
wire n_1431;
wire n_31988;
wire FE_RN_1605_0;
wire n_29155;
wire n_5323;
wire n_647;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_4_;
wire n_11121;
wire FE_RN_268_0;
wire n_32201;
wire n_35929;
wire n_23161;
wire n_27586;
wire n_2680;
wire n_26445;
wire n_34086;
wire n_4766;
wire n_45755;
wire n_36126;
wire n_34638;
wire n_14898;
wire n_29920;
wire n_34769;
wire n_16563;
wire n_8774;
wire n_18938;
wire delay_add_ln22_unr23_stage9_stallmux_q_9_;
wire n_39812;
wire FE_OCP_RBN3131_n_43762;
wire n_11665;
wire FE_OCP_RBN2654_n_9198;
wire n_46956;
wire n_6214;
wire n_11607;
wire n_41416;
wire n_24766;
wire n_39513;
wire n_13707;
wire n_20871;
wire n_25577;
wire FE_OCP_RBN3111_n_43871;
wire n_478;
wire n_11713;
wire n_39045;
wire n_45516;
wire newNet_2182;
wire n_42994;
wire n_40969;
wire n_37416;
wire n_20963;
wire n_22766;
wire n_5821;
wire n_151;
wire FE_RN_1848_0;
wire n_34136;
wire newNet_140;
wire n_11807;
wire n_7692;
wire n_38758;
wire n_37967;
wire FE_OCP_RBN3097_n_6313;
wire n_527;
wire n_16887;
wire n_47005;
wire n_36276;
wire FE_RN_1741_0;
wire n_36298;
wire n_35252;
wire n_40756;
wire n_5802;
wire n_28816;
wire newNet_3185;
wire n_15123;
wire n_26226;
wire n_13303;
wire n_16991;
wire newNet_1319;
wire FE_OCPN1247_n_43120;
wire beta_12;
wire n_14359;
wire n_25106;
wire FE_OCP_RBN2667_n_4158;
wire n_45321;
wire n_41542;
wire n_33717;
wire n_33898;
wire n_19781;
wire n_44672;
wire FE_OCP_RBN3005_n_11087;
wire n_1869;
wire n_26127;
wire n_19919;
wire n_32493;
wire n_39816;
wire n_28280;
wire n_40868;
wire n_20732;
wire newNet_726;
wire n_3346;
wire n_32721;
wire n_39553;
wire n_9465;
wire FE_OCP_RBN2573_n_29922;
wire n_29637;
wire n_27724;
wire n_18727;
wire n_26670;
wire n_36081;
wire n_18982;
wire n_13612;
wire n_28757;
wire n_991;
wire n_39751;
wire n_166;
wire n_41921;
wire n_32112;
wire n_31562;
wire n_16484;
wire n_39199;
wire n_29229;
wire n_22994;
wire n_24389;
wire n_18888;
wire delay_sub_ln23_0_unr23_stage8_stallmux_q;
wire n_41033;
wire n_8576;
wire n_29861;
wire n_35112;
wire n_40394;
wire n_20767;
wire n_3724;
wire FE_OCPN1434_n_30614;
wire n_2902;
wire n_40382;
wire FE_OCP_RBN3631_n_20504;
wire n_11876;
wire n_14259;
wire FE_OCP_RBN3551_n_44575;
wire n_827;
wire FE_OCPN3181_FE_OCP_RBN2831_n_10198;
wire n_3509;
wire n_26312;
wire n_3594;
wire n_7415;
wire n_25679;
wire n_25027;
wire n_28740;
wire n_36419;
wire n_10409;
wire n_15224;
wire n_2855;
wire newNet_352;
wire n_28899;
wire n_8477;
wire n_40828;
wire FE_RN_1690_0;
wire n_13728;
wire n_7172;
wire n_1994;
wire n_41661;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_14_;
wire newNet_267;
wire n_8491;
wire n_44051;
wire n_31626;
wire n_13310;
wire n_34500;
wire FE_RN_252_0;
wire FE_OCP_RBN2372_n_8221;
wire n_2583;
wire n_7388;
wire n_7472;
wire n_39678;
wire n_14758;
wire n_23779;
wire n_37989;
wire n_39001;
wire FE_OCP_RBN3713_n_31466;
wire n_36888;
wire FE_RN_1319_0;
wire n_26655;
wire n_36841;
wire n_40261;
wire n_23638;
wire n_30203;
wire newNet_2335;
wire n_34428;
wire n_975;
wire FE_OCP_RBN2646_n_47015;
wire n_24612;
wire n_19618;
wire n_34334;
wire n_2541;
wire n_15743;
wire newNet_52;
wire n_15908;
wire newNet_2395;
wire n_38639;
wire newNet_1288;
wire FE_RN_4_0;
wire n_9339;
wire newNet_1701;
wire newNet_393;
wire n_27783;
wire n_22485;
wire n_14911;
wire FE_OCP_RBN2783_n_9859;
wire n_32970;
wire n_10005;
wire newNet_1982;
wire n_30677;
wire n_34118;
wire n_40084;
wire n_44443;
wire n_27868;
wire n_3830;
wire n_9749;
wire n_32412;
wire n_4729;
wire n_36388;
wire FE_OCP_RBN1351_n_19148;
wire n_42071;
wire n_24864;
wire FE_OCP_RBN2979_n_5656;
wire n_21363;
wire n_35354;
wire newNet_3465;
wire n_7985;
wire n_36492;
wire n_4117;
wire n_34521;
wire n_931;
wire n_31748;
wire newNet_1709;
wire n_26192;
wire n_43629;
wire n_21263;
wire n_10527;
wire n_43464;
wire n_26953;
wire n_18052;
wire n_22153;
wire n_43067;
wire n_35441;
wire n_30316;
wire newNet_3002;
wire n_35614;
wire n_12962;
wire n_23032;
wire n_41721;
wire n_5400;
wire n_2986;
wire n_23592;
wire newNet_1725;
wire n_31313;
wire n_5783;
wire n_29793;
wire FE_OCP_RBN2793_n_10106;
wire n_21861;
wire n_31939;
wire n_10170;
wire n_19758;
wire n_19255;
wire n_2200;
wire n_2786;
wire n_207;
wire n_29175;
wire n_42746;
wire n_41746;
wire n_15191;
wire n_1977;
wire n_3606;
wire FE_RN_234_0;
wire n_8321;
wire beta_27;
wire n_35726;
wire n_22399;
wire n_29148;
wire newNet_2924;
wire n_41859;
wire n_27201;
wire n_40944;
wire n_20205;
wire n_31582;
wire n_45825;
wire n_25972;
wire FE_OCPN891_n_7802;
wire FE_OFN799_n_46285;
wire FE_OCP_RBN1138_n_11779;
wire n_33904;
wire n_27654;
wire n_10615;
wire FE_OCP_RBN2968_n_26398;
wire n_27245;
wire FE_OCP_RBN2282_n_29111;
wire n_30343;
wire n_7874;
wire n_24989;
wire n_4876;
wire n_27614;
wire n_1905;
wire newNet_1907;
wire n_6373;
wire n_26143;
wire n_29053;
wire n_13407;
wire n_13029;
wire n_33596;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_7_;
wire n_15747;
wire n_4472;
wire FE_RN_1870_0;
wire n_31255;
wire n_18844;
wire n_2758;
wire n_28535;
wire n_17958;
wire n_31066;
wire n_32227;
wire n_11005;
wire FE_OCPN1786_n_30134;
wire n_28147;
wire n_41044;
wire n_16268;
wire n_41790;
wire FE_RN_194_0;
wire n_33042;
wire FE_OCP_RBN3496_n_13818;
wire n_25890;
wire newNet_2780;
wire n_27499;
wire n_14133;
wire n_23675;
wire FE_OCP_RBN2607_n_3807;
wire n_43848;
wire n_42911;
wire n_9077;
wire n_46939;
wire n_3141;
wire n_17672;
wire FE_OCP_RBN1371_n_20763;
wire n_37662;
wire n_3825;
wire n_5695;
wire n_30371;
wire n_38158;
wire n_45889;
wire n_38733;
wire n_16830;
wire newNet_1838;
wire n_30068;
wire n_29258;
wire n_13974;
wire FE_OCP_RBN2585_n_9009;
wire FE_OCP_RBN2148_FE_OCPN861_n_45450;
wire n_30444;
wire n_12134;
wire n_43701;
wire n_1445;
wire n_40530;
wire n_17334;
wire n_12020;
wire n_1240;
wire n_29450;
wire n_887;
wire FE_OCP_RBN2278_n_24173;
wire n_31705;
wire n_24782;
wire n_18162;
wire n_20269;
wire FE_OCPN885_n_42216;
wire n_3683;
wire n_32662;
wire n_11641;
wire n_31839;
wire n_26279;
wire n_13944;
wire n_24800;
wire FE_OCP_RBN3221_n_22068;
wire n_22446;
wire n_4615;
wire n_13031;
wire n_39294;
wire n_12818;
wire newNet_2491;
wire n_36350;
wire n_33974;
wire n_14480;
wire n_25952;
wire n_27965;
wire n_35341;
wire n_26608;
wire FE_RN_10_0;
wire n_40924;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_16_;
wire n_31908;
wire n_33035;
wire n_40017;
wire n_42354;
wire n_30663;
wire n_8045;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_26_;
wire n_3412;
wire n_42088;
wire n_32953;
wire n_12978;
wire n_4193;
wire n_17963;
wire n_41276;
wire n_14620;
wire n_7435;
wire newNet_2815;
wire n_11405;
wire n_46252;
wire mux_while_ln12_psv_q_8_;
wire n_38174;
wire FE_RN_1482_0;
wire n_11994;
wire newNet_62;
wire n_36861;
wire n_19270;
wire n_20286;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_13_;
wire n_23089;
wire n_1230;
wire n_14689;
wire n_25468;
wire n_19005;
wire n_9956;
wire n_27455;
wire n_32296;
wire n_45224;
wire n_821;
wire n_10210;
wire FE_RN_1383_0;
wire newNet_2498;
wire newNet_2276;
wire newNet_2047;
wire n_43492;
wire n_4053;
wire newNet_2642;
wire n_39429;
wire n_8114;
wire newNet_2693;
wire n_36782;
wire n_40323;
wire n_9420;
wire n_40214;
wire n_14013;
wire n_31271;
wire n_2068;
wire n_2961;
wire n_29362;
wire n_31541;
wire n_37759;
wire n_42164;
wire FE_OCP_RBN3252_delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire n_13004;
wire n_28037;
wire n_43887;
wire n_6765;
wire n_904;
wire newNet_185;
wire n_30890;
wire n_40585;
wire n_36415;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_21_;
wire n_26924;
wire newNet_3692;
wire n_4321;
wire newNet_3274;
wire n_3233;
wire n_19253;
wire n_43021;
wire FE_RN_1055_0;
wire newNet_1486;
wire n_35836;
wire n_39460;
wire n_30621;
wire n_1263;
wire n_21803;
wire FE_OCP_RBN2002_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_26345;
wire n_2721;
wire n_27306;
wire n_1376;
wire n_41788;
wire n_40280;
wire n_734;
wire n_36933;
wire n_10159;
wire n_25602;
wire n_36014;
wire n_2691;
wire n_16411;
wire n_44958;
wire n_41219;
wire n_9735;
wire newNet_824;
wire FE_OCP_RBN3062_FE_RN_640_0;
wire n_16527;
wire n_35697;
wire n_43885;
wire n_1027;
wire n_12579;
wire n_16064;
wire n_43537;
wire n_5905;
wire n_7230;
wire FE_RN_203_0;
wire n_35891;
wire FE_OCP_RBN3837_n_19513;
wire n_25718;
wire n_31518;
wire newNet_2649;
wire n_29897;
wire n_38631;
wire n_16719;
wire newNet_1469;
wire FE_OCP_RBN2582_n_3734;
wire n_5062;
wire n_15592;
wire n_17250;
wire n_31449;
wire newNet_3394;
wire n_8155;
wire n_7334;
wire n_33799;
wire n_7049;
wire n_111;
wire n_73;
wire n_17398;
wire n_31762;
wire n_32124;
wire n_24222;
wire n_33942;
wire n_14295;
wire n_16585;
wire n_37676;
wire FE_OCP_RBN3361_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_RN_1359_0;
wire n_32608;
wire FE_OCP_RBN2579_n_3734;
wire newNet_1443;
wire FE_OCP_RBN2404_n_24638;
wire FE_RN_933_0;
wire n_29490;
wire n_38136;
wire n_11217;
wire n_15515;
wire FE_RN_247_0;
wire n_6203;
wire n_34298;
wire n_41827;
wire FE_RN_1499_0;
wire n_14233;
wire n_42681;
wire FE_OCP_RBN3722_n_39913;
wire n_31417;
wire n_4436;
wire n_2644;
wire n_23740;
wire n_19272;
wire n_2693;
wire n_7521;
wire FE_RN_1288_0;
wire n_1832;
wire n_11071;
wire FE_OCP_RBN2446_n_29684;
wire n_13475;
wire n_26137;
wire newNet_1407;
wire n_19213;
wire n_8855;
wire n_13502;
wire n_23668;
wire n_16833;
wire n_17305;
wire n_6858;
wire n_16535;
wire n_12535;
wire newNet_2266;
wire n_18619;
wire FE_OCPN1506_n_17680;
wire newNet_1669;
wire n_21999;
wire n_3083;
wire n_19594;
wire n_28315;
wire n_16438;
wire n_28159;
wire n_29538;
wire n_29743;
wire newNet_1;
wire n_14055;
wire n_8960;
wire n_3897;
wire n_34656;
wire n_13791;
wire newNet_994;
wire FE_OCP_RBN3632_n_20568;
wire newNet_3135;
wire n_7707;
wire n_30394;
wire n_43691;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_23_;
wire n_4485;
wire n_13299;
wire n_31389;
wire FE_OCP_RBN3004_n_10930;
wire n_27057;
wire n_5928;
wire n_14145;
wire n_35376;
wire n_14636;
wire n_46181;
wire n_13193;
wire n_15347;
wire n_32185;
wire n_12364;
wire n_28956;
wire n_40712;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_12_;
wire n_15055;
wire n_4253;
wire n_28769;
wire n_8504;
wire n_29319;
wire n_4910;
wire n_21808;
wire n_42420;
wire newNet_3686;
wire n_3656;
wire n_43339;
wire delay_add_ln22_unr20_stage8_stallmux_q_20_;
wire FE_OCP_RBN3666_n_10106;
wire FE_OCPN960_n_3951;
wire FE_RN_1460_0;
wire n_38564;
wire n_39252;
wire n_39698;
wire n_42607;
wire n_20643;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_11_;
wire n_27634;
wire n_19743;
wire n_20539;
wire n_28126;
wire n_20093;
wire n_4064;
wire n_30922;
wire n_11357;
wire n_23615;
wire n_41160;
wire FE_OCP_RBN2538_n_3645;
wire n_8676;
wire FE_OCP_RBN2920_n_31107;
wire n_38927;
wire n_20470;
wire n_42551;
wire FE_RN_1367_0;
wire n_35323;
wire n_42110;
wire n_21687;
wire newNet_86;
wire n_34869;
wire n_24757;
wire n_14802;
wire n_35328;
wire n_20415;
wire n_10201;
wire n_39379;
wire n_15918;
wire n_35428;
wire n_40078;
wire n_21517;
wire FE_OCP_RBN2560_n_3437;
wire n_15006;
wire n_31360;
wire n_20016;
wire n_6979;
wire FE_OCP_RBN2239_n_44881;
wire n_13289;
wire n_38156;
wire n_24670;
wire n_20515;
wire n_20056;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_3_;
wire n_38443;
wire n_43590;
wire FE_OCP_RBN2969_n_26398;
wire n_43341;
wire n_370;
wire n_29122;
wire n_22383;
wire n_7135;
wire n_3401;
wire n_37841;
wire n_26059;
wire mux_while_ln12_psv_q_6_;
wire n_1105;
wire n_43689;
wire n_43793;
wire n_42531;
wire FE_OCP_RBN2512_n_19884;
wire n_172;
wire n_35396;
wire newNet_470;
wire n_10416;
wire n_43675;
wire n_24741;
wire n_12176;
wire n_38288;
wire n_23583;
wire n_1142;
wire n_4519;
wire n_6502;
wire n_11681;
wire n_26519;
wire n_18495;
wire n_31091;
wire n_39965;
wire FE_RN_929_0;
wire newNet_2011;
wire n_24963;
wire n_28504;
wire newNet_1021;
wire n_29313;
wire n_3227;
wire n_27511;
wire n_35360;
wire n_664;
wire n_28709;
wire FE_OCP_RBN2537_n_3645;
wire n_23229;
wire n_29092;
wire newNet_738;
wire n_9989;
wire n_17926;
wire n_31059;
wire n_27905;
wire n_11282;
wire n_33206;
wire n_7158;
wire n_41286;
wire newNet_2309;
wire newNet_414;
wire n_29465;
wire FE_OCP_RBN2416_n_8293;
wire n_15651;
wire newNet_1530;
wire n_15667;
wire n_3748;
wire n_43518;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_26_;
wire n_33675;
wire n_27040;
wire n_32746;
wire FE_RN_158_0;
wire n_12155;
wire n_25234;
wire n_10714;
wire n_19538;
wire n_22052;
wire n_24696;
wire n_7412;
wire n_43589;
wire newNet_846;
wire n_30082;
wire newNet_1526;
wire n_33978;
wire n_42558;
wire newNet_2885;
wire n_549;
wire delay_xor_ln22_unr21_stage8_stallmux_q_2_;
wire n_9431;
wire n_7167;
wire n_15135;
wire n_43626;
wire newNet_611;
wire n_24299;
wire n_40491;
wire n_13230;
wire n_29137;
wire n_38887;
wire n_42490;
wire n_5991;
wire n_23409;
wire n_24733;
wire delay_add_ln22_unr8_stage4_stallmux_q_23_;
wire n_14592;
wire FE_OCP_RBN3213_n_44365;
wire n_26240;
wire n_41632;
wire n_37372;
wire n_38430;
wire n_14299;
wire n_7160;
wire n_42590;
wire n_18432;
wire n_8264;
wire n_33882;
wire n_15421;
wire n_7748;
wire n_29835;
wire n_43255;
wire newNet_108;
wire FE_OCP_RBN2311_n_41420;
wire n_13086;
wire n_3032;
wire n_11231;
wire n_2638;
wire n_5620;
wire n_6443;
wire FE_RN_30_0;
wire n_2387;
wire n_3105;
wire n_24993;
wire n_23142;
wire n_653;
wire n_28455;
wire n_15971;
wire n_9193;
wire n_46200;
wire n_38455;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_8_;
wire n_7630;
wire n_16226;
wire n_33704;
wire n_27731;
wire n_33946;
wire newNet_2021;
wire n_28178;
wire n_40784;
wire n_23889;
wire n_18478;
wire n_19111;
wire n_33518;
wire n_9007;
wire newNet_2697;
wire newNet_904;
wire n_31021;
wire n_41421;
wire newNet_2624;
wire n_22486;
wire n_43039;
wire n_17688;
wire n_3214;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_17_;
wire newNet_2225;
wire newNet_1864;
wire n_37703;
wire n_29673;
wire n_38292;
wire n_43645;
wire n_19225;
wire n_41141;
wire n_7054;
wire n_1192;
wire n_52;
wire n_13014;
wire n_17373;
wire n_42048;
wire n_34465;
wire n_9331;
wire n_29756;
wire n_16155;
wire FE_OCP_DRV_N3157_n_27062;
wire n_43025;
wire n_35870;
wire n_21708;
wire n_39890;
wire newNet_1049;
wire n_2965;
wire n_30035;
wire n_34063;
wire n_7931;
wire n_40629;
wire n_32571;
wire n_25631;
wire n_34793;
wire n_29732;
wire FE_RN_900_0;
wire n_2977;
wire n_27518;
wire n_7447;
wire n_33552;
wire n_23948;
wire n_17039;
wire n_34855;
wire n_33777;
wire n_21745;
wire newNet_94;
wire n_7656;
wire n_4713;
wire n_36386;
wire newNet_3312;
wire n_19009;
wire n_5963;
wire n_9166;
wire n_8351;
wire n_16998;
wire n_41381;
wire n_29011;
wire n_7561;
wire FE_OCP_RBN2779_n_15595;
wire n_18811;
wire n_41487;
wire n_23692;
wire n_31301;
wire n_381;
wire n_36985;
wire n_27702;
wire n_15394;
wire newNet_2936;
wire n_43655;
wire n_25825;
wire FE_RN_1124_0;
wire FE_RN_1424_0;
wire n_12983;
wire n_30600;
wire n_35990;
wire FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire FE_OCPN1525_n_26587;
wire FE_OCP_RBN3337_n_44610;
wire n_29930;
wire n_43739;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_22_;
wire n_32961;
wire delay_xor_ln22_unr18_stage7_stallmux_q_3_;
wire newNet_581;
wire FE_RN_755_0;
wire newNet_439;
wire n_11130;
wire newNet_1584;
wire FE_OCP_RBN3020_n_39942;
wire n_18897;
wire n_34284;
wire n_5565;
wire n_15969;
wire n_23627;
wire FE_OCPN906_n_44561;
wire n_30014;
wire n_33560;
wire n_24058;
wire n_30322;
wire newNet_1376;
wire FE_OCP_RBN3571_n_44563;
wire n_34358;
wire n_43268;
wire n_40679;
wire n_9617;
wire delay_add_ln22_unr11_stage5_stallmux_q_3_;
wire n_21497;
wire n_32409;
wire n_23439;
wire n_25250;
wire FE_OCP_RBN3128_n_32266;
wire n_5612;
wire n_1909;
wire n_35279;
wire n_22081;
wire n_41925;
wire n_7519;
wire n_43394;
wire n_45185;
wire newNet_3454;
wire n_34586;
wire n_33090;
wire n_2365;
wire newNet_2092;
wire n_27403;
wire newNet_2056;
wire n_15083;
wire n_36427;
wire n_12632;
wire n_22442;
wire cos_out_25;
wire n_2538;
wire n_12099;
wire n_42805;
wire n_24322;
wire newNet_3595;
wire n_12007;
wire n_43761;
wire n_19954;
wire n_32049;
wire n_28849;
wire n_39078;
wire FE_RN_315_0;
wire FE_RN_83_0;
wire n_12774;
wire n_32210;
wire n_27540;
wire n_1393;
wire delay_xor_ln22_unr18_stage7_stallmux_q_2_;
wire n_16418;
wire n_32586;
wire n_2714;
wire FE_RN_1268_0;
wire FE_RN_1252_0;
wire n_20799;
wire newNet_142;
wire n_36203;
wire FE_OCP_RBN2775_n_10100;
wire n_15520;
wire n_30953;
wire newNet_2618;
wire n_34291;
wire n_25091;
wire n_34965;
wire newNet_969;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_8_;
wire FE_OCP_RBN3052_n_39913;
wire n_24808;
wire n_18392;
wire n_23882;
wire n_13639;
wire n_5399;
wire n_8891;
wire n_42117;
wire n_1057;
wire newNet_1751;
wire newNet_3398;
wire n_31445;
wire n_9158;
wire n_23205;
wire n_32997;
wire FE_OCP_RBN2320_n_2382;
wire n_45619;
wire n_7559;
wire newNet_3288;
wire delay_add_ln22_unr2_stage2_stallmux_q_1_;
wire n_28471;
wire FE_OCP_RBN2926_n_16446;
wire n_25117;
wire n_16685;
wire FE_OCP_RBN2841_n_4784;
wire n_13793;
wire n_13358;
wire n_24532;
wire n_19794;
wire n_34005;
wire n_27485;
wire n_16595;
wire n_36021;
wire n_8906;
wire n_40699;
wire n_35167;
wire newNet_2004;
wire n_21102;
wire n_8893;
wire n_35015;
wire n_44216;
wire delay_add_ln22_unr20_stage8_stallmux_q_10_;
wire n_43372;
wire n_14566;
wire n_15527;
wire n_20666;
wire n_35037;
wire n_34927;
wire n_6680;
wire n_8355;
wire n_13519;
wire n_28690;
wire FE_OCP_RBN1370_n_20763;
wire n_109;
wire n_725;
wire FE_OCP_RBN2880_n_21132;
wire n_24859;
wire n_41563;
wire newNet_273;
wire n_5060;
wire n_14605;
wire n_4301;
wire n_29047;
wire n_9531;
wire n_19812;
wire n_3536;
wire newNet_442;
wire n_13383;
wire n_25036;
wire n_19933;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_13_;
wire FE_RN_927_0;
wire n_36158;
wire n_13622;
wire FE_OCP_RBN2693_n_15083;
wire n_19494;
wire n_40488;
wire n_37413;
wire newNet_2539;
wire n_15571;
wire n_26178;
wire n_6121;
wire n_35125;
wire n_26502;
wire newNet_3199;
wire n_12092;
wire n_4024;
wire newNet_3566;
wire n_37935;
wire n_9657;
wire n_22306;
wire n_4156;
wire n_4509;
wire n_13805;
wire delay_xor_ln22_unr12_stage5_stallmux_q_13_;
wire n_42589;
wire n_3200;
wire newNet_808;
wire FE_RN_211_0;
wire FE_RN_1171_0;
wire n_3230;
wire n_19621;
wire n_9543;
wire n_17450;
wire n_24463;
wire n_25675;
wire n_1544;
wire n_5866;
wire n_9633;
wire n_32911;
wire n_11966;
wire n_22109;
wire n_43030;
wire n_39249;
wire n_4398;
wire n_8965;
wire delay_xor_ln21_unr3_stage2_stallmux_q_1_;
wire FE_RN_696_0;
wire FE_OCP_RBN2472_n_8664;
wire n_20117;
wire n_34783;
wire n_27914;
wire n_38591;
wire n_13436;
wire n_18425;
wire n_26719;
wire n_3444;
wire n_31524;
wire n_29287;
wire n_4699;
wire n_5531;
wire n_35162;
wire FE_OCPN997_n_44460;
wire FE_OCP_RBN1840_n_19528;
wire FE_OCP_RBN2758_FE_RN_722_0;
wire n_27560;
wire n_21301;
wire n_37881;
wire n_23126;
wire n_420;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_12_;
wire n_2521;
wire n_704;
wire n_23112;
wire n_16003;
wire n_45815;
wire n_11061;
wire n_25903;
wire n_2466;
wire n_19521;
wire FE_OCP_RBN3076_FE_OFN807_n_46195;
wire n_6927;
wire n_25547;
wire n_41220;
wire newNet_2688;
wire n_36505;
wire n_42307;
wire n_22965;
wire n_14716;
wire n_36083;
wire n_39746;
wire n_43348;
wire n_21956;
wire n_26897;
wire n_29436;
wire n_36670;
wire n_7260;
wire n_12187;
wire n_5350;
wire n_1409;
wire n_26772;
wire n_33760;
wire n_37771;
wire newNet_2232;
wire n_4241;
wire n_12461;
wire n_39532;
wire n_30727;
wire n_22517;
wire n_5435;
wire n_35512;
wire newNet_2919;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_18_;
wire newNet_838;
wire newNet_2902;
wire n_28004;
wire n_42968;
wire newNet_2165;
wire FE_OFN753_n_44461;
wire n_19119;
wire n_18911;
wire n_31840;
wire n_27391;
wire n_29004;
wire n_19851;
wire n_7863;
wire n_8225;
wire newNet_498;
wire n_6900;
wire FE_OCP_RBN3823_n_44061;
wire n_21963;
wire n_13642;
wire n_1623;
wire n_18555;
wire n_24826;
wire n_6169;
wire n_24121;
wire n_20122;
wire n_21552;
wire n_21562;
wire n_17326;
wire n_32057;
wire n_18068;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_22_;
wire n_43540;
wire newNet_2755;
wire n_38228;
wire n_43016;
wire FE_OCP_RBN3546_n_44575;
wire n_30654;
wire n_20694;
wire n_15678;
wire n_21256;
wire FE_RN_731_0;
wire n_21918;
wire n_36164;
wire n_41529;
wire FE_OCP_RBN2820_n_4872;
wire n_20019;
wire delay_xor_ln21_unr9_stage4_stallmux_q_4_;
wire n_20439;
wire n_28886;
wire n_1125;
wire FE_RN_669_0;
wire n_8626;
wire n_15212;
wire n_40552;
wire n_24499;
wire n_20172;
wire n_43164;
wire n_18421;
wire n_23548;
wire n_9210;
wire newNet_3294;
wire n_15601;
wire n_7539;
wire n_7467;
wire n_13926;
wire sin_out_12;
wire n_38778;
wire n_17746;
wire FE_OCPN1460_n_37232;
wire n_37761;
wire n_7809;
wire n_7218;
wire n_9528;
wire n_18923;
wire newNet_1152;
wire n_12062;
wire n_46195;
wire n_4583;
wire FE_OCPN1512_n_22280;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_30_;
wire n_5603;
wire beta_1;
wire n_2602;
wire n_23267;
wire n_25661;
wire n_13997;
wire n_31321;
wire n_34489;
wire n_41553;
wire n_12257;
wire newNet_2415;
wire newNet_3626;
wire n_26214;
wire n_32591;
wire n_30424;
wire n_21067;
wire newNet_2582;
wire n_7333;
wire n_26004;
wire n_33159;
wire n_18043;
wire n_13332;
wire n_28658;
wire n_41693;
wire n_14915;
wire n_28487;
wire n_24231;
wire FE_OCP_RBN2546_n_44944;
wire n_14648;
wire n_25453;
wire n_42214;
wire newNet_3570;
wire n_24072;
wire n_14378;
wire n_27779;
wire n_34058;
wire n_8376;
wire n_10895;
wire n_16927;
wire n_8051;
wire n_43718;
wire n_26659;
wire n_15876;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_23_;
wire n_46361;
wire n_10733;
wire newNet_2835;
wire FE_RN_207_0;
wire n_20265;
wire n_32204;
wire n_37602;
wire n_4692;
wire n_30402;
wire newNet_1957;
wire n_799;
wire n_5160;
wire n_41003;
wire n_3789;
wire n_38804;
wire n_31177;
wire FE_OCP_RBN1323_n_29056;
wire n_11019;
wire n_13442;
wire n_24302;
wire n_40297;
wire n_27276;
wire newNet_1967;
wire FE_OCP_RBN2143_FE_OCPN861_n_45450;
wire n_21336;
wire n_21324;
wire FE_OCPN1236_n_32791;
wire n_31319;
wire n_32811;
wire n_37152;
wire n_8828;
wire n_14064;
wire newNet_2481;
wire n_19125;
wire n_2120;
wire n_13750;
wire n_36394;
wire n_41056;
wire n_15887;
wire n_29537;
wire FE_OCP_RBN2957_n_26231;
wire n_3252;
wire n_12356;
wire n_35184;
wire n_8836;
wire n_17285;
wire newNet_2868;
wire FE_OCP_RBN2316_n_41420;
wire n_37029;
wire n_36100;
wire n_6207;
wire FE_RN_971_0;
wire n_16690;
wire n_29903;
wire n_17485;
wire n_37812;
wire n_12164;
wire n_35136;
wire n_42857;
wire newNet_3743;
wire n_32191;
wire n_41734;
wire n_26429;
wire n_186;
wire n_22475;
wire n_12286;
wire n_14202;
wire FE_RN_1389_0;
wire n_33664;
wire n_37203;
wire FE_RN_27_0;
wire n_37686;
wire n_10958;
wire n_21376;
wire n_38892;
wire n_15817;
wire n_34685;
wire n_10823;
wire n_3470;
wire n_12922;
wire n_40233;
wire n_3620;
wire n_12881;
wire n_6834;
wire n_16986;
wire n_44066;
wire n_37368;
wire n_36121;
wire n_2426;
wire newNet_2487;
wire n_6363;
wire newNet_513;
wire n_39575;
wire n_845;
wire n_46994;
wire n_34758;
wire n_19646;
wire n_22469;
wire n_2436;
wire n_23956;
wire n_39364;
wire n_9341;
wire n_1858;
wire n_36355;
wire n_21422;
wire newNet_2221;
wire newNet_1246;
wire n_31241;
wire n_6173;
wire n_18860;
wire n_730;
wire n_26890;
wire n_2915;
wire n_11899;
wire n_27401;
wire n_13144;
wire FE_RN_1542_0;
wire n_18084;
wire n_23335;
wire newNet_1076;
wire FE_OFN837_n_4298;
wire n_2270;
wire n_6472;
wire n_43435;
wire n_36005;
wire newNet_1935;
wire n_14985;
wire n_28056;
wire n_37595;
wire n_3822;
wire n_8818;
wire n_20174;
wire newNet_2317;
wire n_9904;
wire FE_RN_802_0;
wire FE_RN_422_0;
wire n_38233;
wire n_9092;
wire FE_RN_1326_0;
wire n_24544;
wire n_7105;
wire n_22793;
wire delay_add_ln22_unr14_stage6_stallmux_q_27_;
wire n_12486;
wire n_17087;
wire n_27438;
wire n_32293;
wire FE_OCP_RBN2380_n_3502;
wire newNet_3427;
wire n_5878;
wire n_41656;
wire FE_OCP_RBN1846_n_22068;
wire n_26645;
wire FE_RN_935_0;
wire n_17070;
wire n_44058;
wire n_21017;
wire n_7141;
wire n_35338;
wire n_25220;
wire n_34359;
wire n_4333;
wire FE_RN_1548_0;
wire FE_OCP_RBN2822_n_10023;
wire n_28118;
wire newNet_1537;
wire n_16305;
wire n_30719;
wire n_22472;
wire newNet_1554;
wire n_17531;
wire n_29698;
wire n_33075;
wire FE_RN_225_0;
wire n_18322;
wire n_21836;
wire n_27327;
wire n_39212;
wire n_12127;
wire FE_OCP_RBN2356_n_13858;
wire n_22056;
wire n_42339;
wire n_15932;
wire n_35768;
wire n_26232;
wire n_26904;
wire n_42976;
wire FE_RN_1153_0;
wire n_9929;
wire n_20631;
wire n_36571;
wire n_10768;
wire n_41956;
wire n_21171;
wire FE_OCP_RBN1919_n_22476;
wire n_32899;
wire n_22421;
wire newNet_2285;
wire n_641;
wire n_18759;
wire n_10644;
wire FE_OCP_RBN1334_n_20249;
wire n_11063;
wire n_9282;
wire n_43828;
wire n_20428;
wire n_5421;
wire n_44623;
wire n_4447;
wire n_22602;
wire n_13319;
wire newNet_3434;
wire n_4788;
wire n_8123;
wire n_22985;
wire n_47175;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_19_;
wire n_18216;
wire n_18195;
wire n_41491;
wire n_9266;
wire n_1999;
wire n_9376;
wire n_83;
wire n_41135;
wire FE_RN_1079_0;
wire n_14412;
wire n_29256;
wire n_33226;
wire n_41646;
wire n_37122;
wire n_20084;
wire n_19844;
wire n_7263;
wire n_9374;
wire n_27855;
wire n_8424;
wire n_30530;
wire n_40740;
wire n_17127;
wire n_10431;
wire n_41725;
wire n_18119;
wire n_8157;
wire n_14724;
wire n_39643;
wire FE_OCP_RBN2184_FE_RN_464_0;
wire n_33613;
wire n_22679;
wire newNet_661;
wire n_22014;
wire n_16602;
wire n_37212;
wire n_2260;
wire n_9961;
wire delay_add_ln22_unr11_stage5_stallmux_q_8_;
wire n_26614;
wire n_7026;
wire n_23404;
wire n_39437;
wire n_17493;
wire n_23044;
wire n_6803;
wire n_18532;
wire n_30148;
wire n_38657;
wire n_43462;
wire n_28743;
wire n_12265;
wire n_32503;
wire n_31853;
wire n_1667;
wire n_16181;
wire n_35645;
wire newNet_2905;
wire n_18901;
wire n_36737;
wire n_14577;
wire n_2689;
wire n_39727;
wire n_33479;
wire n_41674;
wire n_22910;
wire newNet_631;
wire n_15496;
wire n_37801;
wire FE_OCP_RBN3850_n_20290;
wire FE_RN_1313_0;
wire n_8931;
wire n_28134;
wire n_33010;
wire n_38521;
wire n_7684;
wire n_41478;
wire FE_OCP_RBN2650_n_9042;
wire n_16588;
wire n_35770;
wire n_38276;
wire n_42834;
wire n_28541;
wire n_30513;
wire FE_OCPN929_n_44083;
wire n_36826;
wire n_14907;
wire newNet_280;
wire n_6404;
wire n_18123;
wire n_35389;
wire newNet_659;
wire n_17797;
wire n_40519;
wire n_19374;
wire delay_add_ln22_unr2_stage2_stallmux_q_11_;
wire n_6348;
wire FE_OCP_RBN3472_n_7886;
wire n_4944;
wire n_26130;
wire n_40068;
wire n_41296;
wire n_23846;
wire n_7952;
wire n_6181;
wire n_43485;
wire n_34789;
wire n_41676;
wire FE_RN_1746_0;
wire n_20275;
wire n_30005;
wire n_31842;
wire n_17681;
wire n_36899;
wire n_39526;
wire newNet_1657;
wire n_37078;
wire n_8342;
wire n_28195;
wire n_30811;
wire n_3900;
wire n_38793;
wire n_21254;
wire n_9228;
wire n_15056;
wire n_21751;
wire n_32083;
wire n_33784;
wire n_6571;
wire n_3425;
wire n_37728;
wire n_15162;
wire n_4495;
wire n_17358;
wire FE_OCP_RBN3714_n_31466;
wire n_36578;
wire n_14380;
wire n_1563;
wire n_10444;
wire n_34150;
wire n_31697;
wire n_26102;
wire n_38574;
wire n_12238;
wire FE_OCP_RBN1130_n_24179;
wire n_30777;
wire n_14465;
wire n_28512;
wire n_5988;
wire n_40284;
wire FE_OCP_RBN2747_n_9584;
wire FE_OCPN955_n_44460;
wire FE_RN_558_0;
wire n_8443;
wire n_19893;
wire n_36041;
wire n_7884;
wire n_11568;
wire n_40450;
wire n_7962;
wire FE_OCP_RBN3500_n_8187;
wire n_14244;
wire newNet_787;
wire n_35931;
wire FE_OCP_RBN3017_n_31117;
wire n_41154;
wire n_8940;
wire n_30851;
wire n_35927;
wire n_32252;
wire FE_OCP_RBN2549_n_44944;
wire n_17300;
wire n_18649;
wire n_47245;
wire n_14478;
wire n_23061;
wire n_4460;
wire newNet_1509;
wire n_37861;
wire n_7549;
wire n_37196;
wire n_24638;
wire n_39347;
wire n_40013;
wire n_18629;
wire n_40764;
wire FE_RN_470_0;
wire n_32325;
wire n_8530;
wire n_15045;
wire n_19557;
wire n_37891;
wire n_30767;
wire n_30119;
wire n_37403;
wire n_26305;
wire n_5732;
wire n_21644;
wire n_29200;
wire n_12128;
wire newNet_2548;
wire n_840;
wire n_30437;
wire n_306;
wire n_9047;
wire n_41300;
wire n_23810;
wire n_37115;
wire n_32364;
wire FE_RN_561_0;
wire n_35458;
wire n_18835;
wire n_23134;
wire n_38673;
wire newNet_2712;
wire n_788;
wire n_21043;
wire n_5389;
wire n_3759;
wire n_11209;
wire n_14553;
wire n_2744;
wire n_5567;
wire n_26839;
wire n_37624;
wire n_35713;
wire n_839;
wire n_13697;
wire n_9476;
wire FE_OCP_RBN3607_n_8981;
wire n_23046;
wire newNet_156;
wire n_30198;
wire n_23453;
wire n_6188;
wire n_36968;
wire n_19453;
wire n_38329;
wire n_15362;
wire newNet_3369;
wire n_38385;
wire newNet_3382;
wire n_10577;
wire n_4319;
wire n_14632;
wire n_8687;
wire n_31615;
wire n_24701;
wire newNet_1330;
wire n_19202;
wire n_4772;
wire n_14920;
wire n_39058;
wire n_28591;
wire n_37293;
wire n_29112;
wire newNet_477;
wire n_22734;
wire newNet_1314;
wire n_12048;
wire n_40703;
wire n_26816;
wire FE_OCP_RBN2702_n_4041;
wire n_24917;
wire n_33505;
wire n_21157;
wire n_32513;
wire n_41765;
wire n_2301;
wire n_12854;
wire n_46232;
wire n_6665;
wire n_8031;
wire n_38968;
wire n_14301;
wire n_34919;
wire n_38492;
wire n_22342;
wire n_20607;
wire n_3357;
wire n_45503;
wire newNet_1146;
wire n_10088;
wire newNet_3681;
wire n_26509;
wire n_41817;
wire n_17142;
wire n_4969;
wire n_17522;
wire n_3395;
wire FE_OCP_RBN2428_n_8300;
wire FE_OCP_RBN2144_FE_OCPN861_n_45450;
wire n_6733;
wire n_32118;
wire n_41990;
wire n_25098;
wire n_36996;
wire n_28943;
wire n_38012;
wire FE_OCP_RBN3078_FE_OFN807_n_46195;
wire newNet_533;
wire FE_OCP_RBN1204_n_26121;
wire n_8518;
wire n_36629;
wire n_31392;
wire n_46947;
wire n_1609;
wire FE_OFN2_n_43918;
wire n_2742;
wire n_31013;
wire newNet_1846;
wire n_2623;
wire n_11039;
wire n_21894;
wire newNet_3041;
wire n_19056;
wire FE_OCP_RBN2483_n_14326;
wire n_18993;
wire n_14369;
wire n_43595;
wire n_5349;
wire n_8437;
wire n_24017;
wire n_39141;
wire n_41317;
wire n_21492;
wire n_24030;
wire n_20803;
wire n_11153;
wire n_462;
wire n_38660;
wire n_25588;
wire n_24001;
wire n_30215;
wire n_39787;
wire n_6435;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_7_;
wire FE_OCP_RBN2942_n_5454;
wire newNet_3232;
wire newNet_2858;
wire n_4017;
wire n_2826;
wire n_31786;
wire n_414;
wire FE_OCPN986_n_28402;
wire n_4726;
wire newNet_2098;
wire n_15620;
wire n_38959;
wire n_5667;
wire n_31719;
wire n_46253;
wire newNet_2857;
wire n_866;
wire n_5503;
wire FE_RN_1666_0;
wire newNet_386;
wire n_43696;
wire n_34762;
wire n_1631;
wire FE_RN_255_0;
wire n_23713;
wire n_13127;
wire n_19876;
wire n_23004;
wire FE_OCP_RBN3419_n_12739;
wire FE_OCP_RBN2153_n_32772;
wire n_13956;
wire FE_RN_1191_0;
wire n_25533;
wire n_6999;
wire n_26558;
wire FE_OCP_RBN1199_n_25763;
wire n_17789;
wire n_9963;
wire n_33062;
wire n_16385;
wire n_12969;
wire delay_xor_ln22_unr18_stage7_stallmux_q_12_;
wire n_3814;
wire n_9588;
wire n_28406;
wire n_11537;
wire n_2506;
wire n_10276;
wire n_16560;
wire n_20953;
wire FE_OCP_RBN2158_n_1614;
wire n_7452;
wire n_24848;
wire n_35967;
wire n_11755;
wire n_19419;
wire n_34249;
wire n_36260;
wire n_26997;
wire n_5885;
wire n_10423;
wire n_23006;
wire n_43360;
wire n_7376;
wire n_875;
wire n_25728;
wire n_27492;
wire n_1455;
wire newNet_401;
wire n_18286;
wire n_26928;
wire n_41137;
wire newNet_1478;
wire n_17208;
wire newNet_3373;
wire n_37907;
wire n_1829;
wire n_20191;
wire n_34225;
wire n_6510;
wire n_37482;
wire FE_RN_1173_0;
wire n_40041;
wire delay_add_ln22_unr20_stage8_stallmux_q_8_;
wire n_3240;
wire n_7003;
wire n_22456;
wire n_22539;
wire n_17643;
wire n_9387;
wire n_27972;
wire n_6541;
wire n_41972;
wire n_2668;
wire n_1844;
wire n_18668;
wire n_27959;
wire n_34231;
wire n_6938;
wire FE_RN_460_0;
wire n_28252;
wire n_30028;
wire n_30332;
wire n_39108;
wire n_43571;
wire n_21817;
wire n_36231;
wire n_40374;
wire n_19902;
wire n_34985;
wire FE_OCPN3772_n_15371;
wire newNet_1827;
wire n_10986;
wire n_38821;
wire FE_OCP_RBN3535_n_13765;
wire n_36685;
wire FE_RN_235_0;
wire n_12546;
wire n_30164;
wire newNet_1384;
wire n_34707;
wire newNet_858;
wire n_350;
wire n_40573;
wire n_41064;
wire newNet_2698;
wire newNet_2529;
wire n_40309;
wire FE_RN_1615_0;
wire n_33731;
wire n_42575;
wire n_43149;
wire n_19264;
wire newNet_2250;
wire FE_OCP_RBN3479_n_3006;
wire n_20317;
wire n_33530;
wire n_6987;
wire n_6087;
wire n_10927;
wire n_35887;
wire FE_RN_156_0;
wire FE_OCP_RBN2207_n_12907;
wire n_29336;
wire n_8566;
wire n_26497;
wire FE_RN_1058_0;
wire n_9555;
wire sin_out_28;
wire n_6105;
wire newNet_33;
wire newNet_291;
wire n_27159;
wire n_39088;
wire n_34875;
wire n_38912;
wire newNet_1435;
wire n_9742;
wire n_18709;
wire n_27239;
wire n_28961;
wire n_43274;
wire n_26725;
wire n_43870;
wire n_942;
wire n_35242;
wire n_6519;
wire n_34433;
wire n_18712;
wire n_19938;
wire n_1538;
wire n_36315;
wire newNet_3389;
wire n_18374;
wire n_19967;
wire n_15475;
wire n_6064;
wire n_28679;
wire n_25045;
wire n_24139;
wire n_23577;
wire newNet_716;
wire n_11344;
wire n_41103;
wire n_38336;
wire n_2163;
wire n_24579;
wire n_35708;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_15_;
wire n_19639;
wire n_18440;
wire n_25472;
wire n_8053;
wire n_10947;
wire n_38218;
wire n_38239;
wire n_19013;
wire n_6589;
wire n_9567;
wire n_18319;
wire n_28923;
wire n_31079;
wire n_11439;
wire n_42545;
wire n_14612;
wire n_5974;
wire FE_OCPN1779_n_24097;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_24_;
wire n_42413;
wire n_13278;
wire n_36019;
wire n_28067;
wire n_41868;
wire n_2909;
wire n_24202;
wire n_11254;
wire n_27672;
wire n_18345;
wire n_1882;
wire n_18368;
wire FE_OCP_RBN3569_n_9188;
wire n_12116;
wire n_42814;
wire FE_OCP_RBN3426_n_44881;
wire newNet_1238;
wire n_21765;
wire n_11224;
wire n_17609;
wire newNet_3678;
wire n_36338;
wire n_42061;
wire n_22033;
wire n_42090;
wire n_38473;
wire n_903;
wire n_29942;
wire n_36871;
wire n_27810;
wire n_11628;
wire n_37304;
wire n_8077;
wire n_10311;
wire n_33374;
wire n_43688;
wire FE_RN_869_0;
wire n_10462;
wire n_2343;
wire newNet_2629;
wire n_31351;
wire n_42565;
wire newNet_1523;
wire n_17600;
wire n_40539;
wire n_4007;
wire n_35387;
wire n_31107;
wire n_14979;
wire n_23690;
wire newNet_1761;
wire n_32818;
wire n_38270;
wire n_37395;
wire newNet_451;
wire n_21214;
wire n_12438;
wire n_10779;
wire n_1759;
wire n_35344;
wire n_36810;
wire n_29658;
wire n_3332;
wire n_8715;
wire n_24436;
wire newNet_1849;
wire n_35621;
wire FE_RN_978_0;
wire delay_xor_ln23_unr6_stage3_stallmux_q;
wire n_3775;
wire n_32538;
wire n_14685;
wire n_37277;
wire n_8162;
wire FE_OCP_RBN3119_n_22755;
wire n_17192;
wire n_24204;
wire n_868;
wire FE_OCPN3173_n_38799;
wire n_2992;
wire n_13970;
wire delay_add_ln22_unr11_stage5_stallmux_q_6_;
wire n_12745;
wire n_18111;
wire n_38552;
wire n_41134;
wire n_7581;
wire newNet_857;
wire n_38422;
wire n_1047;
wire n_39233;
wire n_4454;
wire n_1062;
wire FE_RN_1260_0;
wire n_23642;
wire n_30626;
wire n_2719;
wire n_21159;
wire n_2889;
wire n_30997;
wire n_27456;
wire n_40161;
wire newNet_1303;
wire n_19224;
wire n_14027;
wire FE_OCP_RBN3408_n_28597;
wire n_2234;
wire n_29741;
wire newNet_2943;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_5_;
wire n_23153;
wire n_35850;
wire n_10981;
wire n_4427;
wire n_7006;
wire n_15503;
wire n_42570;
wire n_33211;
wire n_2217;
wire n_30771;
wire n_7606;
wire FE_RN_827_0;
wire n_41762;
wire n_3257;
wire n_35643;
wire FE_OCP_RBN2212_n_37720;
wire n_22444;
wire n_25785;
wire n_26973;
wire n_32558;
wire n_20195;
wire n_44849;
wire n_16447;
wire n_1271;
wire n_29219;
wire n_41507;
wire FE_RN_400_0;
wire n_5314;
wire n_37432;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_1_;
wire n_35367;
wire n_6349;
wire n_29097;
wire n_42533;
wire n_44850;
wire n_1175;
wire n_1039;
wire n_7117;
wire n_15797;
wire n_3806;
wire n_13356;
wire n_12443;
wire n_2970;
wire n_36300;
wire FE_OCP_RBN2376_n_29480;
wire FE_OCP_RBN3545_n_44575;
wire newNet_5;
wire n_7371;
wire newNet_1430;
wire FE_OFN3_n_43918;
wire n_30894;
wire n_16258;
wire n_35566;
wire n_32263;
wire FE_OCP_RBN3497_n_13818;
wire n_485;
wire n_24090;
wire newNet_2610;
wire n_17200;
wire n_884;
wire delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire n_38183;
wire FE_RN_1681_0;
wire FE_RN_452_0;
wire n_13939;
wire n_6620;
wire FE_OCP_RBN3306_n_44722;
wire FE_RN_334_0;
wire n_14677;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_8_;
wire n_3527;
wire n_21105;
wire FE_OCPN1393_n_962;
wire n_8075;
wire n_38529;
wire n_33172;
wire n_19562;
wire n_42362;
wire newNet_3728;
wire n_16370;
wire n_28977;
wire n_38499;
wire n_10437;
wire FE_OCPN1748_n_23354;
wire n_4257;
wire n_38471;
wire n_33485;
wire newNet_2523;
wire n_25451;
wire n_35369;
wire newNet_293;
wire n_42771;
wire newNet_936;
wire n_35330;
wire n_4963;
wire n_35763;
wire FE_OCP_RBN3488_n_3390;
wire n_624;
wire n_8904;
wire newNet_3627;
wire n_18895;
wire n_11686;
wire newNet_3146;
wire n_29056;
wire n_40254;
wire n_17177;
wire n_45521;
wire n_37484;
wire FE_OCP_RBN2856_n_10176;
wire delay_xor_ln21_unr6_stage3_stallmux_q_3_;
wire n_28967;
wire FE_RN_1546_0;
wire n_15833;
wire n_17380;
wire n_6243;
wire n_11248;
wire n_4826;
wire n_29712;
wire n_31860;
wire FE_OCP_RBN1699_n_19353;
wire n_16550;
wire FE_OCPN1459_n_37232;
wire n_36859;
wire n_7226;
wire n_29507;
wire n_24181;
wire n_35594;
wire n_19973;
wire n_35627;
wire n_8401;
wire n_26826;
wire n_37295;
wire n_42370;
wire n_16617;
wire FE_OCP_RBN3439_n_33803;
wire FE_OCP_RBN2201_n_12808;
wire FE_OCPN886_n_42367;
wire FE_OCP_RBN1353_n_33584;
wire n_9842;
wire n_1871;
wire n_26122;
wire n_13681;
wire n_32274;
wire FE_OCPN1419_n_14003;
wire n_8112;
wire n_37210;
wire n_12830;
wire n_15823;
wire n_23802;
wire n_12543;
wire n_23432;
wire n_19589;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_25_;
wire newNet_3174;
wire n_36995;
wire n_23644;
wire FE_RN_1503_0;
wire n_531;
wire newNet_485;
wire newNet_878;
wire n_30936;
wire n_9337;
wire n_2947;
wire n_11268;
wire newNet_1144;
wire n_23070;
wire n_6730;
wire n_28273;
wire n_36931;
wire FE_OCP_RBN2283_n_33846;
wire n_21064;
wire n_1627;
wire n_13064;
wire n_19957;
wire n_21898;
wire n_16549;
wire n_21526;
wire n_24907;
wire n_43839;
wire newNet_2791;
wire n_41535;
wire n_24660;
wire delay_add_ln22_unr20_stage8_stallmux_q_3_;
wire n_1924;
wire n_12133;
wire n_5226;
wire FE_OCPN917_n_46991;
wire newNet_1598;
wire n_40171;
wire n_13699;
wire n_5563;
wire n_23123;
wire FE_OCP_RBN2171_n_32892;
wire FE_OCPN1455_n_18860;
wire n_20279;
wire newNet_152;
wire FE_OCPN849_n_2306;
wire n_29611;
wire newNet_482;
wire n_13196;
wire n_17263;
wire n_24045;
wire n_33246;
wire n_14951;
wire n_787;
wire n_255;
wire n_4914;
wire FE_RN_347_0;
wire newNet_304;
wire n_25706;
wire n_5132;
wire n_4946;
wire newNet_3181;
wire newNet_3362;
wire n_34600;
wire n_25399;
wire newNet_1068;
wire n_13738;
wire n_38361;
wire FE_OCP_RBN2743_n_15319;
wire FE_RN_986_0;
wire n_14085;
wire FE_RN_1439_0;
wire n_19229;
wire n_35249;
wire n_18370;
wire n_32103;
wire n_40709;
wire n_2054;
wire n_21758;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_7_;
wire delay_xor_ln22_unr21_stage8_stallmux_q_3_;
wire n_9411;
wire n_7717;
wire n_2167;
wire n_26805;
wire n_29242;
wire n_39943;
wire delay_add_ln22_unr27_stage10_stallmux_q_27_;
wire n_2816;
wire n_29786;
wire n_16031;
wire n_38163;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_28_;
wire newNet_96;
wire n_23002;
wire n_21871;
wire n_37975;
wire n_19358;
wire newNet_307;
wire n_4313;
wire n_9634;
wire n_9586;
wire n_27797;
wire n_16343;
wire n_21631;
wire n_23343;
wire n_26448;
wire n_8183;
wire newNet_3705;
wire n_44430;
wire n_19203;
wire n_36285;
wire n_13928;
wire n_9551;
wire n_37846;
wire n_6579;
wire n_31458;
wire n_20430;
wire FE_RN_108_0;
wire n_24938;
wire n_33609;
wire n_33507;
wire n_42223;
wire n_26749;
wire n_5834;
wire n_16676;
wire newNet_1294;
wire n_29681;
wire n_34570;
wire n_36449;
wire n_41128;
wire n_21777;
wire n_18767;
wire n_4505;
wire n_6081;
wire n_21627;
wire n_7138;
wire n_11674;
wire n_11161;
wire n_27386;
wire n_28182;
wire n_17894;
wire delay_xor_ln22_unr18_stage7_stallmux_q_5_;
wire n_18446;
wire FE_OCPN3762_n_34222;
wire FE_OCPN1256_n_13831;
wire FE_OCP_RBN2861_n_10399;
wire n_729;
wire n_12840;
wire n_42547;
wire n_9468;
wire delay_add_ln22_unr11_stage5_stallmux_q_19_;
wire n_23811;
wire newNet_2453;
wire n_5545;
wire n_22009;
wire n_36607;
wire n_17224;
wire n_3979;
wire n_29758;
wire n_41184;
wire n_13510;
wire n_41450;
wire n_2189;
wire newNet_3605;
wire n_27749;
wire n_8474;
wire FE_RN_1468_0;
wire n_1004;
wire FE_RN_198_0;
wire n_14616;
wire newNet_2112;
wire n_41294;
wire n_18137;
wire FE_OCP_RBN2169_n_32892;
wire n_7545;
wire n_32256;
wire n_40778;
wire n_1094;
wire n_30003;
wire n_1901;
wire n_30468;
wire newNet_1998;
wire n_15644;
wire n_40231;
wire n_31733;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_17_;
wire n_18956;
wire n_21576;
wire n_12993;
wire n_1295;
wire n_1488;
wire n_41151;
wire n_31618;
wire n_34286;
wire n_32715;
wire n_22923;
wire n_22568;
wire n_15869;
wire n_27772;
wire n_12715;
wire newNet_3027;
wire n_12449;
wire n_3076;
wire n_29169;
wire n_26086;
wire FE_RN_428_0;
wire n_17559;
wire n_35719;
wire n_24686;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_15_;
wire n_39910;
wire n_32449;
wire n_42486;
wire n_14326;
wire n_3117;
wire n_2071;
wire n_3948;
wire n_7551;
wire n_42216;
wire n_8902;
wire n_29695;
wire n_41623;
wire newNet_712;
wire newNet_2987;
wire n_37156;
wire newNet_249;
wire n_20637;
wire n_35452;
wire n_31148;
wire n_28733;
wire n_10404;
wire n_34833;
wire n_35049;
wire n_41808;
wire n_12727;
wire n_11825;
wire n_22340;
wire n_40338;
wire sin_out_7;
wire n_1713;
wire n_39515;
wire n_15387;
wire FE_RN_1150_0;
wire n_43442;
wire n_42258;
wire n_7827;
wire n_1725;
wire n_5721;
wire FE_OCP_RBN3413_n_12739;
wire n_37406;
wire n_39305;
wire n_28068;
wire n_27081;
wire n_8777;
wire n_4673;
wire n_16798;
wire n_41326;
wire n_7258;
wire newNet_2770;
wire n_38732;
wire n_23447;
wire n_43853;
wire n_13534;
wire n_42003;
wire n_14905;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_5_;
wire newNet_2854;
wire n_25740;
wire n_7980;
wire n_10371;
wire n_35284;
wire n_37194;
wire newNet_2784;
wire n_28925;
wire n_6254;
wire n_35526;
wire FE_RN_1434_0;
wire n_41588;
wire n_27625;
wire FE_RN_1215_0;
wire n_2347;
wire n_39349;
wire n_43106;
wire n_16424;
wire n_42833;
wire n_3426;
wire n_3961;
wire newNet_2574;
wire newNet_1017;
wire FE_OCPN1411_n_21007;
wire n_20884;
wire newNet_2809;
wire n_6842;
wire newNet_1338;
wire n_17641;
wire n_8986;
wire newNet_3385;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_4_;
wire n_30128;
wire FE_OCPN916_n_46991;
wire n_43789;
wire n_14930;
wire n_9430;
wire n_15385;
wire n_41930;
wire n_7109;
wire n_35502;
wire n_2919;
wire n_12506;
wire n_7885;
wire n_17998;
wire newNet_1642;
wire n_23214;
wire n_367;
wire n_15935;
wire n_19465;
wire n_29114;
wire n_34319;
wire n_31644;
wire n_23497;
wire n_1492;
wire FE_OCPN880_n_31944;
wire newNet_1939;
wire n_481;
wire n_19473;
wire n_27423;
wire FE_OCP_RBN2717_n_14982;
wire n_15900;
wire n_40602;
wire n_23605;
wire n_34315;
wire n_27785;
wire newNet_1139;
wire n_1752;
wire n_17725;
wire n_19939;
wire n_31795;
wire n_27153;
wire n_28628;
wire n_7453;
wire n_43548;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_8_;
wire n_3301;
wire n_36657;
wire n_8200;
wire FE_RN_151_0;
wire n_43616;
wire n_46984;
wire n_12635;
wire n_1715;
wire n_41866;
wire delay_add_ln22_unr14_stage6_stallmux_q_25_;
wire n_22587;
wire n_31951;
wire n_31535;
wire n_22508;
wire n_42876;
wire n_4991;
wire n_25081;
wire n_26613;
wire newNet_947;
wire n_26680;
wire n_5166;
wire n_5224;
wire n_10674;
wire n_36336;
wire FE_OCP_RBN3834_n_19241;
wire n_25933;
wire n_46413;
wire newNet_3568;
wire n_29038;
wire n_12122;
wire n_19168;
wire n_42782;
wire n_4784;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_17_;
wire n_8588;
wire n_25545;
wire n_31935;
wire n_37111;
wire n_43529;
wire newNet_333;
wire n_39032;
wire n_9284;
wire newNet_3006;
wire newNet_2715;
wire n_10763;
wire n_21077;
wire n_7458;
wire n_11907;
wire n_36559;
wire n_10001;
wire n_3581;
wire n_23027;
wire n_41050;
wire n_19627;
wire n_41974;
wire n_28265;
wire FE_OCP_RBN2123_n_45224;
wire n_16016;
wire n_28600;
wire n_35597;
wire n_27649;
wire n_45212;
wire n_33971;
wire FE_OCPN961_n_28506;
wire n_23887;
wire n_40544;
wire n_34241;
wire n_40279;
wire n_15248;
wire n_34380;
wire n_309;
wire n_22304;
wire n_13040;
wire FE_OCP_DRV_N1535_n_12633;
wire n_23090;
wire n_14248;
wire newNet_1951;
wire n_11459;
wire n_11310;
wire n_19536;
wire n_6819;
wire n_16028;
wire newNet_45;
wire n_7796;
wire n_19853;
wire n_22080;
wire newNet_633;
wire n_28421;
wire n_29448;
wire newNet_1797;
wire n_18574;
wire n_5468;
wire n_10381;
wire n_31622;
wire FE_OCP_DRV_N1586_n_35594;
wire n_22918;
wire newNet_3417;
wire newNet_2438;
wire n_11638;
wire n_16758;
wire n_21175;
wire n_30376;
wire n_307;
wire n_2272;
wire n_18544;
wire n_43166;
wire newNet_3430;
wire n_24737;
wire n_8544;
wire FE_RN_213_0;
wire delay_xor_ln22_unr9_stage4_stallmux_q_19_;
wire FE_OFN349_n_8981;
wire n_26920;
wire newNet_1035;
wire n_13047;
wire n_5113;
wire n_41909;
wire n_29605;
wire n_24761;
wire n_30326;
wire n_26418;
wire n_42774;
wire FE_RN_985_0;
wire n_33829;
wire n_32000;
wire n_27645;
wire n_22580;
wire newNet_2565;
wire n_4011;
wire n_39770;
wire newNet_3024;
wire newNet_231;
wire n_35289;
wire newNet_2137;
wire n_44511;
wire n_20809;
wire n_34943;
wire n_30026;
wire n_4448;
wire n_3387;
wire n_21891;
wire n_2132;
wire n_4581;
wire n_25717;
wire n_26709;
wire n_19450;
wire n_30807;
wire n_26814;
wire n_16933;
wire n_8366;
wire n_10035;
wire n_31260;
wire newNet_25;
wire n_23898;
wire n_40457;
wire n_43837;
wire n_39459;
wire n_6170;
wire n_43238;
wire n_7300;
wire n_2831;
wire n_11794;
wire n_47013;
wire n_8046;
wire n_8976;
wire n_33835;
wire FE_RN_1811_0;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_18_;
wire n_12219;
wire n_29425;
wire n_9269;
wire n_17472;
wire n_15110;
wire newNet_160;
wire n_20901;
wire n_6119;
wire FE_OCPN1053_n_14098;
wire newNet_2840;
wire newNet_3043;
wire n_2778;
wire n_32790;
wire n_8811;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_0_;
wire n_22018;
wire n_23115;
wire n_37019;
wire FE_OCP_RBN1158_n_18517;
wire n_33729;
wire n_32180;
wire n_42662;
wire FE_OCP_RBN2722_n_4219;
wire newNet_2489;
wire n_7506;
wire n_28935;
wire newNet_2666;
wire n_15566;
wire n_22219;
wire n_34188;
wire n_7210;
wire n_28012;
wire n_19720;
wire n_11245;
wire n_14208;
wire n_37830;
wire n_38322;
wire n_5717;
wire n_4096;
wire n_2664;
wire n_9625;
wire n_1054;
wire n_24977;
wire n_34851;
wire FE_OCP_RBN3271_n_45224;
wire n_38410;
wire n_1675;
wire n_10705;
wire n_20077;
wire n_14655;
wire n_12197;
wire n_46359;
wire n_39310;
wire n_17486;
wire n_8011;
wire FE_OCP_RBN2634_n_30213;
wire n_5600;
wire n_11065;
wire n_30968;
wire n_36973;
wire n_12249;
wire FE_OCP_RBN2959_n_26231;
wire n_30144;
wire newNet_3105;
wire n_35237;
wire n_41738;
wire n_8293;
wire n_22246;
wire n_39567;
wire n_14794;
wire n_6110;
wire n_8055;
wire n_9552;
wire delay_xor_ln22_unr12_stage5_stallmux_q_1_;
wire n_5456;
wire n_18069;
wire n_19645;
wire n_835;
wire delay_xor_ln22_unr6_stage3_stallmux_q_22_;
wire n_5539;
wire n_29494;
wire n_2174;
wire n_43710;
wire n_8151;
wire n_38769;
wire n_33406;
wire n_5340;
wire n_5105;
wire n_20015;
wire n_26015;
wire n_7560;
wire n_38165;
wire n_13001;
wire n_16127;
wire FE_RN_292_0;
wire n_33568;
wire n_29708;
wire newNet_3753;
wire FE_RN_32_0;
wire n_9615;
wire n_8213;
wire n_16008;
wire n_2397;
wire FE_RN_1418_0;
wire n_23685;
wire n_3482;
wire n_17043;
wire n_25823;
wire FE_OCPN948_n_41382;
wire newNet_3460;
wire n_17747;
wire n_22041;
wire n_34582;
wire n_38193;
wire n_739;
wire FE_OCP_RBN3446_n_37945;
wire n_2117;
wire n_41862;
wire n_24249;
wire n_35936;
wire n_36152;
wire n_1136;
wire n_16486;
wire n_26025;
wire n_9523;
wire n_12887;
wire delay_xor_ln22_unr15_stage6_stallmux_q_3_;
wire n_17960;
wire FE_OFN809_n_36594;
wire n_38128;
wire n_18255;
wire n_22463;
wire n_17947;
wire n_32840;
wire n_35447;
wire n_4863;
wire n_4819;
wire n_11936;
wire n_47025;
wire newNet_3123;
wire n_24659;
wire n_42350;
wire n_11016;
wire n_27295;
wire newNet_1914;
wire n_10966;
wire n_30867;
wire n_30453;
wire n_3459;
wire n_34967;
wire newNet_1231;
wire n_25733;
wire n_37820;
wire n_20898;
wire n_43132;
wire newNet_3531;
wire newNet_3323;
wire n_18394;
wire n_35578;
wire FE_RN_1498_0;
wire n_40150;
wire n_6903;
wire n_6952;
wire FE_RN_481_0;
wire n_26799;
wire FE_RN_1269_0;
wire n_16491;
wire newNet_3682;
wire n_34701;
wire n_21259;
wire delay_xor_ln22_unr12_stage5_stallmux_q_2_;
wire n_31869;
wire FE_OCPN860_n_12880;
wire n_27395;
wire n_28475;
wire n_38962;
wire n_12293;
wire n_40288;
wire n_9628;
wire n_44267;
wire delay_add_ln22_unr20_stage8_stallmux_q_14_;
wire n_41748;
wire n_21877;
wire n_6684;
wire FE_RN_221_0;
wire n_28248;
wire FE_OCP_RBN2682_n_35139;
wire n_36484;
wire FE_RN_1426_0;
wire n_26717;
wire newNet_833;
wire n_14157;
wire n_22039;
wire n_26055;
wire n_22372;
wire n_27264;
wire delay_add_ln22_unr11_stage5_stallmux_q_10_;
wire newNet_2725;
wire n_1545;
wire FE_OCPN1038_n_28318;
wire n_27629;
wire n_40054;
wire n_40970;
wire n_33876;
wire n_18586;
wire n_30097;
wire n_2449;
wire n_18183;
wire n_38681;
wire n_41893;
wire n_10081;
wire n_11947;
wire n_39995;
wire n_26871;
wire n_46160;
wire n_31286;
wire n_13646;
wire newNet_3226;
wire n_10067;
wire FE_OCP_RBN2242_n_13017;
wire newNet_3064;
wire n_18239;
wire n_21995;
wire n_4598;
wire n_25692;
wire n_40831;
wire n_12416;
wire newNet_3613;
wire n_15204;
wire n_36831;
wire n_42328;
wire n_42247;
wire n_28367;
wire FE_OCP_RBN1376_n_20889;
wire n_43204;
wire n_25777;
wire FE_OCPN3758_n_2346;
wire n_41454;
wire newNet_508;
wire n_14141;
wire n_36543;
wire n_12215;
wire FE_OCP_RBN2255_n_37844;
wire n_27727;
wire n_40148;
wire n_5277;
wire n_2477;
wire n_13393;
wire n_13895;
wire n_8121;
wire n_23736;
wire n_16310;
wire n_27075;
wire n_795;
wire n_28255;
wire n_30898;
wire newNet_2063;
wire n_6673;
wire n_3465;
wire n_7058;
wire n_39579;
wire n_1461;
wire n_8640;
wire n_21595;
wire FE_RN_1053_0;
wire n_32659;
wire n_43692;
wire n_13452;
wire n_955;
wire n_5148;
wire n_14391;
wire newNet_2752;
wire n_26171;
wire n_16869;
wire n_30881;
wire n_22271;
wire n_39162;
wire FE_RN_680_0;
wire n_2670;
wire n_5883;
wire newNet_1647;
wire cos_out_24;
wire n_35829;
wire n_21216;
wire n_13640;
wire n_8639;
wire n_4220;
wire n_14717;
wire FE_OCP_RBN1925_cordic_combinational_sub_ln23_0_unr12_z_0__;
wire FE_RN_842_0;
wire n_45502;
wire delay_sub_ln22_unr24_stage9_stallmux_q_1_;
wire n_19324;
wire n_7064;
wire n_23910;
wire n_20231;
wire newNet_612;
wire n_14773;
wire newNet_337;
wire FE_RN_812_0;
wire n_38786;
wire n_40425;
wire newNet_2237;
wire n_34545;
wire n_2456;
wire n_11167;
wire n_34182;
wire n_12168;
wire newNet_3738;
wire n_15911;
wire n_29736;
wire n_20170;
wire FE_RN_393_0;
wire n_13922;
wire n_430;
wire n_2629;
wire newNet_802;
wire n_9896;
wire n_27712;
wire n_42471;
wire n_37315;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_18_;
wire n_27966;
wire n_6822;
wire n_26393;
wire n_38300;
wire n_7753;
wire n_47195;
wire n_39503;
wire n_15494;
wire n_42803;
wire n_17795;
wire n_3721;
wire n_13472;
wire n_44829;
wire n_32531;
wire n_37364;
wire FE_RN_1667_0;
wire n_10295;
wire newNet_1379;
wire n_40468;
wire n_2431;
wire n_8160;
wire n_5022;
wire n_17750;
wire newNet_3593;
wire n_11132;
wire n_29474;
wire n_32063;
wire n_10720;
wire n_43456;
wire n_37716;
wire n_4347;
wire n_21387;
wire n_3097;
wire n_37427;
wire n_33131;
wire FE_OCP_RBN2286_n_2433;
wire n_14128;
wire n_14601;
wire n_17291;
wire n_5743;
wire n_43425;
wire n_18633;
wire delay_add_ln22_unr23_stage9_stallmux_q_15_;
wire n_19185;
wire n_25183;
wire n_13012;
wire n_7;
wire n_28098;
wire n_2042;
wire n_26872;
wire n_1633;
wire n_35485;
wire n_5410;
wire n_15721;
wire n_11084;
wire n_4546;
wire n_9082;
wire n_5728;
wire n_33443;
wire n_22720;
wire n_42233;
wire n_11596;
wire n_26833;
wire n_29600;
wire n_46369;
wire newNet_2368;
wire n_29167;
wire n_32823;
wire n_39331;
wire delay_sub_ln23_0_unr25_stage9_stallmux_q;
wire n_15425;
wire n_23475;
wire n_14576;
wire newNet_1755;
wire n_18435;
wire n_43420;
wire n_475;
wire n_7845;
wire FE_OCP_RBN1339_n_32653;
wire newNet_1819;
wire n_15446;
wire n_423;
wire n_43861;
wire n_1395;
wire n_21430;
wire n_17868;
wire n_12096;
wire n_8359;
wire n_45895;
wire n_26098;
wire n_2652;
wire n_15632;
wire n_10814;
wire n_9372;
wire n_13264;
wire FE_RN_49_0;
wire newNet_1156;
wire n_36829;
wire n_22482;
wire n_33267;
wire n_1479;
wire newNet_1633;
wire n_20366;
wire FE_RN_1461_0;
wire n_13082;
wire n_26983;
wire newNet_1349;
wire n_3440;
wire n_10191;
wire n_30692;
wire n_32897;
wire n_40131;
wire n_27092;
wire newNet_1080;
wire n_32833;
wire n_33990;
wire n_17355;
wire n_33497;
wire n_40499;
wire n_33089;
wire n_20985;
wire n_23191;
wire n_194;
wire n_275;
wire newNet_2080;
wire n_16454;
wire n_19172;
wire n_36537;
wire n_16925;
wire n_39905;
wire n_44355;
wire n_43699;
wire FE_OCP_RBN2222_n_13010;
wire newNet_2016;
wire n_26592;
wire n_26756;
wire n_375;
wire FE_RN_629_0;
wire n_30011;
wire n_34782;
wire n_46973;
wire newNet_2519;
wire n_2345;
wire n_31034;
wire FE_OCP_RBN1377_n_20889;
wire FE_OCP_RBN3716_n_39913;
wire n_19010;
wire n_7091;
wire n_23661;
wire newNet_3671;
wire newNet_3285;
wire n_25437;
wire newNet_3012;
wire n_4989;
wire n_34741;
wire n_142;
wire n_36037;
wire n_6582;
wire FE_OCP_RBN1153_n_29053;
wire n_23847;
wire n_40820;
wire n_16141;
wire n_26783;
wire n_10249;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_18_;
wire FE_OCP_RBN2552_n_44921;
wire n_35199;
wire n_1198;
wire n_3874;
wire n_8093;
wire n_38884;
wire newNet_2551;
wire n_25072;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_15_;
wire newNet_2822;
wire n_28454;
wire n_34473;
wire FE_OCPN1854_n_13366;
wire n_22470;
wire n_1250;
wire n_12987;
wire n_27688;
wire FE_OCP_RBN3401_n_37670;
wire n_2424;
wire n_31527;
wire n_36695;
wire n_24369;
wire FE_RN_684_0;
wire n_15669;
wire n_12158;
wire n_22959;
wire delay_add_ln22_unr17_stage7_stallmux_q_14_;
wire n_42113;
wire n_41397;
wire n_36717;
wire n_17588;
wire n_18231;
wire n_18885;
wire n_45332;
wire n_26762;
wire n_30385;
wire n_4953;
wire n_19023;
wire n_260;
wire n_25161;
wire n_20103;
wire n_28745;
wire n_19704;
wire FE_OCP_DRV_N1543_n_18854;
wire newNet_3459;
wire n_15785;
wire n_7291;
wire n_40763;
wire n_35820;
wire n_12349;
wire n_30285;
wire n_27899;
wire n_38820;
wire n_1380;
wire n_35849;
wire FE_OCP_RBN3464_n_7886;
wire n_26384;
wire n_6596;
wire n_25004;
wire n_11346;
wire n_14010;
wire n_25254;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_29_;
wire n_43254;
wire newNet_382;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_2_;
wire n_16785;
wire n_33844;
wire n_35212;
wire newNet_1936;
wire n_747;
wire n_47200;
wire n_4807;
wire n_11843;
wire n_9738;
wire n_16643;
wire n_19525;
wire n_34671;
wire n_27575;
wire n_8371;
wire n_40090;
wire n_9834;
wire n_34561;
wire n_32099;
wire n_19075;
wire n_9880;
wire FE_RN_778_0;
wire n_23460;
wire FE_OCP_RBN3296_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire n_43288;
wire newNet_111;
wire n_31369;
wire n_22715;
wire newNet_104;
wire n_24541;
wire delay_add_ln22_unr23_stage9_stallmux_q_11_;
wire n_38799;
wire n_40721;
wire FE_OFN795_n_45813;
wire n_15021;
wire n_10226;
wire n_16137;
wire n_26620;
wire n_21206;
wire n_20661;
wire n_12093;
wire n_44029;
wire n_45863;
wire n_10897;
wire n_28828;
wire n_15132;
wire n_21677;
wire n_29323;
wire n_13234;
wire n_441;
wire newNet_2052;
wire n_11394;
wire n_14121;
wire n_32783;
wire FE_OCPN1249_n_44267;
wire n_6240;
wire n_22864;
wire n_2195;
wire n_14800;
wire n_16779;
wire n_212;
wire newNet_37;
wire n_21002;
wire n_14870;
wire n_11785;
wire n_11760;
wire n_36425;
wire n_25943;
wire n_3375;
wire n_36773;
wire n_17685;
wire n_6872;
wire n_34726;
wire n_2367;
wire n_38171;
wire n_31676;
wire newNet_3051;
wire n_28382;
wire n_13232;
wire n_37376;
wire n_9493;
wire n_25964;
wire n_33884;
wire newNet_2928;
wire newNet_1308;
wire n_4015;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_16_;
wire FE_OCPN964_n_27287;
wire n_9982;
wire n_39764;
wire n_4075;
wire n_19117;
wire n_20951;
wire n_3350;
wire n_41225;
wire n_19928;
wire newNet_3652;
wire n_39878;
wire n_36110;
wire n_25632;
wire n_23207;
wire n_43174;
wire n_37643;
wire FE_RN_1765_0;
wire n_24699;
wire n_32677;
wire n_18748;
wire newNet_3352;
wire n_43260;
wire n_21314;
wire n_18871;
wire n_8759;
wire n_39639;
wire n_37108;
wire n_34539;
wire n_2278;
wire n_15801;
wire FE_OCP_RBN2843_n_10326;
wire n_2674;
wire n_12408;
wire n_29761;
wire newNet_2284;
wire n_4430;
wire newNet_1382;
wire n_2940;
wire n_32162;
wire n_13833;
wire n_24745;
wire FE_OCP_RBN3356_delay_xor_ln22_unr28_stage10_stallmux_q_0_;
wire n_32548;
wire n_11731;
wire n_17634;
wire n_15985;
wire n_6418;
wire n_28149;
wire n_6279;
wire n_35923;
wire n_6964;
wire n_6679;
wire n_25884;
wire n_8916;
wire n_42985;
wire n_8644;
wire n_17118;
wire n_27954;
wire newNet_1002;
wire n_38110;
wire n_13760;
wire n_33851;
wire n_10095;
wire n_40535;
wire n_3089;
wire n_35188;
wire n_38432;
wire newNet_3139;
wire newNet_1804;
wire n_32132;
wire n_4491;
wire n_16450;
wire n_29827;
wire newNet_189;
wire n_28801;
wire n_38208;
wire n_1766;
wire FE_OCPN1782_FE_OCP_RBN1701_n_19353;
wire n_27051;
wire n_46147;
wire n_29458;
wire newNet_799;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_22_;
wire n_32114;
wire n_32379;
wire n_23383;
wire n_42953;
wire n_30584;
wire n_5976;
wire n_11990;
wire n_43584;
wire newNet_1177;
wire FE_RN_653_0;
wire n_47271;
wire n_6689;
wire n_5500;
wire n_19278;
wire FE_RN_170_0;
wire newNet_3014;
wire n_20531;
wire n_947;
wire n_40470;
wire newNet_1409;
wire n_37619;
wire n_2588;
wire n_13059;
wire n_6288;
wire n_32827;
wire n_38242;
wire n_28558;
wire n_40940;
wire n_19990;
wire FE_RN_62_0;
wire n_25538;
wire n_9444;
wire n_40178;
wire n_26837;
wire FE_OCP_RBN3044_n_46337;
wire n_21603;
wire n_12837;
wire n_3065;
wire FE_RN_1454_0;
wire n_37789;
wire n_19548;
wire n_32273;
wire n_9740;
wire n_42451;
wire n_43597;
wire n_2160;
wire n_27544;
wire n_6627;
wire FE_RN_1420_0;
wire n_39203;
wire n_35546;
wire newNet_2260;
wire n_7641;
wire n_7757;
wire n_22389;
wire n_23595;
wire n_7178;
wire n_13818;
wire n_14770;
wire n_25900;
wire FE_OCPN1020_n_23078;
wire FE_OCP_RBN3719_n_39913;
wire n_9029;
wire n_22333;
wire n_34883;
wire n_36612;
wire n_23398;
wire newNet_1851;
wire n_13821;
wire n_17530;
wire n_20114;
wire FE_OCP_RBN1726_n_20924;
wire n_33242;
wire n_43778;
wire n_39012;
wire n_2105;
wire n_9992;
wire newNet_1901;
wire n_22927;
wire n_43846;
wire n_26679;
wire FE_RN_782_0;
wire newNet_776;
wire newNet_939;
wire n_24283;
wire FE_OCPN1035_n_28288;
wire n_12577;
wire n_15464;
wire n_20862;
wire n_22359;
wire n_3187;
wire n_24443;
wire n_8533;
wire n_40928;
wire n_32804;
wire n_935;
wire n_45145;
wire FE_OCP_RBN3218_n_21358;
wire newNet_2536;
wire FE_OFN766_n_15670;
wire n_43683;
wire n_46347;
wire n_20184;
wire n_13779;
wire n_33594;
wire FE_OCP_RBN2378_n_29480;
wire n_25371;
wire n_35497;
wire FE_RN_769_0;
wire newNet_1123;
wire n_18199;
wire newNet_864;
wire n_17182;
wire n_29845;
wire n_17212;
wire n_20736;
wire newNet_3420;
wire n_878;
wire beta_9;
wire n_36058;
wire n_35688;
wire n_4853;
wire n_27003;
wire n_28918;
wire n_31469;
wire n_9866;
wire n_28539;
wire n_30310;
wire n_40981;
wire FE_OCP_RBN3712_n_31466;
wire n_6374;
wire n_22179;
wire n_12401;
wire n_22044;
wire n_5476;
wire n_37118;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_4_;
wire n_12515;
wire n_33812;
wire n_8590;
wire n_28039;
wire n_2124;
wire n_24912;
wire n_37217;
wire n_1448;
wire n_32309;
wire n_27227;
wire n_31127;
wire n_25002;
wire newNet_3164;
wire n_42196;
wire n_12017;
wire FE_RN_340_0;
wire newNet_2652;
wire n_44761;
wire n_43883;
wire FE_OCP_RBN1678_n_44847;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_11_;
wire n_21725;
wire n_412;
wire newNet_1557;
wire FE_OCP_RBN2156_n_1602;
wire n_6947;
wire n_15469;
wire n_18894;
wire newNet_1664;
wire n_17615;
wire FE_RN_1015_0;
wire n_2238;
wire n_9874;
wire n_15881;
wire n_43345;
wire n_36593;
wire n_490;
wire n_19215;
wire n_20474;
wire n_25714;
wire n_17739;
wire n_34009;
wire n_38214;
wire n_27851;
wire n_1264;
wire n_12101;
wire n_33068;
wire n_18327;
wire n_28294;
wire n_26107;
wire newNet_2860;
wire n_33782;
wire n_14965;
wire n_41879;
wire n_38197;
wire n_354;
wire newNet_3159;
wire n_18337;
wire FE_OCP_RBN3565_n_29857;
wire n_37091;
wire FE_OCP_RBN2913_n_30949;
wire n_37231;
wire n_21887;
wire n_43065;
wire n_14652;
wire n_34776;
wire n_1038;
wire n_16253;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_9_;
wire n_39983;
wire n_8998;
wire n_3646;
wire n_12034;
wire n_23560;
wire n_26329;
wire newNet_1981;
wire n_13482;
wire n_36630;
wire n_34634;
wire n_25626;
wire n_17277;
wire n_24900;
wire n_20289;
wire n_15927;
wire n_35425;
wire n_26724;
wire newNet_322;
wire n_3410;
wire n_322;
wire n_41948;
wire n_18498;
wire n_5129;
wire n_40366;
wire n_37637;
wire n_32631;
wire newNet_1370;
wire newNet_3117;
wire n_20012;
wire n_29749;
wire n_25116;
wire n_10031;
wire n_11684;
wire n_2905;
wire n_22338;
wire n_43639;
wire newNet_1465;
wire n_7665;
wire n_13316;
wire n_18613;
wire n_36040;
wire n_18467;
wire n_15059;
wire n_36122;
wire n_10787;
wire n_6747;
wire n_22828;
wire n_1235;
wire n_31422;
wire n_18096;
wire FE_OFN834_n_2285;
wire newNet_3244;
wire n_2897;
wire n_42063;
wire n_14681;
wire n_31540;
wire n_38034;
wire n_21616;
wire n_36490;
wire n_34032;
wire n_32755;
wire n_6992;
wire n_29655;
wire n_40513;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_10_;
wire n_32300;
wire n_40582;
wire n_11124;
wire FE_OCPN1524_n_45072;
wire n_14869;
wire n_28652;
wire n_17317;
wire n_18075;
wire FE_OCP_RBN2642_n_34921;
wire FE_OCP_RBN3621_n_15135;
wire n_41076;
wire n_6210;
wire n_41172;
wire n_39737;
wire n_2213;
wire n_8972;
wire n_26790;
wire n_22992;
wire newNet_2431;
wire FE_RN_60_0;
wire n_20332;
wire n_969;
wire n_22857;
wire n_7131;
wire n_44441;
wire n_4515;
wire n_1863;
wire newNet_1098;
wire n_13224;
wire n_28076;
wire n_36912;
wire n_27207;
wire n_27345;
wire n_35403;
wire n_10222;
wire n_26007;
wire FE_RN_1512_0;
wire n_7631;
wire n_42464;
wire n_357;
wire n_38616;
wire n_25594;
wire n_42010;
wire n_17965;
wire n_39852;
wire newNet_601;
wire n_33222;
wire n_35810;
wire n_14291;
wire n_46938;
wire n_14998;
wire n_22416;
wire n_23689;
wire n_5787;
wire FE_OCPN908_n_23227;
wire n_5056;
wire n_13493;
wire n_28793;
wire n_14070;
wire n_776;
wire n_39953;
wire newNet_657;
wire n_439;
wire n_36566;
wire n_15553;
wire n_1671;
wire n_2332;
wire n_40249;
wire n_16436;
wire n_18080;
wire n_15241;
wire FE_OCPN1753_n_7225;
wire n_44624;
wire n_10036;
wire n_3919;
wire n_38909;
wire n_5697;
wire n_27719;
wire n_25882;
wire n_34802;
wire n_18822;
wire n_33926;
wire FE_RN_444_0;
wire n_10759;
wire n_589;
wire n_4234;
wire n_12796;
wire n_18578;
wire n_8320;
wire n_29254;
wire n_37548;
wire n_25868;
wire n_36169;
wire n_2019;
wire n_30646;
wire newNet_1030;
wire newNet_13;
wire n_16359;
wire n_11975;
wire delay_add_ln22_unr17_stage7_stallmux_q_7_;
wire n_11753;
wire n_45824;
wire newNet_2951;
wire n_9704;
wire n_45899;
wire n_44055;
wire FE_RN_721_0;
wire n_9062;
wire n_31954;
wire n_31667;
wire n_23507;
wire FE_RN_1545_0;
wire n_14098;
wire newNet_219;
wire n_7037;
wire newNet_1932;
wire n_22425;
wire n_26759;
wire n_22391;
wire n_11314;
wire FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_28779;
wire n_20058;
wire n_15676;
wire n_3192;
wire newNet_3669;
wire n_24869;
wire newNet_3486;
wire n_10592;
wire n_16244;
wire n_18404;
wire n_43392;
wire n_1112;
wire n_11870;
wire delay_xor_ln22_unr9_stage4_stallmux_q_16_;
wire n_41823;
wire newNet_954;
wire newNet_724;
wire n_35736;
wire n_22742;
wire n_7418;
wire n_18350;
wire n_38763;
wire FE_OCP_RBN1364_n_20412;
wire n_21164;
wire n_19596;
wire n_35461;
wire n_2178;
wire n_32376;
wire newNet_2205;
wire n_26135;
wire n_3718;
wire n_25819;
wire n_27413;
wire n_38399;
wire n_33022;
wire n_28340;
wire FE_OCP_RBN2755_n_30558;
wire newNet_2419;
wire n_15077;
wire n_20689;
wire n_31876;
wire n_20920;
wire n_32976;
wire FE_RN_95_0;
wire n_29479;
wire FE_RN_399_0;
wire n_47187;
wire n_5093;
wire n_3107;
wire n_4130;
wire newNet_2641;
wire n_31030;
wire n_37244;
wire n_38568;
wire newNet_146;
wire tau_clk;
wire n_41635;
wire n_2282;
wire n_21269;
wire n_10008;
wire FE_OCP_RBN1214_n_31847;
wire n_35489;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_5_;
wire n_3662;
wire n_21902;
wire delay_add_ln22_unr2_stage2_stallmux_q_25_;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_28_;
wire n_32602;
wire newNet_2273;
wire FE_RN_551_0;
wire n_47248;
wire n_26689;
wire n_2607;
wire n_15749;
wire n_973;
wire n_19923;
wire n_29621;
wire FE_RN_537_0;
wire n_21705;
wire n_37341;
wire n_29704;
wire n_17648;
wire n_43632;
wire n_41643;
wire n_5031;
wire n_29874;
wire n_1072;
wire n_9556;
wire n_16667;
wire n_22127;
wire FE_RN_1734_0;
wire n_39900;
wire newNet_579;
wire n_24969;
wire n_43082;
wire n_32646;
wire FE_RN_1596_0;
wire delay_add_ln22_unr11_stage5_stallmux_q_15_;
wire n_42239;
wire n_10218;
wire n_39321;
wire n_7594;
wire n_1807;
wire n_25773;
wire FE_OCP_RBN2689_n_38870;
wire n_34421;
wire n_31573;
wire n_8840;
wire n_11605;
wire n_8232;
wire n_5065;
wire FE_OCP_RBN1131_n_24179;
wire n_18980;
wire n_30197;
wire n_25642;
wire FE_OCPN1394_n_962;
wire n_34139;
wire n_32346;
wire newNet_2349;
wire n_32722;
wire n_11367;
wire FE_RN_1775_0;
wire n_2885;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_20_;
wire n_39492;
wire FE_RN_1705_0;
wire FE_RN_601_0;
wire n_1972;
wire n_20508;
wire n_458;
wire n_35717;
wire FE_OCPN1241_n_7721;
wire n_8230;
wire n_13782;
wire n_43481;
wire n_21572;
wire newNet_1325;
wire n_40079;
wire n_21480;
wire n_35827;
wire FE_OCP_RBN2393_n_8288;
wire n_23038;
wire newNet_2931;
wire n_30673;
wire n_3986;
wire n_31741;
wire newNet_741;
wire n_10168;
wire n_41897;
wire n_35480;
wire n_43460;
wire n_379;
wire n_44823;
wire newNet_132;
wire n_6729;
wire n_7088;
wire n_27796;
wire n_44420;
wire newNet_1729;
wire n_25505;
wire delay_add_ln22_unr14_stage6_stallmux_q_23_;
wire n_752;
wire n_37778;
wire n_43746;
wire n_33048;
wire n_41031;
wire n_17322;
wire n_40617;
wire n_15195;
wire n_27506;
wire n_29799;
wire n_31836;
wire n_41358;
wire n_39603;
wire n_15538;
wire n_7894;
wire n_26221;
wire n_3505;
wire n_18511;
wire n_23361;
wire n_5320;
wire n_34573;
wire n_21923;
wire n_7060;
wire n_3725;
wire FE_OCP_RBN3063_n_11325;
wire n_33623;
wire n_34153;
wire FE_OCP_RBN2895_n_39575;
wire n_30170;
wire newNet_1643;
wire n_81;
wire n_5559;
wire n_25574;
wire n_33524;
wire n_28286;
wire n_27751;
wire delay_xor_ln22_unr15_stage6_stallmux_q_14_;
wire n_12130;
wire newNet_2507;
wire n_7573;
wire n_41782;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_24_;
wire n_15512;
wire n_26713;
wire n_14057;
wire n_32221;
wire n_38050;
wire n_41548;
wire n_22768;
wire n_22481;
wire n_3720;
wire n_28527;
wire newNet_2798;
wire n_40560;
wire n_13025;
wire n_10470;
wire newNet_2394;
wire newNet_889;
wire FE_RN_143_0;
wire n_23657;
wire n_5809;
wire n_18624;
wire n_45204;
wire n_36252;
wire n_46184;
wire n_29388;
wire n_37983;
wire n_34415;
wire n_5513;
wire n_19328;
wire n_4088;
wire newNet_2777;
wire n_40637;
wire n_29170;
wire n_46164;
wire n_30763;
wire n_31001;
wire FE_RN_745_0;
wire n_16296;
wire n_15374;
wire n_19745;
wire n_25749;
wire n_46227;
wire FE_OCP_DRV_N1558_n_19590;
wire n_26511;
wire n_19161;
wire FE_RN_1401_0;
wire n_3672;
wire n_32606;
wire n_10354;
wire n_27520;
wire n_960;
wire n_37069;
wire n_25686;
wire n_7470;
wire n_12608;
wire n_39357;
wire newNet_1765;
wire n_27323;
wire delay_add_ln22_unr23_stage9_stallmux_q_26_;
wire n_15293;
wire n_34746;
wire n_42895;
wire n_38267;
wire n_29553;
wire n_45741;
wire FE_RN_1399_0;
wire newNet_2326;
wire n_37171;
wire n_43478;
wire n_37497;
wire newNet_2192;
wire FE_RN_752_0;
wire n_29782;
wire n_30051;
wire n_32589;
wire delay_xor_ln21_unr3_stage2_stallmux_q_21_;
wire n_3578;
wire n_35448;
wire newNet_529;
wire n_2244;
wire n_6128;
wire n_19462;
wire n_18225;
wire n_30520;
wire n_40141;
wire n_20759;
wire n_3299;
wire n_22319;
wire n_37148;
wire n_28320;
wire n_41405;
wire n_14274;
wire n_21749;
wire n_7077;
wire n_7972;
wire n_29641;
wire n_21272;
wire n_16052;
wire n_30988;
wire n_40932;
wire n_7732;
wire n_16498;
wire n_1529;
wire n_13175;
wire n_27088;
wire n_11435;
wire n_9308;
wire n_14152;
wire n_37842;
wire n_42129;
wire n_39674;
wire n_42335;
wire n_2330;
wire n_30090;
wire newNet_2044;
wire newNet_702;
wire newNet_951;
wire n_26434;
wire n_42268;
wire n_34640;
wire newNet_1078;
wire n_7325;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_22_;
wire newNet_2676;
wire n_37419;
wire n_40441;
wire n_27781;
wire n_46175;
wire n_22821;
wire n_12524;
wire newNet_3508;
wire n_31770;
wire newNet_2818;
wire delay_xor_ln21_unr9_stage4_stallmux_q_1_;
wire n_13706;
wire n_40502;
wire n_20690;
wire n_33105;
wire newNet_2769;
wire FE_RN_977_0;
wire n_36665;
wire n_2470;
wire n_13199;
wire delay_add_ln22_unr8_stage4_stallmux_q_16_;
wire n_5201;
wire n_38974;
wire n_15319;
wire n_9108;
wire n_20354;
wire n_46217;
wire n_14193;
wire n_31214;
wire newNet_2971;
wire n_18178;
wire n_32693;
wire n_21953;
wire n_11045;
wire n_17092;
wire n_22835;
wire n_14740;
wire n_10375;
wire n_24494;
wire newNet_1140;
wire n_22317;
wire n_24417;
wire n_19882;
wire n_23586;
wire n_28234;
wire n_3014;
wire n_14837;
wire n_7347;
wire n_25968;
wire FE_OCP_RBN2678_n_9247;
wire n_4653;
wire n_30799;
wire n_1875;
wire n_23019;
wire newNet_370;
wire n_33398;
wire n_19833;
wire n_41096;
wire n_16505;
wire n_17455;
wire n_23276;
wire FE_OCP_RBN2719_n_9182;
wire n_10799;
wire n_40007;
wire n_35260;
wire n_12386;
wire FE_RN_1343_0;
wire newNet_56;
wire n_13243;
wire n_38467;
wire n_29233;
wire n_6168;
wire newNet_3196;
wire newNet_3101;
wire newNet_803;
wire n_1337;
wire n_43243;
wire n_26589;
wire n_19456;
wire n_38587;
wire n_28998;
wire FE_OCP_RBN3559_n_8809;
wire n_12313;
wire newNet_974;
wire n_33533;
wire n_39753;
wire newNet_1244;
wire n_28639;
wire n_43359;
wire n_43557;
wire n_34054;
wire n_2493;
wire FE_OCP_RBN2386_n_8342;
wire n_13180;
wire n_29669;
wire n_3337;
wire n_33763;
wire newNet_1884;
wire n_32791;
wire n_16362;
wire n_6159;
wire n_30545;
wire n_5930;
wire n_27014;
wire n_34856;
wire n_7918;
wire n_31207;
wire beta_6;
wire n_8910;
wire n_38084;
wire n_23576;
wire n_6766;
wire n_20314;
wire n_2340;
wire n_7187;
wire FE_RN_490_0;
wire n_6892;
wire FE_OCPN999_n_19311;
wire n_10741;
wire n_27595;
wire n_310;
wire n_32237;
wire n_41259;
wire n_15088;
wire n_221;
wire n_26237;
wire n_44869;
wire n_14210;
wire n_20708;
wire n_25351;
wire n_36763;
wire n_2156;
wire n_26693;
wire newNet_3445;
wire newNet_3089;
wire n_38624;
wire n_9346;
wire n_3363;
wire n_24424;
wire n_22542;
wire FE_RN_1856_0;
wire n_2599;
wire n_28873;
wire n_7241;
wire delay_add_ln22_unr27_stage10_stallmux_q_22_;
wire FE_OCP_RBN2486_n_3498;
wire n_714;
wire n_32652;
wire newNet_3110;
wire n_40849;
wire n_17704;
wire delay_xor_ln22_unr6_stage3_stallmux_q_3_;
wire n_23242;
wire n_43152;
wire n_34484;
wire n_39126;
wire n_20974;
wire n_24839;
wire n_38079;
wire newNet_2428;
wire n_11374;
wire n_46247;
wire FE_RN_578_0;
wire n_38419;
wire n_3043;
wire n_2570;
wire n_11818;
wire n_18966;
wire n_14782;
wire newNet_2743;
wire n_1000;
wire n_27738;
wire FE_RN_1094_0;
wire n_38696;
wire sin_out_24;
wire n_2519;
wire n_28448;
wire n_1014;
wire n_32469;
wire n_21453;
wire n_5192;
wire n_36098;
wire FE_OCPN1485_n_27315;
wire n_8770;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_30_;
wire n_13942;
wire n_29462;
wire n_6961;
wire n_31183;
wire n_5537;
wire n_37354;
wire n_8649;
wire n_29549;
wire FE_OCPN869_n_16086;
wire n_6518;
wire n_23852;
wire n_4757;
wire n_32978;
wire n_45135;
wire n_9351;
wire FE_OFN49_n_1045;
wire n_39039;
wire n_7907;
wire n_32894;
wire newNet_3543;
wire n_12454;
wire n_10179;
wire n_23534;
wire FE_RN_803_0;
wire FE_OCP_RBN3613_n_20249;
wire n_2085;
wire n_33901;
wire n_32427;
wire n_12067;
wire n_45813;
wire n_7709;
wire n_9570;
wire n_13616;
wire newNet_2978;
wire n_5581;
wire n_45871;
wire n_10806;
wire n_2702;
wire n_23536;
wire delay_xor_ln22_unr3_stage2_stallmux_q_0_;
wire n_32814;
wire n_38020;
wire n_21961;
wire n_43714;
wire n_17248;
wire n_32190;
wire n_14730;
wire n_41842;
wire n_24980;
wire n_169;
wire n_688;
wire n_19017;
wire n_36520;
wire n_8270;
wire FE_OFN827_n_1941;
wire n_25488;
wire n_42179;
wire n_31805;
wire FE_OFN220_n_35655;
wire FE_OCP_RBN2046_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire n_8737;
wire n_38008;
wire n_25262;
wire n_39860;
wire n_11424;
wire n_42585;
wire n_38580;
wire n_3891;
wire n_16936;
wire n_32775;
wire FE_RN_1457_0;
wire newNet_421;
wire newNet_345;
wire n_34120;
wire n_35913;
wire n_21471;
wire n_35269;
wire n_1932;
wire n_7144;
wire n_12452;
wire n_33037;
wire n_28485;
wire newNet_3216;
wire newNet_2376;
wire n_2841;
wire n_17622;
wire n_36691;
wire n_37128;
wire newNet_338;
wire n_14206;
wire n_5907;
wire n_13653;
wire n_25166;
wire FE_OCPN1474_n_24624;
wire FE_OCPN1467_n_12968;
wire newNet_2216;
wire n_7647;
wire n_21540;
wire n_34827;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_1_;
wire n_44812;
wire n_41686;
wire n_19673;
wire n_46354;
wire n_42295;
wire n_3403;
wire n_20327;
wire n_19624;
wire FE_RN_728_0;
wire n_19846;
wire n_19981;
wire FE_RN_1100_0;
wire n_22439;
wire FE_RN_1850_0;
wire n_43765;
wire n_29587;
wire n_28021;
wire n_30652;
wire n_23959;
wire n_37266;
wire n_21283;
wire n_36877;
wire n_29393;
wire n_26251;
wire FE_OCP_DRV_N3151_n_13264;
wire n_36478;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_23_;
wire n_1755;
wire newNet_2999;
wire n_7307;
wire n_32749;
wire n_14007;
wire n_46990;
wire n_24237;
wire n_31484;
wire n_30151;
wire n_40379;
wire n_7427;
wire n_6855;
wire n_32864;
wire n_4537;
wire n_7728;
wire n_35139;
wire n_1744;
wire n_17354;
wire n_44453;
wire delay_xor_ln22_unr12_stage5_stallmux_q_9_;
wire n_3858;
wire n_7862;
wire n_15454;
wire newNet_1875;
wire n_8951;
wire n_46154;
wire n_42554;
wire n_3847;
wire n_34917;
wire newNet_564;
wire n_10410;
wire n_33892;
wire n_37273;
wire newNet_489;
wire n_35611;
wire FE_RN_1590_0;
wire n_6547;
wire n_16024;
wire n_37189;
wire n_37691;
wire n_4874;
wire newNet_1519;
wire newNet_2994;
wire n_33000;
wire n_46342;
wire n_8584;
wire n_38798;
wire delay_xor_ln22_unr9_stage4_stallmux_q_8_;
wire n_43773;
wire n_28175;
wire n_3557;
wire n_25461;
wire newNet_2383;
wire n_36464;
wire n_12689;
wire n_32470;
wire n_4450;
wire n_43918;
wire FE_RN_1061_0;
wire n_38426;
wire n_10818;
wire n_30185;
wire n_2372;
wire n_8063;
wire FE_OCPN1233_n_2414;
wire n_15406;
wire n_35562;
wire newNet_1206;
wire n_38629;
wire n_10636;
wire FE_RN_376_0;
wire FE_RN_1790_0;
wire newNet_2703;
wire newNet_1947;
wire n_9925;
wire n_1324;
wire n_8142;
wire n_16705;
wire FE_RN_1385_0;
wire n_34778;
wire n_293;
wire n_17929;
wire n_33341;
wire delay_xor_ln21_unr18_stage7_stallmux_q_11_;
wire n_5875;
wire n_28491;
wire n_24887;
wire FE_RN_702_0;
wire n_9937;
wire n_32259;
wire n_12161;
wire n_31195;
wire n_13162;
wire n_32354;
wire n_11798;
wire n_36136;
wire n_40083;
wire n_27790;
wire n_30534;
wire FE_OCP_RBN3286_n_44365;
wire n_22907;
wire n_7806;
wire n_40349;
wire n_46942;
wire n_1248;
wire n_14761;
wire n_28501;
wire newNet_3338;
wire n_39028;
wire newNet_1978;
wire n_40118;
wire delay_xor_ln21_unr9_stage4_stallmux_q_19_;
wire n_39975;
wire n_10919;
wire n_18693;
wire n_23602;
wire n_41792;
wire n_33772;
wire newNet_1057;
wire n_13950;
wire n_19405;
wire n_30389;
wire newNet_2038;
wire n_31586;
wire newNet_1343;
wire n_32669;
wire newNet_1674;
wire n_42764;
wire n_20078;
wire n_43213;
wire n_42204;
wire n_8708;
wire n_37738;
wire n_454;
wire n_267;
wire n_41144;
wire n_43364;
wire n_30225;
wire FE_OCP_RBN2789_n_4294;
wire n_34321;
wire FE_OCP_RBN1343_n_19077;
wire n_8209;
wire n_28821;
wire n_12151;
wire n_6005;
wire FE_RN_1039_0;
wire n_42408;
wire n_38525;
wire n_39065;
wire n_40165;
wire n_26850;
wire n_9290;
wire n_5888;
wire n_22020;
wire n_42082;
wire newNet_262;
wire n_30419;
wire delay_add_ln22_unr20_stage8_stallmux_q_5_;
wire n_47006;
wire n_36326;
wire FE_OCP_RBN2867_n_16088;
wire n_39384;
wire newNet_1362;
wire FE_OCP_RBN2752_n_15461;
wire n_31949;
wire n_28746;
wire FE_OCP_RBN3039_n_46337;
wire n_19977;
wire n_34443;
wire n_41770;
wire n_40357;
wire n_27145;
wire n_27304;
wire n_19332;
wire newNet_81;
wire n_26126;
wire n_16760;
wire n_30086;
wire n_37920;
wire n_37895;
wire n_19519;
wire FE_RN_743_0;
wire newNet_3471;
wire n_40901;
wire n_987;
wire n_18688;
wire n_3693;
wire n_6062;
wire n_13019;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_2_;
wire n_6368;
wire n_23145;
wire n_32989;
wire n_9390;
wire n_41347;
wire n_18815;
wire FE_RN_2_0;
wire FE_RN_204_0;
wire n_26901;
wire n_31210;
wire n_37420;
wire FE_RN_22_0;
wire n_11273;
wire n_46250;
wire newNet_3450;
wire n_8478;
wire n_1792;
wire n_9046;
wire n_39685;
wire n_10611;
wire FE_RN_1201_0;
wire n_30956;
wire n_7995;
wire n_30845;
wire n_21406;
wire FE_OCP_RBN3029_n_39942;
wire n_7988;
wire n_42940;
wire newNet_2795;
wire n_39299;
wire n_13152;
wire n_9485;
wire n_16898;
wire n_39396;
wire n_27110;
wire n_18134;
wire n_20836;
wire n_26217;
wire n_134;
wire n_26572;
wire n_12996;
wire n_20412;
wire FE_RN_699_0;
wire n_36595;
wire n_37567;
wire n_40430;
wire n_33639;
wire n_3051;
wire newNet_1476;
wire n_41531;
wire n_4666;
wire n_2405;
wire n_36186;
wire newNet_44;
wire n_28721;
wire n_20046;
wire newNet_932;
wire newNet_2357;
wire n_16177;
wire newNet_584;
wire FE_RN_186_0;
wire n_42977;
wire n_41116;
wire n_24087;
wire newNet_2627;
wire n_13099;
wire n_32459;
wire n_37080;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_4_;
wire n_40314;
wire n_12629;
wire n_12904;
wire n_35258;
wire n_24561;
wire n_39871;
wire newNet_1808;
wire n_43603;
wire n_13204;
wire n_8496;
wire n_34492;
wire n_43825;
wire n_24514;
wire n_8187;
wire FE_RN_327_0;
wire FE_OCP_RBN2878_n_15553;
wire n_31614;
wire FE_RN_1181_0;
wire n_36726;
wire n_7315;
wire n_9811;
wire n_9053;
wire FE_RN_1291_0;
wire n_12076;
wire n_27872;
wire n_3416;
wire n_36413;
wire n_32714;
wire n_27539;
wire n_19606;
wire newNet_2241;
wire FE_OCP_RBN1328_n_36489;
wire FE_OCP_RBN1178_n_18981;
wire n_29301;
wire newNet_2600;
wire n_25909;
wire n_46363;
wire n_6313;
wire n_21395;
wire n_42706;
wire FE_RN_1226_0;
wire n_17225;
wire FE_RN_1466_0;
wire n_16900;
wire n_43208;
wire n_10656;
wire n_40591;
wire n_15041;
wire n_12652;
wire n_16849;
wire newNet_2124;
wire n_4611;
wire n_33868;
wire FE_OCP_RBN2615_n_35005;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_3_;
wire n_18915;
wire n_2389;
wire n_42166;
wire n_16555;
wire FE_OCP_DRV_N1546_n_18860;
wire n_20977;
wire n_30852;
wire n_8599;
wire n_43612;
wire n_29583;
wire n_33562;
wire n_33015;
wire newNet_1740;
wire n_32407;
wire n_36316;
wire n_18609;
wire n_10708;
wire FE_OCPN1773_n_30210;
wire n_43465;
wire n_36247;
wire n_34816;
wire n_22765;
wire n_17657;
wire n_26732;
wire n_32226;
wire delay_xor_ln21_unr6_stage3_stallmux_q_15_;
wire n_25444;
wire FE_OFN1_n_43918;
wire newNet_2060;
wire FE_OCP_RBN1189_n_14911;
wire n_36059;
wire n_39750;
wire n_8869;
wire n_16950;
wire n_274;
wire FE_RN_1836_0;
wire newNet_780;
wire newNet_575;
wire n_13007;
wire newNet_353;
wire newNet_2334;
wire n_1617;
wire n_5792;
wire n_24392;
wire FE_OCP_RBN3007_n_31117;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_17_;
wire newNet_3709;
wire n_21306;
wire delay_add_ln22_unr23_stage9_stallmux_q_13_;
wire n_736;
wire beta_2;
wire n_26336;
wire n_28148;
wire n_34000;
wire n_40750;
wire n_43144;
wire n_1586;
wire n_33862;
wire FE_OCP_RBN2257_n_37844;
wire n_36952;
wire n_47176;
wire FE_RN_1509_0;
wire n_7768;
wire n_13253;
wire n_19154;
wire n_19905;
wire n_41321;
wire n_19284;
wire n_2830;
wire newNet_99;
wire n_165;
wire n_23955;
wire FE_RN_1696_0;
wire n_41660;
wire n_22795;
wire n_24350;
wire n_20612;
wire n_3754;
wire n_30836;
wire n_39552;
wire n_26671;
wire n_363;
wire n_19439;
wire n_32153;
wire n_36082;
wire n_31123;
wire n_29375;
wire n_25820;
wire FE_OCPN1862_n_30319;
wire n_34450;
wire n_17592;
wire n_147;
wire n_17169;
wire newNet_2138;
wire n_28025;
wire n_41187;
wire n_31980;
wire n_30931;
wire n_1197;
wire n_41108;
wire newNet_1255;
wire n_32912;
wire delay_add_ln22_unr17_stage7_stallmux_q_15_;
wire n_28121;
wire newNet_594;
wire n_36299;
wire delay_xor_ln22_unr15_stage6_stallmux_q_13_;
wire n_42993;
wire n_1432;
wire n_29433;
wire n_12618;
wire n_9361;
wire n_14349;
wire n_19732;
wire n_9748;
wire n_31843;
wire n_349;
wire n_42060;
wire n_40069;
wire n_30610;
wire n_13981;
wire n_40958;
wire n_10488;
wire n_42097;
wire n_39687;
wire n_16817;
wire n_39525;
wire n_14706;
wire n_46966;
wire n_16838;
wire n_18939;
wire FE_RN_655_0;
wire n_23493;
wire n_26083;
wire FE_OFN798_n_46285;
wire n_39512;
wire n_38205;
wire newNet_1995;
wire FE_OCPN1383_n_18345;
wire n_27764;
wire n_25400;
wire FE_OCP_RBN3069_n_43230;
wire n_17344;
wire n_27605;
wire n_35472;
wire n_152;
wire n_5465;
wire FE_RN_689_0;
wire n_30219;
wire n_39718;
wire n_16804;
wire n_14608;
wire n_32186;
wire newNet_1816;
wire newNet_913;
wire newNet_788;
wire newNet_385;
wire n_7490;
wire FE_RN_1834_0;
wire n_35767;
wire n_42013;
wire n_32507;
wire newNet_2412;
wire n_13638;
wire FE_OCP_RBN3668_n_20812;
wire FE_RN_1293_0;
wire n_17444;
wire n_9089;
wire n_34385;
wire n_42163;
wire n_10386;
wire n_4200;
wire n_10481;
wire n_2018;
wire delay_add_ln22_unr5_stage3_stallmux_q_5_;
wire n_13792;
wire delay_add_ln22_unr14_stage6_stallmux_q_2_;
wire n_41798;
wire newNet_879;
wire n_16189;
wire n_36424;
wire n_28511;
wire n_38860;
wire newNet_2302;
wire n_3985;
wire n_43543;
wire n_19789;
wire n_1778;
wire n_41673;
wire n_3831;
wire n_30540;
wire n_39259;
wire n_34714;
wire n_31314;
wire n_2137;
wire n_22398;
wire n_41284;
wire n_11064;
wire n_26623;
wire FE_OCPN3186_FE_OCP_RBN1140_n_25816;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_12_;
wire n_5330;
wire n_27498;
wire n_36393;
wire newNet_3612;
wire n_6601;
wire newNet_3269;
wire FE_RN_1764_0;
wire n_9377;
wire n_28381;
wire n_34105;
wire n_28625;
wire n_24064;
wire n_40684;
wire FE_RN_1011_0;
wire n_22495;
wire n_21837;
wire n_2962;
wire n_29140;
wire n_22567;
wire n_6036;
wire n_17629;
wire n_38405;
wire n_7414;
wire n_916;
wire n_35457;
wire n_37743;
wire n_21178;
wire FE_OFN800_n_46285;
wire n_43850;
wire FE_OCPN1229_n_46101;
wire n_27615;
wire n_20632;
wire n_22672;
wire n_22011;
wire n_37711;
wire n_41977;
wire n_37544;
wire n_17088;
wire n_30258;
wire n_3480;
wire n_35648;
wire n_39215;
wire n_8549;
wire n_14323;
wire n_16509;
wire FE_OCP_RBN2864_n_39523;
wire n_34836;
wire n_14958;
wire newNet_3357;
wire FE_OCP_RBN3570_n_9188;
wire n_42387;
wire newNet_3150;
wire n_20954;
wire FE_OCP_RBN2792_n_9910;
wire n_31430;
wire FE_OCP_RBN2339_n_29385;
wire FE_OCP_RBN3653_n_10100;
wire n_2688;
wire n_11006;
wire n_38476;
wire newNet_1501;
wire n_21978;
wire FE_RN_1441_0;
wire n_3277;
wire n_20177;
wire n_11775;
wire n_19617;
wire n_31627;
wire n_15490;
wire n_29692;
wire n_20499;
wire n_3004;
wire n_41269;
wire FE_RN_1862_0;
wire n_15495;
wire FE_OCP_DRV_N1582_n_35500;
wire n_23181;
wire n_23869;
wire FE_RN_1296_0;
wire n_4336;
wire n_2930;
wire FE_RN_1471_0;
wire n_30465;
wire n_46228;
wire n_26956;
wire n_10597;
wire n_42817;
wire n_42153;
wire delay_add_ln22_unr8_stage4_stallmux_q_6_;
wire n_20395;
wire n_24908;
wire n_5430;
wire FE_OCP_RBN2944_FE_RN_1269_0;
wire n_10765;
wire n_26278;
wire FE_OCP_RBN3505_n_13860;
wire n_28515;
wire n_41402;
wire FE_OCPN931_n_40736;
wire n_1976;
wire n_12157;
wire n_45136;
wire FE_OCP_RBN3824_n_44061;
wire newNet_2967;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_27_;
wire n_3243;
wire n_28862;
wire newNet_2467;
wire n_22343;
wire n_33528;
wire n_24865;
wire n_26838;
wire n_38735;
wire n_42873;
wire FE_OCP_RBN3841_n_19419;
wire n_5377;
wire delay_add_ln22_unr5_stage3_stallmux_q_25_;
wire n_21694;
wire n_41745;
wire n_19836;
wire n_2785;
wire n_21735;
wire n_1478;
wire n_8205;
wire n_11251;
wire newNet_141;
wire n_33464;
wire n_6489;
wire n_2500;
wire n_14919;
wire n_38659;
wire FE_RN_1518_0;
wire n_30129;
wire n_34155;
wire n_10164;
wire n_26891;
wire n_8526;
wire FE_OCPN1511_n_22280;
wire n_29543;
wire n_25802;
wire n_2202;
wire n_14245;
wire n_17362;
wire n_10002;
wire n_35854;
wire n_2076;
wire n_38575;
wire FE_RN_1591_0;
wire n_3607;
wire n_42310;
wire n_7395;
wire n_15641;
wire n_32762;
wire n_32005;
wire delay_add_ln22_unr17_stage7_stallmux_q_31_;
wire n_43096;
wire newNet_315;
wire newNet_678;
wire newNet_7;
wire n_34978;
wire newNet_3702;
wire n_32579;
wire newNet_2152;
wire n_14184;
wire n_16288;
wire n_42367;
wire n_30405;
wire n_42105;
wire n_39931;
wire FE_RN_1824_0;
wire FE_OCP_RBN2243_n_13017;
wire n_28346;
wire n_41218;
wire FE_RN_979_0;
wire n_8977;
wire n_6065;
wire n_16750;
wire n_29816;
wire n_10508;
wire n_23659;
wire n_30622;
wire n_29944;
wire n_32496;
wire n_25585;
wire n_26557;
wire FE_OCP_RBN1327_n_36489;
wire n_42594;
wire n_35835;
wire newNet_3275;
wire n_879;
wire n_28115;
wire n_34874;
wire n_148;
wire n_42089;
wire n_38881;
wire FE_OCPN1463_n_29630;
wire FE_OCP_RBN1724_n_21004;
wire FE_RN_43_0;
wire FE_RN_441_0;
wire n_41824;
wire newNet_2512;
wire n_3154;
wire n_26757;
wire delay_xor_ln22_unr21_stage8_stallmux_q_9_;
wire n_23086;
wire n_11223;
wire n_11429;
wire n_39239;
wire n_29530;
wire n_38498;
wire n_35521;
wire newNet_1391;
wire n_45890;
wire delay_xor_ln21_unr15_stage6_stallmux_q_9_;
wire n_42530;
wire n_16406;
wire newNet_666;
wire n_33840;
wire n_34612;
wire n_30358;
wire n_16442;
wire n_15341;
wire n_8088;
wire n_24203;
wire n_37248;
wire FE_RN_882_0;
wire newNet_3393;
wire n_4486;
wire n_41810;
wire n_37105;
wire n_23211;
wire n_34299;
wire n_34394;
wire n_21722;
wire n_35571;
wire n_13684;
wire n_14042;
wire n_36339;
wire n_38917;
wire FE_OCPN3783_n_16463;
wire FE_RN_1541_0;
wire FE_OCP_RBN2998_n_11004;
wire n_1773;
wire n_6583;
wire beta_21;
wire n_43493;
wire n_40993;
wire n_40044;
wire n_19182;
wire n_41131;
wire n_2550;
wire n_1456;
wire n_2221;
wire n_20555;
wire n_26806;
wire n_7706;
wire n_42419;
wire n_32555;
wire n_28108;
wire delay_xor_ln22_unr12_stage5_stallmux_q_19_;
wire n_33476;
wire FE_OCP_RBN3442_n_37945;
wire n_29259;
wire n_1887;
wire n_39167;
wire n_33488;
wire n_15231;
wire FE_OCP_RBN1378_n_20889;
wire n_40333;
wire n_35888;
wire n_10898;
wire n_47026;
wire n_18346;
wire n_43874;
wire newNet_77;
wire n_25710;
wire n_37612;
wire n_29428;
wire n_21888;
wire newNet_1277;
wire n_6142;
wire FE_RN_1464_0;
wire n_7335;
wire n_13288;
wire newNet_1155;
wire newNet_1431;
wire n_8113;
wire FE_OCP_RBN2445_n_29684;
wire n_46180;
wire FE_RN_835_0;
wire n_2667;
wire n_36045;
wire FE_OCPN1032_n_28448;
wire newNet_290;
wire n_10687;
wire n_469;
wire n_6084;
wire n_16419;
wire n_4422;
wire n_6941;
wire FE_OFN813_n_2540;
wire n_31176;
wire n_7390;
wire n_35241;
wire n_22913;
wire n_18667;
wire n_21165;
wire n_29769;
wire n_4968;
wire n_26097;
wire newNet_849;
wire n_5744;
wire FE_RN_1708_0;
wire n_29339;
wire FE_RN_741_0;
wire n_859;
wire n_4443;
wire n_1727;
wire delay_add_ln22_unr20_stage8_stallmux_q_13_;
wire n_11154;
wire FE_RN_564_0;
wire n_8677;
wire n_22865;
wire FE_OCP_RBN3099_n_32001;
wire n_11387;
wire n_16384;
wire n_26905;
wire newNet_2408;
wire n_204;
wire n_4600;
wire n_9798;
wire n_13419;
wire n_24924;
wire FE_RN_69_0;
wire n_13281;
wire n_27422;
wire n_15627;
wire n_40984;
wire n_24277;
wire n_4684;
wire n_3462;
wire n_21686;
wire n_27635;
wire FE_OCP_RBN3487_n_2438;
wire n_11475;
wire n_5857;
wire FE_OCP_DRV_N1545_n_18860;
wire delay_xor_ln21_unr9_stage4_stallmux_q_3_;
wire n_23716;
wire n_2069;
wire n_35794;
wire n_44100;
wire newNet_2019;
wire n_20057;
wire n_34126;
wire n_9774;
wire n_15351;
wire n_41180;
wire n_18998;
wire n_5268;
wire n_37329;
wire newNet_1217;
wire FE_OCP_RBN2198_n_41256;
wire n_43089;
wire n_28648;
wire n_31671;
wire n_32542;
wire n_14897;
wire newNet_229;
wire n_16009;
wire FE_OCP_RBN3049_n_11329;
wire delay_add_ln22_unr5_stage3_stallmux_q_24_;
wire n_6859;
wire n_2975;
wire n_23647;
wire n_21787;
wire n_32820;
wire n_36441;
wire newNet_2183;
wire FE_OCPN1799_FE_OFN780_n_17093;
wire n_45304;
wire n_15063;
wire n_25518;
wire n_23007;
wire n_1288;
wire n_20804;
wire n_33308;
wire FE_OCP_RBN3724_n_16975;
wire n_22066;
wire FE_RN_1046_0;
wire n_10876;
wire n_38444;
wire n_38342;
wire n_2344;
wire FE_OCP_RBN2411_n_13960;
wire n_26049;
wire FE_OCP_RBN1380_n_21240;
wire newNet_3020;
wire n_22757;
wire n_28545;
wire n_8602;
wire n_29456;
wire FE_OCP_RBN3701_n_31064;
wire newNet_1022;
wire n_12910;
wire n_39880;
wire n_39769;
wire FE_OCPN1528_n_26296;
wire n_37648;
wire FE_OCP_RBN2767_n_4376;
wire n_173;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_10_;
wire n_3226;
wire n_12817;
wire n_41079;
wire n_23942;
wire FE_RN_477_0;
wire n_4923;
wire n_15666;
wire n_47241;
wire n_23238;
wire newNet_2535;
wire FE_OCP_RBN2844_n_10326;
wire n_18618;
wire n_23590;
wire n_10531;
wire n_32674;
wire FE_RN_489_0;
wire n_32898;
wire n_34657;
wire n_16333;
wire FE_RN_1477_0;
wire newNet_456;
wire n_10944;
wire n_27233;
wire n_27638;
wire n_21980;
wire newNet_2948;
wire n_4620;
wire delay_add_ln22_unr17_stage7_stallmux_q_10_;
wire delay_add_ln22_unr14_stage6_stallmux_q_31_;
wire n_6847;
wire n_45716;
wire n_21814;
wire n_2901;
wire n_12534;
wire n_31014;
wire n_5879;
wire FE_OCP_RBN2824_n_10068;
wire n_20650;
wire n_19707;
wire n_35335;
wire FE_OCP_RBN3222_n_22068;
wire FE_OCP_DRV_N3742_n_25400;
wire n_40176;
wire n_29722;
wire n_18039;
wire n_23693;
wire n_32145;
wire n_32021;
wire n_35377;
wire newNet_1573;
wire n_7114;
wire n_22106;
wire n_20092;
wire n_20962;
wire n_17682;
wire n_29790;
wire FE_OCP_RBN3365_n_44722;
wire FE_OCP_RBN2859_n_10399;
wire n_38366;
wire n_29776;
wire n_41713;
wire n_26233;
wire n_39044;
wire newNet_1408;
wire n_41316;
wire FE_OCP_RBN2352_n_38534;
wire n_39711;
wire n_4479;
wire n_2706;
wire n_8610;
wire n_20664;
wire n_42355;
wire n_27486;
wire n_41206;
wire n_35953;
wire n_38903;
wire n_25092;
wire n_22113;
wire FE_RN_1561_0;
wire n_4995;
wire n_32966;
wire n_14532;
wire FE_RN_467_0;
wire n_14641;
wire n_40072;
wire delay_xor_ln21_unr15_stage6_stallmux_q_12_;
wire FE_RN_42_0;
wire n_12663;
wire n_11113;
wire n_23762;
wire n_12986;
wire n_16355;
wire n_32886;
wire newNet_2699;
wire n_1172;
wire n_34587;
wire n_42342;
wire n_31929;
wire newNet_874;
wire n_24115;
wire n_42789;
wire n_18391;
wire n_3448;
wire n_19114;
wire n_20032;
wire n_4248;
wire n_26300;
wire n_22840;
wire n_17335;
wire n_19849;
wire n_33253;
wire n_39477;
wire n_40197;
wire n_19653;
wire n_15686;
wire FE_OCPN3177_n_21901;
wire newNet_1034;
wire n_2235;
wire n_763;
wire n_13794;
wire n_6262;
wire n_8096;
wire n_15772;
wire FE_OCP_RBN2332_n_29380;
wire n_14921;
wire n_16636;
wire n_38712;
wire n_35030;
wire n_40463;
wire n_2676;
wire n_34169;
wire n_34210;
wire newNet_3714;
wire n_39336;
wire n_25335;
wire n_11180;
wire n_14563;
wire n_8753;
wire n_42550;
wire n_17033;
wire newNet_1322;
wire FE_RN_523_0;
wire n_4215;
wire n_17152;
wire n_34848;
wire FE_OFN777_n_17093;
wire n_31308;
wire n_4302;
wire n_11131;
wire n_19098;
wire n_32465;
wire n_9391;
wire n_4830;
wire n_15337;
wire n_18784;
wire n_35507;
wire newNet_3282;
wire n_1707;
wire FE_OCP_RBN2602_n_39126;
wire n_23901;
wire n_6442;
wire n_3740;
wire delay_add_ln22_unr14_stage6_stallmux_q_3_;
wire n_7481;
wire n_34552;
wire newNet_534;
wire n_1239;
wire FE_OCP_RBN2694_n_15083;
wire n_1131;
wire n_18354;
wire n_4734;
wire FE_OCPN1413_n_19715;
wire FE_OCPN858_n_45697;
wire n_5077;
wire n_14664;
wire n_31902;
wire n_31051;
wire n_36621;
wire newNet_732;
wire n_17644;
wire n_35174;
wire n_32788;
wire n_20857;
wire n_5760;
wire n_8743;
wire newNet_2369;
wire n_35700;
wire n_27706;
wire n_32094;
wire n_19340;
wire n_15109;
wire n_18898;
wire n_23057;
wire n_3251;
wire n_5082;
wire n_10579;
wire n_38691;
wire n_20214;
wire n_34745;
wire n_41617;
wire n_18735;
wire n_19715;
wire n_6343;
wire n_35788;
wire newNet_3453;
wire n_17329;
wire n_18718;
wire n_18602;
wire n_35060;
wire newNet_599;
wire n_1552;
wire n_21504;
wire newNet_1923;
wire n_42806;
wire n_20854;
wire n_42304;
wire n_10245;
wire n_18845;
wire n_13865;
wire n_19854;
wire n_26993;
wire newNet_1832;
wire n_20729;
wire FE_OCP_RBN3547_n_44575;
wire n_23463;
wire newNet_1048;
wire n_2620;
wire n_18437;
wire n_2128;
wire n_9848;
wire n_26307;
wire FE_RN_1206_0;
wire n_29832;
wire delay_add_ln22_unr8_stage4_stallmux_q_18_;
wire newNet_893;
wire n_7614;
wire n_5999;
wire n_25251;
wire n_36962;
wire n_12694;
wire n_3355;
wire n_28135;
wire n_17096;
wire n_38425;
wire n_34179;
wire FE_OCP_RBN3407_n_28597;
wire FE_OCP_RBN2327_n_29378;
wire n_27211;
wire n_35748;
wire FE_OCP_RBN2600_n_34388;
wire newNet_122;
wire n_30262;
wire n_17428;
wire n_24006;
wire FE_OCPN3771_n_8669;
wire n_41293;
wire n_29744;
wire n_22139;
wire n_3929;
wire n_46209;
wire n_6752;
wire n_31005;
wire n_34060;
wire newNet_48;
wire n_58;
wire n_12867;
wire n_6875;
wire n_18434;
wire n_35946;
wire FE_OCPUNCON1808_n_31435;
wire newNet_2910;
wire n_36934;
wire newNet_434;
wire n_38309;
wire FE_RN_968_0;
wire n_43455;
wire n_22621;
wire n_37707;
wire n_9016;
wire FE_OCPN1767_n_29715;
wire n_11786;
wire n_17494;
wire n_453;
wire newNet_3311;
wire n_11584;
wire FE_RN_1798_0;
wire n_11299;
wire n_12464;
wire n_17020;
wire n_40156;
wire n_7448;
wire n_18013;
wire n_17923;
wire n_16726;
wire n_35569;
wire newNet_1696;
wire n_31934;
wire n_16943;
wire newNet_1619;
wire n_9698;
wire newNet_1793;
wire newNet_2598;
wire n_40223;
wire n_4078;
wire n_8184;
wire n_37970;
wire newNet_2872;
wire FE_RN_1540_0;
wire n_4814;
wire n_43428;
wire n_8175;
wire n_10314;
wire n_9126;
wire n_9002;
wire n_5144;
wire newNet_2228;
wire n_7933;
wire n_31455;
wire n_636;
wire n_12476;
wire n_19028;
wire n_29755;
wire n_7495;
wire n_35969;
wire n_11464;
wire n_13557;
wire n_5169;
wire n_1087;
wire n_46418;
wire FE_RN_942_0;
wire n_23220;
wire n_14573;
wire n_47333;
wire delay_add_ln22_unr17_stage7_stallmux_q_28_;
wire n_7936;
wire n_39271;
wire n_23544;
wire n_28848;
wire n_32389;
wire n_32994;
wire n_36577;
wire n_32628;
wire n_22949;
wire FE_OCP_RBN3698_n_35543;
wire n_43588;
wire n_2510;
wire newNet_1268;
wire n_19046;
wire n_39661;
wire n_26665;
wire n_23104;
wire n_263;
wire FE_RN_1368_0;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_16_;
wire n_42172;
wire n_3700;
wire n_33963;
wire n_43489;
wire n_29581;
wire n_35844;
wire n_37733;
wire n_40420;
wire n_43519;
wire n_32416;
wire n_41984;
wire n_19539;
wire newNet_3408;
wire n_1200;
wire n_21998;
wire n_32845;
wire n_26248;
wire n_25073;
wire n_2095;
wire n_1083;
wire n_5061;
wire n_11325;
wire n_9762;
wire n_105;
wire n_7434;
wire newNet_1197;
wire n_36208;
wire n_19383;
wire n_16746;
wire n_19083;
wire n_22879;
wire n_32249;
wire n_10622;
wire n_27;
wire n_31230;
wire n_36034;
wire n_43368;
wire n_26116;
wire n_19505;
wire newNet_377;
wire n_11901;
wire n_28643;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_26_;
wire n_28045;
wire n_33438;
wire n_34794;
wire FE_OCPN1044_n_20307;
wire n_4541;
wire n_27066;
wire n_27406;
wire n_12211;
wire n_31391;
wire n_46997;
wire n_31078;
wire n_17133;
wire n_34404;
wire newNet_1911;
wire n_7128;
wire newNet_3171;
wire n_25429;
wire FE_OCP_RBN2437_n_8402;
wire n_4650;
wire n_5010;
wire n_11960;
wire n_700;
wire FE_RN_1756_0;
wire n_42116;
wire n_16163;
wire n_7567;
wire n_43515;
wire n_9095;
wire newNet_1938;
wire FE_RN_1282_0;
wire n_14887;
wire n_18944;
wire n_1109;
wire n_21317;
wire n_34842;
wire FE_OCPN1732_n_34369;
wire n_28027;
wire n_17237;
wire FE_OCP_DRV_N1578_n_33904;
wire n_15818;
wire n_11835;
wire FE_RN_1339_0;
wire n_259;
wire n_1851;
wire n_41087;
wire n_16571;
wire n_30897;
wire n_31581;
wire n_29017;
wire n_34809;
wire n_41303;
wire n_37256;
wire newNet_885;
wire n_3651;
wire n_9450;
wire newNet_3044;
wire n_12540;
wire n_26149;
wire n_26654;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_24_;
wire n_29715;
wire n_33407;
wire n_35552;
wire newNet_3069;
wire n_6800;
wire n_627;
wire n_38993;
wire n_1358;
wire n_32475;
wire n_21759;
wire n_33832;
wire n_270;
wire newNet_1306;
wire FE_OCP_RBN2453_n_38537;
wire n_17908;
wire n_10953;
wire n_5208;
wire newNet_1891;
wire n_28684;
wire n_29098;
wire n_4860;
wire n_8268;
wire FE_OCP_RBN2118_n_45224;
wire n_43642;
wire n_31490;
wire n_12321;
wire n_21798;
wire FE_RN_804_0;
wire n_400;
wire n_43259;
wire n_9835;
wire n_41690;
wire n_9616;
wire n_33668;
wire n_43862;
wire n_31164;
wire newNet_708;
wire n_30425;
wire n_6257;
wire n_8432;
wire n_12360;
wire n_41504;
wire n_17482;
wire newNet_2471;
wire n_33238;
wire FE_OCPN884_n_42216;
wire n_34300;
wire n_41735;
wire n_7288;
wire n_22476;
wire newNet_935;
wire n_30711;
wire n_3816;
wire n_10341;
wire n_792;
wire n_39721;
wire n_20206;
wire n_41002;
wire n_37331;
wire FE_RN_1310_0;
wire n_46192;
wire n_10892;
wire n_37825;
wire n_4592;
wire n_23875;
wire n_36986;
wire n_10808;
wire n_31254;
wire n_26295;
wire n_16092;
wire n_9627;
wire n_9620;
wire n_11358;
wire n_37512;
wire n_18048;
wire FE_RN_313_0;
wire n_25208;
wire newNet_517;
wire n_41995;
wire n_3304;
wire n_22309;
wire n_7657;
wire n_11671;
wire n_25377;
wire n_33218;
wire n_7215;
wire n_19765;
wire n_26424;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_1_;
wire n_339;
wire n_34096;
wire n_32742;
wire n_24002;
wire n_17866;
wire newNet_270;
wire n_16494;
wire FE_OCP_RBN2425_n_47023;
wire n_7356;
wire n_13228;
wire n_6147;
wire n_36684;
wire n_37472;
wire n_7735;
wire n_10157;
wire n_40919;
wire n_13322;
wire n_25416;
wire n_5459;
wire n_24616;
wire n_37303;
wire newNet_3266;
wire n_11419;
wire FE_OCPN967_n_19342;
wire n_11913;
wire n_16734;
wire n_15094;
wire FE_OCP_RBN3590_n_47014;
wire newNet_1787;
wire n_199;
wire n_21049;
wire n_42860;
wire n_36704;
wire n_5156;
wire n_32452;
wire n_43233;
wire n_1042;
wire n_28989;
wire n_37151;
wire n_27337;
wire n_18516;
wire n_593;
wire n_16921;
wire n_35065;
wire n_27430;
wire n_19120;
wire n_42306;
wire n_121;
wire n_22773;
wire n_24685;
wire n_280;
wire n_679;
wire n_28246;
wire n_897;
wire delay_add_ln22_unr5_stage3_stallmux_q_14_;
wire n_24402;
wire n_37311;
wire n_1517;
wire n_25911;
wire n_42927;
wire n_38160;
wire n_5351;
wire n_1166;
wire n_25366;
wire n_12188;
wire n_17005;
wire n_19845;
wire n_44352;
wire n_25705;
wire n_17548;
wire FE_RN_1699_0;
wire n_7323;
wire n_18232;
wire n_25112;
wire n_42329;
wire n_27134;
wire n_37505;
wire n_32058;
wire n_43856;
wire n_25467;
wire n_38532;
wire delay_xor_ln22_unr3_stage2_stallmux_q_4_;
wire n_11142;
wire FE_OCP_DRV_N1541_n_26125;
wire n_3169;
wire n_13302;
wire FE_OCP_RBN3616_n_20249;
wire n_6935;
wire n_25247;
wire n_30803;
wire n_36199;
wire n_25984;
wire newNet_213;
wire n_36143;
wire n_32328;
wire n_19236;
wire n_31291;
wire FE_RN_1842_0;
wire n_23789;
wire n_7219;
wire newNet_1050;
wire n_18387;
wire n_8634;
wire FE_RN_395_0;
wire n_38230;
wire n_33188;
wire n_20571;
wire n_5881;
wire FE_OCP_RBN3089_FE_OCPN1052_n_31674;
wire n_10392;
wire n_23542;
wire n_13671;
wire n_36698;
wire n_16874;
wire n_31263;
wire n_11049;
wire n_37001;
wire n_43179;
wire n_8617;
wire n_17435;
wire n_8352;
wire n_37365;
wire n_24250;
wire FE_OCP_RBN3685_n_5217;
wire n_29659;
wire FE_OCP_RBN1139_n_25816;
wire n_646;
wire n_23907;
wire n_15114;
wire n_5751;
wire FE_RN_859_0;
wire n_8462;
wire n_7461;
wire n_27076;
wire n_4639;
wire n_22149;
wire n_4881;
wire n_26886;
wire newNet_3550;
wire n_37290;
wire n_11482;
wire n_18599;
wire n_23310;
wire n_25676;
wire n_34684;
wire n_16917;
wire delay_xor_ln21_unr6_stage3_stallmux_q_0_;
wire newNet_3293;
wire n_46424;
wire n_16030;
wire n_46158;
wire delay_xor_ln22_unr6_stage3_stallmux_q_8_;
wire n_24704;
wire FE_OCPN945_n_1780;
wire n_16303;
wire n_14260;
wire n_1953;
wire FE_OCP_RBN2819_n_4872;
wire n_43387;
wire n_8867;
wire newNet_490;
wire n_45828;
wire n_18697;
wire newNet_135;
wire n_5049;
wire n_33984;
wire n_29486;
wire n_11767;
wire n_37014;
wire n_1496;
wire n_36224;
wire n_29518;
wire n_24692;
wire n_39085;
wire n_21197;
wire n_22669;
wire n_12239;
wire n_26417;
wire FE_OCPN890_n_7802;
wire n_18424;
wire n_27865;
wire n_21565;
wire n_25567;
wire n_29280;
wire newNet_649;
wire n_30926;
wire n_36376;
wire n_43229;
wire n_41249;
wire n_20018;
wire n_2396;
wire n_3208;
wire n_14192;
wire FE_OCPN1764_n_13646;
wire n_25757;
wire n_42226;
wire n_36731;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_6_;
wire n_33590;
wire n_10811;
wire n_9119;
wire FE_RN_461_0;
wire n_45623;
wire n_14974;
wire n_25357;
wire newNet_2720;
wire n_7854;
wire n_24190;
wire n_18562;
wire n_25287;
wire n_17367;
wire n_18190;
wire n_25015;
wire n_6048;
wire n_11808;
wire n_10566;
wire n_8668;
wire n_26540;
wire n_43662;
wire n_9285;
wire n_37167;
wire n_11383;
wire n_24054;
wire FE_OCP_RBN3249_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_19497;
wire n_27913;
wire n_6189;
wire n_37581;
wire n_7268;
wire n_479;
wire n_21862;
wire n_29288;
wire FE_OCP_RBN2656_FE_RN_1288_0;
wire n_38674;
wire n_2882;
wire n_160;
wire n_2985;
wire n_25087;
wire delay_xor_ln21_unr6_stage3_stallmux_q_22_;
wire n_29809;
wire FE_RN_1302_0;
wire FE_RN_451_0;
wire n_35393;
wire n_2480;
wire n_36074;
wire n_33118;
wire n_17460;
wire newNet_314;
wire newNet_1508;
wire n_24295;
wire n_34504;
wire n_15990;
wire n_6572;
wire n_29029;
wire n_3991;
wire n_640;
wire n_2755;
wire n_7014;
wire n_8284;
wire n_8752;
wire n_24176;
wire n_33225;
wire newNet_3309;
wire FE_RN_57_0;
wire n_36194;
wire newNet_1359;
wire n_1077;
wire n_6926;
wire n_11162;
wire n_28689;
wire newNet_53;
wire n_17055;
wire n_33043;
wire n_38406;
wire n_33737;
wire n_26208;
wire newNet_2414;
wire n_7922;
wire n_38940;
wire n_37252;
wire n_32157;
wire FE_RN_1707_0;
wire n_19978;
wire n_28088;
wire n_32851;
wire n_1919;
wire n_39191;
wire FE_OCP_RBN3383_n_12365;
wire n_39642;
wire n_1803;
wire n_5301;
wire delay_xor_ln22_unr3_stage2_stallmux_q_28_;
wire n_31854;
wire n_4085;
wire n_12319;
wire newNet_157;
wire n_828;
wire n_24406;
wire n_22420;
wire n_32837;
wire n_46960;
wire n_10058;
wire n_32390;
wire n_29260;
wire FE_OFN826_n_1142;
wire n_9265;
wire n_16088;
wire n_7718;
wire n_20512;
wire n_19579;
wire state_cordic_1_;
wire n_974;
wire FE_RN_382_0;
wire n_22726;
wire n_14109;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_9_;
wire n_12429;
wire n_33599;
wire n_36842;
wire n_26644;
wire n_28750;
wire n_27784;
wire n_19612;
wire n_12487;
wire n_10429;
wire n_46952;
wire FE_OCP_RBN3537_n_8597;
wire n_3970;
wire n_23504;
wire newNet_400;
wire n_14862;
wire n_10195;
wire n_25597;
wire n_29890;
wire n_37988;
wire n_3157;
wire FE_OCP_RBN2557_n_44576;
wire n_10112;
wire FE_OCPN1437_FE_OCP_RBN1330_n_18866;
wire n_29898;
wire n_40959;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_6_;
wire n_6770;
wire n_39000;
wire n_18072;
wire n_42213;
wire newNet_1874;
wire n_14066;
wire n_41814;
wire n_20989;
wire newNet_624;
wire FE_RN_1747_0;
wire n_3575;
wire n_28338;
wire newNet_66;
wire n_23502;
wire n_40303;
wire n_3178;
wire FE_OCP_RBN2823_n_10068;
wire n_6011;
wire n_29065;
wire delay_add_ln22_unr2_stage2_stallmux_q_19_;
wire n_40748;
wire n_21903;
wire FE_OCPN1494_n_23398;
wire n_29361;
wire newNet_1607;
wire n_32125;
wire n_7110;
wire FE_RN_1081_0;
wire n_30192;
wire n_29566;
wire n_28869;
wire n_22745;
wire n_45511;
wire n_32535;
wire n_17828;
wire n_3308;
wire n_16399;
wire n_7473;
wire newNet_544;
wire n_3665;
wire FE_OCP_RBN2507_n_13896;
wire n_15909;
wire n_42037;
wire n_37729;
wire n_13721;
wire n_31701;
wire n_28057;
wire delay_xor_ln22_unr3_stage2_stallmux_q_16_;
wire n_41070;
wire n_34272;
wire delay_xor_ln21_unr12_stage5_stallmux_q_2_;
wire n_25977;
wire n_43291;
wire n_623;
wire n_3701;
wire n_27299;
wire newNet_2107;
wire newNet_1724;
wire n_27017;
wire n_29869;
wire n_39533;
wire FE_OCP_RBN2640_n_34921;
wire n_14994;
wire n_6599;
wire n_39815;
wire n_27397;
wire n_15945;
wire delay_xor_ln21_unr9_stage4_stallmux_q_2_;
wire n_13856;
wire n_45012;
wire FE_RN_484_0;
wire n_41920;
wire n_45474;
wire n_3013;
wire n_34436;
wire n_17880;
wire n_18985;
wire FE_OCPN1427_n_13510;
wire n_10709;
wire n_8176;
wire n_12644;
wire n_17593;
wire n_26931;
wire n_30643;
wire delay_add_ln22_unr20_stage8_stallmux_q_17_;
wire n_8729;
wire n_12393;
wire FE_OCP_DRV_N1610_n_20146;
wire n_19301;
wire n_15196;
wire n_11921;
wire FE_OCP_RBN1688_n_18986;
wire n_1032;
wire n_13404;
wire n_39536;
wire FE_RN_1279_0;
wire n_10772;
wire n_21220;
wire newNet_1203;
wire newNet_698;
wire n_20768;
wire n_25008;
wire n_32504;
wire n_41757;
wire n_1965;
wire n_6386;
wire delay_xor_ln22_unr12_stage5_stallmux_q_14_;
wire FE_RN_630_0;
wire n_25552;
wire n_27534;
wire newNet_1289;
wire n_7051;
wire n_13804;
wire n_33998;
wire n_41663;
wire n_14251;
wire n_35696;
wire n_21804;
wire n_18085;
wire FE_RN_1266_0;
wire n_13698;
wire n_43820;
wire n_8345;
wire n_24147;
wire n_39703;
wire n_38869;
wire n_43434;
wire FE_OFN839_n_4597;
wire n_43574;
wire n_33626;
wire n_7316;
wire n_10473;
wire n_35102;
wire n_7731;
wire n_18641;
wire n_34149;
wire n_15952;
wire n_13652;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_11_;
wire n_4480;
wire n_31872;
wire n_16290;
wire n_24386;
wire n_19787;
wire n_7408;
wire n_29668;
wire n_37238;
wire n_16599;
wire n_26817;
wire FE_OCP_RBN2952_n_21489;
wire n_30886;
wire n_21203;
wire n_16235;
wire n_23637;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_30_;
wire n_19862;
wire n_521;
wire n_36297;
wire n_7171;
wire n_36322;
wire FE_OCPN3170_n_23227;
wire n_12312;
wire n_24700;
wire n_19999;
wire n_14525;
wire n_30412;
wire newNet_2603;
wire n_39811;
wire n_15531;
wire n_9395;
wire n_20301;
wire n_2081;
wire n_14196;
wire n_26831;
wire n_7468;
wire FE_OCP_RBN2960_n_26231;
wire n_12266;
wire n_30514;
wire n_6182;
wire n_35784;
wire n_33785;
wire n_21927;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_18_;
wire n_1860;
wire n_4496;
wire n_3764;
wire n_22543;
wire n_18650;
wire n_15168;
wire n_5247;
wire n_36743;
wire n_30879;
wire n_43796;
wire n_33925;
wire newNet_1702;
wire newNet_1833;
wire FE_OCP_RBN1705_n_21658;
wire n_1836;
wire n_10934;
wire n_20211;
wire n_2738;
wire n_11184;
wire FE_OCP_RBN3051_n_16596;
wire n_43157;
wire FE_RN_1691_0;
wire n_18279;
wire n_7961;
wire n_5558;
wire n_28739;
wire n_19375;
wire n_16314;
wire n_43066;
wire n_28580;
wire n_8191;
wire n_21222;
wire n_28005;
wire FE_RN_5_0;
wire n_4669;
wire n_17252;
wire FE_OCP_RBN2111_n_11548;
wire n_18020;
wire n_35355;
wire n_2536;
wire n_29291;
wire n_5339;
wire n_41120;
wire n_22935;
wire newNet_3337;
wire n_6734;
wire n_41230;
wire n_2660;
wire n_10053;
wire newNet_3138;
wire n_15258;
wire n_10559;
wire n_29400;
wire FE_RN_603_0;
wire FE_OCP_RBN3656_n_25997;
wire n_14335;
wire n_24078;
wire n_22940;
wire n_32144;
wire FE_RN_1492_0;
wire n_44428;
wire newNet_630;
wire n_37386;
wire n_27858;
wire n_47274;
wire n_8981;
wire delay_xor_ln22_unr12_stage5_stallmux_q_10_;
wire n_22095;
wire n_4219;
wire FE_OCPN3187_n_11012;
wire n_27222;
wire FE_OCP_RBN2272_n_13489;
wire n_8509;
wire n_10871;
wire n_13368;
wire n_23111;
wire n_33646;
wire n_3269;
wire n_18157;
wire FE_RN_371_0;
wire n_2699;
wire n_5795;
wire n_4852;
wire n_20311;
wire n_30085;
wire n_2229;
wire FE_RN_26_0;
wire FE_RN_1287_0;
wire n_2205;
wire n_18836;
wire n_5668;
wire FE_OCP_RBN2383_n_8342;
wire n_21346;
wire n_37272;
wire n_36230;
wire n_28555;
wire n_15854;
wire n_21748;
wire n_4435;
wire n_14333;
wire n_33335;
wire n_18201;
wire n_21374;
wire n_16937;
wire FE_OCP_RBN2152_n_22822;
wire n_36617;
wire delay_add_ln22_unr27_stage10_stallmux_q_26_;
wire n_14319;
wire n_35830;
wire n_177;
wire n_14670;
wire n_37939;
wire n_37176;
wire FE_OCP_RBN2335_n_24359;
wire n_19344;
wire n_11694;
wire n_12339;
wire n_1043;
wire newNet_746;
wire n_1874;
wire n_38159;
wire n_31094;
wire n_46344;
wire n_31115;
wire n_34064;
wire n_4275;
wire n_25155;
wire n_7675;
wire n_36633;
wire n_41364;
wire newNet_1770;
wire n_38502;
wire n_40538;
wire n_6565;
wire n_31831;
wire n_19724;
wire n_11216;
wire n_40861;
wire n_39964;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_19_;
wire n_4289;
wire n_24245;
wire n_13719;
wire n_25953;
wire n_20608;
wire n_24444;
wire n_33153;
wire n_11179;
wire n_25490;
wire n_32015;
wire n_36269;
wire n_25817;
wire n_15453;
wire n_12680;
wire FE_OCP_RBN2840_n_4692;
wire n_32549;
wire delay_add_ln22_unr11_stage5_stallmux_q_21_;
wire newNet_2256;
wire n_42679;
wire FE_RN_1558_0;
wire n_36187;
wire FE_RN_1792_0;
wire n_19656;
wire FE_RN_1029_0;
wire n_41472;
wire n_11336;
wire FE_OCP_RBN3492_n_29553;
wire FE_OCP_RBN3477_n_13756;
wire n_8335;
wire newNet_190;
wire n_15000;
wire n_33373;
wire n_9844;
wire n_1162;
wire n_4256;
wire n_33358;
wire n_34412;
wire n_26609;
wire n_9116;
wire n_24608;
wire n_28806;
wire n_3433;
wire n_15409;
wire n_26403;
wire n_12361;
wire n_243;
wire FE_RN_386_0;
wire n_18262;
wire n_29248;
wire n_8724;
wire FE_OCP_RBN1845_n_20910;
wire FE_OCP_RBN2321_n_2638;
wire n_2796;
wire FE_OCPN993_n_15552;
wire FE_RN_1462_0;
wire FE_RN_1642_0;
wire newNet_115;
wire n_24676;
wire FE_RN_685_0;
wire n_38124;
wire n_1268;
wire n_36273;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_11_;
wire FE_RN_1205_0;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_21_;
wire n_40923;
wire n_4879;
wire n_19212;
wire n_24014;
wire n_34926;
wire n_15236;
wire FE_OCP_RBN2221_n_13010;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_29_;
wire n_3435;
wire newNet_993;
wire n_43596;
wire n_3080;
wire n_28277;
wire FE_OCP_RBN3082_n_16977;
wire FE_OCP_RBN1330_n_18866;
wire FE_RN_1726_0;
wire n_19256;
wire n_36925;
wire n_7522;
wire n_822;
wire n_10202;
wire n_12706;
wire delay_add_ln22_unr5_stage3_stallmux_q_11_;
wire n_40859;
wire n_23459;
wire n_41202;
wire FE_RN_106_0;
wire n_8567;
wire n_14552;
wire n_38771;
wire newNet_2863;
wire n_41766;
wire n_27818;
wire n_18324;
wire n_457;
wire n_28295;
wire n_19913;
wire FE_RN_642_0;
wire n_8515;
wire n_41038;
wire n_8747;
wire n_15820;
wire n_7279;
wire FE_RN_1198_0;
wire n_41989;
wire n_39699;
wire n_30731;
wire newNet_182;
wire FE_RN_1521_0;
wire n_42733;
wire n_30377;
wire n_10310;
wire FE_OCP_DRV_N1540_n_35427;
wire n_43888;
wire newNet_2908;
wire n_31402;
wire n_41801;
wire n_8794;
wire FE_RN_779_0;
wire n_8309;
wire n_29771;
wire n_31425;
wire n_40719;
wire n_18318;
wire n_43764;
wire n_37522;
wire n_42242;
wire FE_OCP_RBN1218_n_21088;
wire newNet_1661;
wire n_40328;
wire newNet_1656;
wire n_32245;
wire n_31398;
wire n_43197;
wire n_965;
wire n_28036;
wire n_33967;
wire newNet_2914;
wire n_7124;
wire n_39980;
wire newNet_928;
wire n_30893;
wire n_2102;
wire n_28242;
wire n_8555;
wire n_36816;
wire n_41787;
wire n_4612;
wire newNet_2805;
wire FE_OCP_RBN2220_n_12888;
wire n_27883;
wire n_13217;
wire n_40799;
wire n_5136;
wire n_3347;
wire n_15465;
wire n_15742;
wire n_10163;
wire n_40785;
wire n_26927;
wire n_29025;
wire n_9470;
wire n_21586;
wire n_24840;
wire n_17331;
wire n_38384;
wire n_36942;
wire n_35712;
wire n_882;
wire n_25046;
wire n_25022;
wire n_2998;
wire n_30508;
wire n_37968;
wire FE_OCPN1498_n_26360;
wire n_25163;
wire n_27300;
wire n_35707;
wire n_13977;
wire n_4572;
wire n_30820;
wire n_37062;
wire n_8103;
wire n_15516;
wire n_30333;
wire n_34224;
wire newNet_3114;
wire n_16791;
wire n_28251;
wire n_38668;
wire n_2943;
wire n_35420;
wire n_8219;
wire n_21410;
wire n_29344;
wire n_13766;
wire newNet_3521;
wire n_16625;
wire FE_OCP_RBN3019_n_31117;
wire newNet_1010;
wire n_27284;
wire FE_OCP_RBN3086_n_31819;
wire n_30904;
wire newNet_3374;
wire n_41980;
wire newNet_72;
wire n_25099;
wire n_32922;
wire n_34763;
wire newNet_1839;
wire n_22644;
wire delay_xor_ln21_unr18_stage7_stallmux_q_5_;
wire n_28955;
wire n_12633;
wire n_29529;
wire n_39077;
wire n_5654;
wire FE_RN_1311_0;
wire n_2498;
wire newNet_1477;
wire n_22455;
wire n_28589;
wire n_10713;
wire n_27465;
wire FE_OCP_RBN3711_n_46337;
wire n_42539;
wire n_2286;
wire n_27973;
wire FE_RN_357_0;
wire n_5927;
wire FE_RN_1314_0;
wire n_21850;
wire n_42446;
wire newNet_1621;
wire n_10618;
wire FE_OCP_RBN3387_n_33108;
wire n_39450;
wire n_12760;
wire newNet_830;
wire n_31669;
wire n_43331;
wire newNet_3242;
wire newNet_880;
wire n_11031;
wire n_14409;
wire n_14428;
wire n_40566;
wire newNet_3693;
wire n_20459;
wire n_20959;
wire n_30348;
wire n_7309;
wire n_38373;
wire n_40737;
wire n_36781;
wire n_40710;
wire n_42067;
wire FE_OCP_RBN3597_FE_OCPN1243_n_44460;
wire n_5626;
wire n_10994;
wire n_42197;
wire n_24152;
wire n_2590;
wire n_12857;
wire n_8809;
wire delay_add_ln22_unr5_stage3_stallmux_q_21_;
wire n_43305;
wire n_43273;
wire n_6706;
wire n_46101;
wire n_28680;
wire n_31161;
wire FE_OCP_RBN2987_n_35539;
wire newNet_1483;
wire n_25605;
wire n_37914;
wire n_12069;
wire n_24109;
wire n_5896;
wire n_32800;
wire n_47265;
wire FE_OCP_RBN2589_n_9492;
wire newNet_3279;
wire newNet_1520;
wire n_2651;
wire n_31914;
wire FE_RN_522_0;
wire n_2300;
wire n_28207;
wire n_41964;
wire n_7754;
wire n_24872;
wire n_42509;
wire FE_RN_1849_0;
wire n_18850;
wire newNet_2370;
wire FE_OCP_DRV_N1557_n_19590;
wire newNet_1677;
wire n_34966;
wire n_46352;
wire n_6539;
wire n_38157;
wire n_42906;
wire delay_add_ln22_unr5_stage3_stallmux_q_20_;
wire n_32561;
wire n_37578;
wire FE_RN_697_0;
wire n_19695;
wire FE_RN_1391_0;
wire FE_RN_68_0;
wire n_11953;
wire n_12113;
wire n_38904;
wire n_35956;
wire n_34822;
wire n_24832;
wire n_25879;
wire n_34085;
wire FE_RN_280_0;
wire n_7254;
wire n_40492;
wire FE_OCP_RBN2712_n_35075;
wire n_14396;
wire n_42821;
wire n_28618;
wire n_10918;
wire n_45818;
wire newNet_460;
wire n_33604;
wire n_37032;
wire FE_OCP_RBN2776_n_15110;
wire n_36161;
wire n_35803;
wire delay_add_ln22_unr8_stage4_stallmux_q_15_;
wire n_40040;
wire n_25623;
wire n_9332;
wire newNet_1290;
wire n_12467;
wire n_34324;
wire FE_OCP_RBN3620_n_15135;
wire n_43651;
wire n_1781;
wire n_7134;
wire n_29859;
wire n_32730;
wire newNet_3053;
wire n_36545;
wire n_33495;
wire n_29595;
wire n_36147;
wire n_43817;
wire n_40485;
wire n_20782;
wire n_14063;
wire n_27793;
wire n_26532;
wire FE_OCP_DRV_N3158_n_27062;
wire n_9446;
wire n_19879;
wire n_25107;
wire n_27192;
wire n_34974;
wire n_11756;
wire n_19813;
wire n_10769;
wire n_21964;
wire FE_OCP_RBN1367_n_20763;
wire n_15038;
wire n_43378;
wire n_46151;
wire n_38766;
wire n_10521;
wire n_14418;
wire n_42767;
wire n_2031;
wire n_3404;
wire n_5571;
wire n_39629;
wire n_32230;
wire n_33632;
wire n_35462;
wire n_35673;
wire n_10691;
wire n_39278;
wire newNet_1541;
wire n_23420;
wire n_9955;
wire n_22527;
wire n_34792;
wire n_30655;
wire n_32240;
wire n_8878;
wire newNet_1193;
wire n_17027;
wire FE_RN_501_0;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_16_;
wire n_26639;
wire n_26741;
wire n_10288;
wire n_10045;
wire newNet_2280;
wire n_18172;
wire n_21239;
wire n_41881;
wire n_28890;
wire n_9978;
wire n_13126;
wire n_3698;
wire newNet_3082;
wire n_14889;
wire n_17085;
wire delay_xor_ln21_unr21_stage8_stallmux_q_1_;
wire newNet_3645;
wire FE_OCP_RBN2401_n_13954;
wire n_35093;
wire n_23382;
wire n_6815;
wire n_34706;
wire FE_RN_1175_0;
wire n_43840;
wire n_41372;
wire n_25793;
wire n_16857;
wire n_32657;
wire n_35400;
wire newNet_255;
wire n_23949;
wire n_3832;
wire n_6226;
wire n_23964;
wire newNet_1226;
wire n_33720;
wire newNet_754;
wire n_2800;
wire n_7422;
wire newNet_2891;
wire n_18405;
wire n_35185;
wire n_1787;
wire n_14006;
wire n_35145;
wire n_27743;
wire n_14660;
wire FE_OCPN1754_n_7225;
wire n_4745;
wire n_30240;
wire n_17049;
wire n_15438;
wire n_12039;
wire FE_OCP_RBN2704_n_9411;
wire n_23399;
wire n_42403;
wire n_19386;
wire FE_OCP_RBN3126_n_27632;
wire n_266;
wire n_7672;
wire newNet_1646;
wire n_6861;
wire n_44695;
wire n_389;
wire n_36896;
wire n_5819;
wire n_11281;
wire n_11725;
wire n_38349;
wire newNet_2748;
wire FE_OCPN965_n_47020;
wire n_27906;
wire n_30970;
wire FE_RN_1083_0;
wire n_14988;
wire n_27807;
wire n_31264;
wire n_6323;
wire n_6139;
wire n_41093;
wire FE_OCP_RBN2516_n_8657;
wire n_12518;
wire n_14546;
wire n_23035;
wire n_18963;
wire n_25672;
wire FE_OFN763_n_15670;
wire n_18729;
wire n_742;
wire FE_OCPN1448_n_27463;
wire n_29298;
wire n_14604;
wire n_39582;
wire n_23408;
wire n_1058;
wire n_6043;
wire n_19254;
wire FE_OCPN1763_n_13646;
wire n_24605;
wire n_16107;
wire FE_OCP_RBN3599_FE_OCPN1243_n_44460;
wire n_40647;
wire n_3561;
wire n_21101;
wire n_33326;
wire FE_OCP_RBN1692_n_19052;
wire n_40895;
wire n_2388;
wire n_42854;
wire newNet_1759;
wire n_10865;
wire n_2577;
wire n_9238;
wire newNet_1127;
wire n_1028;
wire n_16596;
wire n_39387;
wire newNet_1054;
wire n_12071;
wire n_10440;
wire n_17113;
wire n_42412;
wire n_1191;
wire n_3317;
wire n_8701;
wire n_35353;
wire n_38033;
wire n_11411;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_18_;
wire n_13732;
wire n_25182;
wire newNet_3245;
wire n_15223;
wire FE_OCP_RBN3269_n_45224;
wire n_37791;
wire FE_OCPN1438_FE_OCP_RBN1330_n_18866;
wire n_35168;
wire n_41942;
wire newNet_1365;
wire n_37245;
wire delay_add_ln22_unr14_stage6_stallmux_q_10_;
wire delay_add_ln22_unr17_stage7_stallmux_q_26_;
wire n_26464;
wire n_14483;
wire n_21489;
wire n_43333;
wire n_1185;
wire n_3140;
wire n_24858;
wire n_27859;
wire n_39509;
wire n_12738;
wire n_17656;
wire n_4340;
wire n_20137;
wire n_42974;
wire n_10223;
wire newNet_966;
wire n_16202;
wire newNet_2005;
wire n_3501;
wire n_7725;
wire n_25855;
wire newNet_2246;
wire n_20722;
wire n_35417;
wire delay_add_ln22_unr11_stage5_stallmux_q_28_;
wire n_4249;
wire n_5368;
wire delay_add_ln22_unr11_stage5_stallmux_q_12_;
wire n_19366;
wire FE_OCP_RBN2802_n_15706;
wire n_803;
wire n_40906;
wire newNet_1861;
wire n_21654;
wire n_17196;
wire n_34199;
wire newNet_3335;
wire FE_OFN810_n_1941;
wire n_43270;
wire n_29304;
wire n_18222;
wire n_36385;
wire n_3951;
wire n_4473;
wire n_23626;
wire n_14118;
wire n_26501;
wire n_39858;
wire n_888;
wire n_28841;
wire n_24644;
wire n_7973;
wire n_3415;
wire n_15739;
wire newNet_1583;
wire n_31570;
wire n_2402;
wire n_33193;
wire FE_OCPN3796_n_26115;
wire n_15487;
wire n_23563;
wire n_2548;
wire n_22061;
wire n_39148;
wire n_2741;
wire n_7859;
wire n_1749;
wire n_31058;
wire n_33281;
wire n_35298;
wire n_40408;
wire n_42637;
wire n_47336;
wire n_10875;
wire n_29952;
wire n_43007;
wire n_2715;
wire n_33561;
wire newNet_1604;
wire n_23928;
wire n_14199;
wire n_4771;
wire n_3802;
wire n_17697;
wire n_17584;
wire n_4730;
wire n_8885;
wire n_17573;
wire n_15084;
wire n_24581;
wire FE_OCP_RBN2927_n_39614;
wire n_12310;
wire FE_OCPN1015_n_32820;
wire n_4933;
wire n_46360;
wire n_41339;
wire newNet_1083;
wire n_43285;
wire n_1908;
wire n_43602;
wire n_12657;
wire n_21561;
wire FE_OFN806_n_46196;
wire n_21302;
wire n_5434;
wire n_34862;
wire FE_RN_1278_0;
wire newNet_361;
wire n_8386;
wire newNet_837;
wire n_33813;
wire FE_RN_466_0;
wire n_11074;
wire n_21180;
wire n_28283;
wire n_24953;
wire n_9685;
wire n_4404;
wire n_23185;
wire n_5590;
wire n_23561;
wire n_15679;
wire n_2089;
wire n_16787;
wire n_30317;
wire n_21932;
wire n_16122;
wire FE_RN_1539_0;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_1_;
wire newNet_2508;
wire n_23531;
wire FE_RN_839_0;
wire n_43017;
wire n_31502;
wire n_33429;
wire newNet_1060;
wire n_8921;
wire n_7061;
wire n_12582;
wire newNet_2356;
wire n_1569;
wire n_41252;
wire n_25521;
wire FE_OCP_DRV_N1594_n_34494;
wire FE_RN_210_0;
wire n_5151;
wire n_30485;
wire n_32318;
wire FE_RN_934_0;
wire n_33158;
wire n_1410;
wire n_39158;
wire n_39121;
wire n_27321;
wire FE_OCPN1489_n_30823;
wire n_2850;
wire n_15954;
wire n_12899;
wire n_43181;
wire n_17604;
wire delay_xor_ln21_unr18_stage7_stallmux_q_8_;
wire delay_xor_ln22_unr6_stage3_stallmux_q_24_;
wire newNet_3638;
wire n_34931;
wire n_16990;
wire n_18529;
wire FE_OCP_RBN2387_n_13860;
wire n_38511;
wire n_32795;
wire n_27109;
wire n_3828;
wire n_36661;
wire n_13996;
wire n_22799;
wire n_41569;
wire n_23731;
wire FE_OCP_RBN3094_n_11475;
wire n_2514;
wire n_9177;
wire n_22884;
wire n_24239;
wire newNet_2164;
wire n_10018;
wire n_32986;
wire FE_RN_576_0;
wire FE_OCP_RBN3726_FE_RN_1787_0;
wire n_21496;
wire n_26454;
wire n_18698;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_4_;
wire FE_OCPN1486_n_27315;
wire n_20616;
wire n_25904;
wire n_21056;
wire n_37869;
wire FE_OCP_RBN3664_n_35326;
wire FE_OCP_RBN2438_n_8402;
wire n_38286;
wire n_39595;
wire n_30760;
wire n_27087;
wire n_40385;
wire n_43031;
wire n_38435;
wire delay_xor_ln22_unr9_stage4_stallmux_q_18_;
wire n_45631;
wire n_24964;
wire n_26778;
wire n_18777;
wire n_22991;
wire n_42379;
wire n_9326;
wire n_18969;
wire n_22856;
wire n_14840;
wire n_17469;
wire n_25290;
wire n_12768;
wire n_44871;
wire n_33112;
wire n_33263;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_2_;
wire n_26433;
wire n_23616;
wire n_7278;
wire n_16435;
wire n_39610;
wire n_1128;
wire n_38312;
wire n_25356;
wire n_33576;
wire newNet_2975;
wire n_4972;
wire n_38448;
wire n_409;
wire n_27832;
wire n_7207;
wire n_12225;
wire n_41290;
wire n_5497;
wire n_38146;
wire n_24668;
wire n_36457;
wire n_31523;
wire n_41047;
wire n_4164;
wire n_39744;
wire n_36178;
wire n_43248;
wire newNet_1424;
wire n_36506;
wire n_4174;
wire newNet_163;
wire n_38;
wire n_38209;
wire n_21685;
wire FE_RN_454_0;
wire newNet_3320;
wire n_9703;
wire n_24597;
wire n_43214;
wire n_7342;
wire n_19885;
wire n_42967;
wire n_17404;
wire n_19601;
wire n_5007;
wire newNet_1174;
wire n_37412;
wire n_42465;
wire n_16533;
wire n_19233;
wire n_39738;
wire n_29841;
wire n_36084;
wire n_29926;
wire n_41221;
wire newNet_3031;
wire n_7646;
wire n_13621;
wire n_5777;
wire FE_OCP_RBN3428_n_12890;
wire n_14493;
wire n_24488;
wire n_2333;
wire n_40888;
wire n_21791;
wire n_28230;
wire n_4112;
wire n_40412;
wire n_36820;
wire n_43123;
wire n_25041;
wire n_16330;
wire n_29689;
wire n_43356;
wire n_43070;
wire n_39726;
wire n_4677;
wire n_21754;
wire n_2435;
wire n_15790;
wire n_28018;
wire n_26368;
wire n_2465;
wire FE_OCP_RBN2997_n_11004;
wire n_42890;
wire n_26653;
wire n_31384;
wire FE_OCP_RBN3456_n_33872;
wire n_2473;
wire n_14155;
wire n_84;
wire n_38998;
wire n_892;
wire n_6698;
wire n_35371;
wire n_41571;
wire n_33124;
wire n_22769;
wire n_24719;
wire newNet_2219;
wire FE_RN_687_0;
wire newNet_1468;
wire n_5918;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_23_;
wire n_29846;
wire FE_OCP_RBN3273_n_45224;
wire n_46224;
wire n_18758;
wire FE_RN_536_0;
wire newNet_1975;
wire n_35268;
wire n_10123;
wire n_42449;
wire n_41873;
wire n_37811;
wire n_25212;
wire n_9718;
wire n_11821;
wire n_10798;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_23_;
wire n_3183;
wire n_15314;
wire n_12565;
wire n_34427;
wire n_31591;
wire n_24375;
wire n_38649;
wire n_26575;
wire n_19891;
wire n_17970;
wire n_9354;
wire n_33205;
wire n_8193;
wire n_5485;
wire n_15296;
wire n_46993;
wire n_30943;
wire n_25241;
wire n_43463;
wire n_5422;
wire n_9276;
wire n_10357;
wire n_23820;
wire n_26370;
wire n_38539;
wire FE_OCP_RBN1683_n_33491;
wire n_38792;
wire n_37519;
wire newNet_1564;
wire n_2147;
wire n_37944;
wire newNet_3218;
wire n_4362;
wire n_2567;
wire newNet_538;
wire n_30550;
wire n_34204;
wire newNet_1245;
wire n_13734;
wire n_16514;
wire n_10451;
wire n_21990;
wire n_25989;
wire n_26038;
wire newNet_2673;
wire n_2025;
wire n_5534;
wire n_5959;
wire n_35522;
wire n_38047;
wire n_42101;
wire FE_OCP_RBN3577_n_4528;
wire n_20218;
wire n_38937;
wire n_19243;
wire n_1327;
wire n_3564;
wire n_8456;
wire n_25418;
wire n_43719;
wire n_17555;
wire n_35974;
wire n_11652;
wire n_40480;
wire newNet_2496;
wire FE_OCP_RBN1722_n_21004;
wire FE_OCP_RBN2587_n_9492;
wire n_34605;
wire n_42366;
wire n_22213;
wire n_8135;
wire FE_RN_1049_0;
wire n_16025;
wire n_4647;
wire n_31760;
wire n_42130;
wire n_5128;
wire newNet_2848;
wire n_20391;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_23_;
wire n_41692;
wire n_40505;
wire n_9787;
wire n_37344;
wire FE_RN_1062_0;
wire n_34420;
wire n_21335;
wire n_20220;
wire n_27921;
wire n_20798;
wire n_20357;
wire FE_RN_1485_0;
wire n_6660;
wire n_33078;
wire FE_OCP_RBN3010_n_31117;
wire n_33546;
wire n_40840;
wire n_1364;
wire n_18490;
wire n_31345;
wire n_37094;
wire newNet_2687;
wire n_14735;
wire n_37045;
wire n_5772;
wire n_4708;
wire n_24301;
wire n_15014;
wire n_5541;
wire n_17902;
wire n_24259;
wire n_72;
wire n_31833;
wire n_38583;
wire FE_OCP_RBN2834_n_39586;
wire n_28856;
wire n_35134;
wire n_1011;
wire FE_RN_739_0;
wire n_1672;
wire n_8843;
wire n_17625;
wire n_13410;
wire n_28107;
wire n_31800;
wire delay_add_ln22_unr27_stage10_stallmux_q_3_;
wire n_20582;
wire n_21543;
wire n_19446;
wire n_40113;
wire n_1514;
wire n_15182;
wire n_21541;
wire n_9693;
wire n_26730;
wire n_37028;
wire FE_RN_1820_0;
wire n_41732;
wire n_30656;
wire newNet_1928;
wire n_38386;
wire n_23903;
wire n_17780;
wire n_4608;
wire n_5243;
wire n_21954;
wire n_33111;
wire n_9747;
wire n_36396;
wire FE_RN_1014_0;
wire FE_RN_529_0;
wire n_6113;
wire n_24427;
wire n_31802;
wire n_37125;
wire n_45872;
wire newNet_3679;
wire n_19367;
wire n_40990;
wire n_2839;
wire n_32077;
wire n_14203;
wire FE_OCP_RBN2147_FE_OCPN861_n_45450;
wire n_31823;
wire n_36438;
wire n_25689;
wire n_29105;
wire n_4697;
wire n_33638;
wire n_43715;
wire n_13582;
wire n_24838;
wire newNet_2223;
wire n_38076;
wire n_9438;
wire n_10936;
wire FE_OCPN3163_n_24117;
wire n_21689;
wire FE_RN_861_0;
wire n_10330;
wire newNet_3480;
wire n_19457;
wire n_14544;
wire n_41032;
wire n_4652;
wire n_6695;
wire n_28646;
wire n_39210;
wire n_5200;
wire n_45748;
wire n_20386;
wire newNet_2448;
wire delay_add_ln22_unr8_stage4_stallmux_q_9_;
wire n_5926;
wire n_8109;
wire FE_RN_192_0;
wire n_12385;
wire n_3534;
wire n_26754;
wire beta_7;
wire newNet_2998;
wire n_4570;
wire n_38060;
wire n_27819;
wire n_39743;
wire n_40098;
wire delay_xor_ln22_unr6_stage3_stallmux_q_23_;
wire n_10152;
wire FE_OCP_RBN2606_FE_OCPN899_n_44593;
wire n_10576;
wire n_34886;
wire n_34873;
wire n_30436;
wire n_11355;
wire n_28606;
wire FE_OCPN1049_n_4459;
wire delay_add_ln22_unr2_stage2_stallmux_q_18_;
wire n_12772;
wire n_37807;
wire n_43112;
wire n_32991;
wire newNet_2612;
wire n_42520;
wire n_31233;
wire FE_RN_795_0;
wire n_36185;
wire n_22612;
wire n_23265;
wire n_40114;
wire n_1585;
wire n_1650;
wire n_1355;
wire n_38237;
wire n_5283;
wire n_32920;
wire n_31224;
wire n_13330;
wire n_34607;
wire n_6598;
wire n_10514;
wire n_24707;
wire n_22559;
wire newNet_1023;
wire FE_RN_787_0;
wire n_4180;
wire n_1045;
wire FE_OCP_RBN1208_n_16814;
wire n_11604;
wire n_36762;
wire n_46168;
wire n_12241;
wire n_42813;
wire delay_add_ln22_unr27_stage10_stallmux_q_4_;
wire n_26415;
wire FE_OCP_RBN1340_n_19077;
wire newNet_695;
wire n_40486;
wire n_30989;
wire newNet_848;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_6_;
wire FE_OCP_RBN1222_n_45522;
wire n_29640;
wire n_39798;
wire n_20560;
wire n_25319;
wire n_7965;
wire n_29527;
wire n_2766;
wire n_35231;
wire n_16306;
wire n_25368;
wire FE_OCP_RBN3661_n_15429;
wire n_40782;
wire n_39543;
wire n_36474;
wire n_45487;
wire n_894;
wire newNet_3730;
wire n_39440;
wire n_39318;
wire n_19804;
wire n_1659;
wire n_1013;
wire n_41943;
wire n_727;
wire n_42200;
wire newNet_1565;
wire n_36570;
wire n_5406;
wire n_18950;
wire newNet_504;
wire delay_add_ln22_unr14_stage6_stallmux_q_12_;
wire n_5193;
wire n_15701;
wire FE_RN_191_0;
wire n_36970;
wire newNet_1273;
wire n_20878;
wire n_20982;
wire n_10550;
wire FE_OCP_RBN2228_n_7598;
wire newNet_705;
wire FE_OCPN1757_n_33213;
wire n_21550;
wire n_32699;
wire n_39362;
wire FE_OCP_RBN3399_n_12751;
wire n_43829;
wire n_3164;
wire n_9713;
wire FE_OCP_RBN2934_n_31010;
wire n_18367;
wire delay_xor_ln21_unr15_stage6_stallmux_q_4_;
wire n_23585;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_16_;
wire FE_OCP_RBN3378_n_40716;
wire n_24598;
wire FE_OCP_RBN2304_n_7817;
wire n_11485;
wire n_26421;
wire n_37017;
wire n_4981;
wire n_10100;
wire n_42668;
wire newNet_2360;
wire n_43236;
wire n_6190;
wire n_26298;
wire n_38742;
wire n_25905;
wire n_40140;
wire n_22878;
wire n_12232;
wire n_15964;
wire newNet_2167;
wire newNet_388;
wire n_175;
wire n_5161;
wire n_41278;
wire n_9281;
wire n_16529;
wire n_8648;
wire n_7350;
wire n_27047;
wire n_39138;
wire n_7099;
wire n_30841;
wire n_2453;
wire n_46216;
wire n_16666;
wire n_22820;
wire n_43391;
wire n_20353;
wire FE_OFN830_n_2540;
wire n_33677;
wire delay_xor_ln21_unr28_stage10_stallmux_q_3_;
wire n_38371;
wire n_43384;
wire n_39754;
wire n_36156;
wire n_24484;
wire FE_OCP_DRV_N1562_n_19562;
wire n_25352;
wire n_4036;
wire n_33414;
wire n_34200;
wire n_31023;
wire newNet_3295;
wire n_3815;
wire n_5138;
wire n_25487;
wire n_38933;
wire n_32688;
wire FE_RN_1106_0;
wire n_5475;
wire FE_OCP_RBN3100_n_22502;
wire n_14622;
wire newNet_899;
wire n_3787;
wire n_37068;
wire n_2127;
wire n_8466;
wire n_19400;
wire n_15023;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_21_;
wire n_12942;
wire n_1566;
wire n_21916;
wire FE_RN_1204_0;
wire n_5674;
wire n_26883;
wire n_35672;
wire newNet_3250;
wire n_29006;
wire n_46422;
wire n_34180;
wire n_2350;
wire n_7212;
wire n_5348;
wire n_12829;
wire n_5265;
wire n_10072;
wire n_12769;
wire newNet_1243;
wire FE_RN_397_0;
wire n_22772;
wire n_2842;
wire newNet_1715;
wire FE_RN_237_0;
wire n_18773;
wire n_35955;
wire newNet_2828;
wire delay_add_ln22_unr27_stage10_stallmux_q_13_;
wire n_13676;
wire newNet_3631;
wire n_41740;
wire n_29906;
wire n_43500;
wire n_3362;
wire FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_29730;
wire newNet_1658;
wire newNet_444;
wire n_12585;
wire n_17234;
wire n_46371;
wire n_34084;
wire n_40444;
wire FE_RN_823_0;
wire n_11819;
wire n_6021;
wire newNet_1042;
wire n_6127;
wire n_1190;
wire n_21660;
wire newNet_3345;
wire n_8007;
wire n_25279;
wire n_37828;
wire n_37163;
wire n_1183;
wire newNet_2626;
wire n_16358;
wire n_1249;
wire n_7488;
wire newNet_3499;
wire n_24110;
wire n_13399;
wire n_20703;
wire newNet_407;
wire n_4643;
wire n_28713;
wire n_26179;
wire FE_OCP_RBN1993_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire n_21351;
wire n_8081;
wire n_25432;
wire n_33392;
wire n_37168;
wire n_38290;
wire FE_OFN788_n_25834;
wire FE_OCP_RBN3484_n_13667;
wire n_23918;
wire n_8143;
wire n_33449;
wire FE_OCPN1041_n_3673;
wire n_31850;
wire FE_OCP_RBN2209_n_18280;
wire n_5176;
wire n_5150;
wire n_37324;
wire n_19878;
wire n_9656;
wire FE_OCP_RBN2176_n_1864;
wire n_42749;
wire FE_RN_944_0;
wire n_7953;
wire n_39937;
wire n_38905;
wire n_27632;
wire delay_add_ln22_unr27_stage10_stallmux_q_12_;
wire newNet_1962;
wire n_10807;
wire n_41759;
wire n_36983;
wire newNet_437;
wire FE_OCP_RBN3617_n_20249;
wire n_18103;
wire n_30512;
wire n_16416;
wire n_8963;
wire n_38726;
wire newNet_243;
wire n_21724;
wire n_5706;
wire n_14246;
wire n_24802;
wire n_23324;
wire n_28379;
wire n_21424;
wire FE_OCP_DRV_N1554_n_19314;
wire n_18260;
wire n_10663;
wire FE_OCP_RBN2399_FE_RN_347_0;
wire n_45069;
wire n_6755;
wire n_17372;
wire n_41620;
wire n_17809;
wire n_8595;
wire n_34121;
wire n_34677;
wire n_33951;
wire n_2878;
wire n_35914;
wire n_37727;
wire FE_OCP_RBN1296_n_30451;
wire n_17577;
wire n_23133;
wire newNet_3287;
wire n_7242;
wire n_32502;
wire n_21486;
wire n_11627;
wire n_18647;
wire n_42414;
wire n_31010;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_26_;
wire n_40401;
wire n_42399;
wire n_6991;
wire n_26657;
wire newNet_2981;
wire n_13754;
wire n_16593;
wire n_30887;
wire n_39309;
wire n_21601;
wire n_455;
wire n_841;
wire n_5386;
wire n_34963;
wire n_9313;
wire n_5395;
wire n_19576;
wire n_11556;
wire n_22355;
wire n_5557;
wire n_19603;
wire n_37739;
wire n_23170;
wire n_8537;
wire n_19445;
wire n_21657;
wire n_10491;
wire FE_OCPN1017_n_23307;
wire n_39539;
wire n_1076;
wire n_43477;
wire n_71;
wire newNet_1473;
wire n_35277;
wire n_5142;
wire n_26705;
wire FE_OCP_RBN2887_n_10570;
wire n_19492;
wire n_30367;
wire n_8611;
wire n_33301;
wire n_5618;
wire n_41489;
wire n_11528;
wire newNet_360;
wire n_4931;
wire n_37588;
wire n_15089;
wire n_20573;
wire FE_OCP_RBN3435_n_29163;
wire n_18715;
wire n_25513;
wire n_5791;
wire n_14160;
wire n_28507;
wire n_38500;
wire delay_xor_ln21_unr6_stage3_stallmux_q_17_;
wire n_39185;
wire FE_OCP_RBN3223_n_22068;
wire n_12281;
wire newNet_462;
wire FE_RN_777_0;
wire n_20121;
wire n_2035;
wire n_19333;
wire n_11052;
wire n_3246;
wire n_40900;
wire newNet_735;
wire n_31019;
wire n_9486;
wire newNet_251;
wire n_23550;
wire n_31910;
wire n_34614;
wire n_23199;
wire n_27483;
wire n_21617;
wire n_24688;
wire n_34683;
wire FE_OCP_RBN2328_n_29378;
wire n_33490;
wire n_29837;
wire newNet_3401;
wire n_7763;
wire FE_OCP_RBN3679_n_21051;
wire n_18949;
wire n_28538;
wire n_22131;
wire n_14926;
wire n_1426;
wire n_9793;
wire n_25970;
wire FE_OCPN1054_n_14098;
wire FE_RN_1562_0;
wire FE_RN_1336_0;
wire FE_OCP_RBN2004_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_5754;
wire n_15522;
wire n_19814;
wire n_27547;
wire n_47258;
wire n_3176;
wire n_9237;
wire n_8936;
wire n_30038;
wire n_39180;
wire n_43451;
wire n_28692;
wire n_42496;
wire n_25122;
wire n_25771;
wire n_12493;
wire n_15576;
wire n_29936;
wire n_8483;
wire n_23427;
wire newNet_1586;
wire n_37863;
wire newNet_40;
wire n_31265;
wire n_34932;
wire n_3205;
wire n_39142;
wire n_4884;
wire n_1080;
wire n_23671;
wire n_21782;
wire n_28040;
wire n_33747;
wire n_21348;
wire n_32792;
wire n_7023;
wire n_10306;
wire FE_RN_281_0;
wire n_3135;
wire n_14408;
wire n_25315;
wire n_27891;
wire n_19059;
wire newNet_926;
wire n_29131;
wire n_41982;
wire n_17870;
wire n_39064;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_17_;
wire n_5318;
wire n_14661;
wire newNet_1450;
wire n_11768;
wire n_13136;
wire n_45817;
wire n_37810;
wire FE_OCP_RBN2115_n_45224;
wire n_40497;
wire n_18450;
wire n_39854;
wire n_32848;
wire n_38666;
wire n_19406;
wire n_37883;
wire n_43865;
wire n_5533;
wire FE_OCP_RBN3526_n_29624;
wire n_1709;
wire n_23105;
wire n_2734;
wire newNet_3491;
wire FE_OCP_RBN2733_n_4219;
wire n_770;
wire n_11754;
wire n_34296;
wire n_29466;
wire n_7161;
wire n_36741;
wire n_40503;
wire newNet_3504;
wire n_24061;
wire n_32479;
wire n_7343;
wire n_35968;
wire n_21819;
wire newNet_1876;
wire n_398;
wire FE_RN_161_0;
wire n_38120;
wire n_22984;
wire n_4157;
wire n_30601;
wire n_24361;
wire n_42489;
wire n_1501;
wire n_17515;
wire n_35766;
wire newNet_1522;
wire n_31113;
wire n_40522;
wire n_35841;
wire n_706;
wire n_42707;
wire n_14494;
wire n_7492;
wire newNet_2511;
wire newNet_3070;
wire n_33137;
wire FE_OCP_RBN2688_n_38870;
wire newNet_3307;
wire n_35555;
wire FE_OCP_RBN3651_n_39249;
wire FE_RN_886_0;
wire n_29404;
wire n_14986;
wire n_43510;
wire n_39276;
wire n_34801;
wire n_39705;
wire n_7858;
wire n_32621;
wire n_15809;
wire delay_add_ln22_unr14_stage6_stallmux_q_5_;
wire newNet_2906;
wire newNet_3489;
wire n_13132;
wire n_19508;
wire n_34724;
wire n_33516;
wire n_10817;
wire n_19022;
wire n_32756;
wire n_22961;
wire n_19847;
wire FE_OCP_RBN3548_n_44575;
wire n_13595;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_22_;
wire n_16899;
wire delay_xor_ln22_unr15_stage6_stallmux_q_5_;
wire n_28457;
wire newNet_1764;
wire n_33123;
wire n_27409;
wire delay_xor_ln22_unr9_stage4_stallmux_q_2_;
wire n_27007;
wire n_35540;
wire n_8263;
wire n_30184;
wire FE_OCP_RBN3578_n_8774;
wire n_47335;
wire n_20326;
wire n_7562;
wire n_25213;
wire FE_OCPN3793_n_31804;
wire n_30706;
wire n_42286;
wire n_31053;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_0_;
wire newNet_1535;
wire n_25955;
wire n_21731;
wire n_29012;
wire n_46157;
wire n_37251;
wire n_6930;
wire n_42714;
wire FE_OCP_RBN3573_n_44563;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_26_;
wire n_20442;
wire newNet_2700;
wire n_3613;
wire newNet_2109;
wire n_24922;
wire n_39406;
wire newNet_1187;
wire n_37541;
wire n_47270;
wire FE_RN_1192_0;
wire delay_xor_ln21_unr28_stage10_stallmux_q_0_;
wire n_41072;
wire n_3241;
wire n_7733;
wire n_43583;
wire newNet_2547;
wire n_911;
wire n_39664;
wire n_33082;
wire n_47177;
wire n_3689;
wire n_20751;
wire n_9333;
wire n_16916;
wire newNet_2177;
wire n_20250;
wire n_21965;
wire FE_RN_1358_0;
wire FE_OCP_RBN1709_n_22150;
wire newNet_1600;
wire n_36589;
wire n_32767;
wire newNet_347;
wire n_6920;
wire n_21738;
wire n_4721;
wire FE_OCPN861_n_45450;
wire n_3358;
wire n_11332;
wire n_23358;
wire n_24791;
wire newNet_2028;
wire n_41636;
wire n_9385;
wire n_22767;
wire n_10078;
wire n_18343;
wire n_10758;
wire newNet_2000;
wire n_959;
wire n_26216;
wire n_33711;
wire n_15060;
wire n_32550;
wire n_33759;
wire n_37306;
wire n_41274;
wire n_3884;
wire n_43503;
wire n_23698;
wire n_7379;
wire newNet_578;
wire n_17251;
wire n_42100;
wire n_11707;
wire n_10913;
wire n_22176;
wire n_4856;
wire FE_RN_1689_0;
wire n_31497;
wire delay_add_ln22_unr8_stage4_stallmux_q_22_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_12_;
wire n_8557;
wire n_877;
wire newNet_3165;
wire n_10505;
wire n_16221;
wire FE_RN_622_0;
wire n_1302;
wire n_38251;
wire n_31099;
wire n_4005;
wire n_323;
wire n_41082;
wire n_12761;
wire n_7531;
wire FE_RN_13_0;
wire newNet_336;
wire n_39425;
wire n_18095;
wire n_27975;
wire n_25272;
wire n_6656;
wire n_32645;
wire n_5147;
wire FE_OCP_RBN2613_n_9075;
wire n_7000;
wire n_18612;
wire n_36062;
wire n_40701;
wire newNet_1466;
wire newNet_3348;
wire newNet_297;
wire n_18524;
wire n_5822;
wire n_15058;
wire n_5672;
wire n_6260;
wire n_39941;
wire delay_add_ln22_unr20_stage8_stallmux_q_11_;
wire n_2149;
wire n_3079;
wire n_35783;
wire n_37500;
wire n_11980;
wire n_37135;
wire newNet_3717;
wire n_10537;
wire n_17443;
wire n_23999;
wire n_14024;
wire n_13210;
wire n_6089;
wire n_22752;
wire n_46949;
wire FE_RN_868_0;
wire FE_OCP_RBN2637_n_38806;
wire n_38106;
wire n_8650;
wire n_5263;
wire n_41287;
wire n_1482;
wire n_22180;
wire n_33361;
wire n_44102;
wire n_36343;
wire n_22339;
wire FE_OCP_RBN2769_n_9892;
wire n_37096;
wire n_6542;
wire n_38306;
wire n_27854;
wire n_37218;
wire n_18591;
wire n_32936;
wire n_18008;
wire n_15473;
wire n_7229;
wire n_31693;
wire n_246;
wire n_47247;
wire FE_RN_700_0;
wire n_20003;
wire newNet_3129;
wire newNet_2010;
wire n_26581;
wire n_8995;
wire n_24984;
wire newNet_1803;
wire n_17649;
wire n_22706;
wire n_27462;
wire n_14694;
wire FE_OCP_RBN1213_n_31847;
wire n_38344;
wire n_693;
wire n_34022;
wire n_32671;
wire n_18924;
wire n_14346;
wire n_15879;
wire n_27957;
wire n_38957;
wire n_18320;
wire FE_OCP_RBN3447_n_37945;
wire n_9759;
wire n_40982;
wire newNet_2651;
wire n_7944;
wire n_34871;
wire n_43682;
wire n_8841;
wire n_26552;
wire n_33252;
wire n_35900;
wire n_944;
wire n_37769;
wire n_24619;
wire n_5210;
wire n_287;
wire n_20957;
wire n_17213;
wire newNet_321;
wire n_24892;
wire n_14439;
wire n_7905;
wire n_43346;
wire n_43871;
wire n_41662;
wire n_1949;
wire n_22737;
wire newNet_539;
wire n_35196;
wire n_9009;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_26_;
wire n_38604;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_30_;
wire n_9565;
wire newNet_3523;
wire n_20477;
wire n_13778;
wire n_5379;
wire n_8409;
wire n_31154;
wire n_6070;
wire n_36353;
wire n_21811;
wire n_26588;
wire n_3193;
wire n_461;
wire n_25625;
wire n_40941;
wire FE_OCP_RBN2700_n_4238;
wire n_24915;
wire n_29247;
wire n_15256;
wire newNet_1316;
wire n_41444;
wire n_10475;
wire n_7123;
wire n_33705;
wire FE_RN_409_0;
wire n_40524;
wire n_43038;
wire n_3091;
wire n_33219;
wire n_40179;
wire newNet_2418;
wire n_22058;
wire newNet_1821;
wire n_34516;
wire n_43522;
wire n_9163;
wire n_25055;
wire n_20653;
wire n_11195;
wire n_2024;
wire n_42587;
wire FE_OCP_RBN3136_n_32380;
wire n_14365;
wire n_18248;
wire n_2625;
wire n_3007;
wire newNet_2696;
wire n_37950;
wire n_34635;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_11_;
wire n_22234;
wire n_21163;
wire n_12080;
wire newNet_835;
wire n_5501;
wire n_10497;
wire n_1620;
wire n_29775;
wire n_2768;
wire n_5418;
wire n_31687;
wire n_27194;
wire n_20115;
wire n_20249;
wire n_22813;
wire n_24754;
wire n_6731;
wire n_31756;
wire n_2739;
wire n_46941;
wire n_42602;
wire n_4277;
wire n_31504;
wire n_21494;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_17_;
wire n_9504;
wire n_7466;
wire FE_RN_1037_0;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_30_;
wire n_43593;
wire n_36924;
wire n_10510;
wire n_10715;
wire n_1407;
wire n_24066;
wire FE_RN_1771_0;
wire n_4704;
wire n_14367;
wire n_28116;
wire newNet_2949;
wire n_18704;
wire n_5589;
wire FE_OCP_RBN3585_n_25295;
wire n_32126;
wire n_4405;
wire n_35380;
wire newNet_1843;
wire newNet_1214;
wire n_24562;
wire n_43541;
wire n_130;
wire n_35709;
wire newNet_176;
wire newNet_2324;
wire n_38145;
wire n_2606;
wire FE_RN_240_0;
wire n_3142;
wire n_17635;
wire FE_OCP_RBN3601_FE_OCPN1243_n_44460;
wire n_21634;
wire n_36628;
wire newNet_2537;
wire n_29588;
wire newNet_812;
wire n_22261;
wire n_27146;
wire n_9032;
wire n_5352;
wire n_934;
wire n_12695;
wire n_34435;
wire n_6985;
wire n_33996;
wire n_1922;
wire newNet_531;
wire n_818;
wire n_31810;
wire n_16846;
wire n_13034;
wire n_40534;
wire n_2852;
wire n_17001;
wire n_1;
wire n_10483;
wire n_17875;
wire n_20151;
wire n_35689;
wire n_32143;
wire n_27582;
wire n_5408;
wire n_5850;
wire n_4425;
wire n_29760;
wire n_38433;
wire n_9481;
wire n_12860;
wire n_39103;
wire n_33207;
wire n_22947;
wire newNet_2709;
wire n_7270;
wire newNet_2355;
wire n_27178;
wire FE_OCP_RBN3412_n_2100;
wire n_21407;
wire n_5274;
wire n_4809;
wire n_23052;
wire n_17103;
wire newNet_1176;
wire n_11007;
wire n_21116;
wire n_29103;
wire n_10989;
wire newNet_718;
wire newNet_417;
wire n_14789;
wire n_38832;
wire n_23118;
wire n_18769;
wire n_13689;
wire n_23711;
wire n_32158;
wire n_28804;
wire n_41255;
wire n_5665;
wire n_11590;
wire n_38402;
wire n_46055;
wire n_28597;
wire n_18994;
wire n_39808;
wire newNet_3725;
wire n_5898;
wire n_34644;
wire n_33802;
wire newNet_851;
wire FE_RN_967_0;
wire n_36891;
wire n_7589;
wire n_33578;
wire n_29160;
wire n_27313;
wire n_6705;
wire newNet_170;
wire n_29750;
wire n_13295;
wire n_4553;
wire n_33627;
wire n_34710;
wire n_37063;
wire n_32034;
wire n_18856;
wire n_26462;
wire n_2795;
wire n_23994;
wire n_3969;
wire n_27882;
wire n_37050;
wire n_40816;
wire n_23362;
wire n_2086;
wire n_31349;
wire FE_OCP_RBN3624_n_38870;
wire n_24359;
wire n_22889;
wire n_35450;
wire n_13973;
wire delay_add_ln22_unr20_stage8_stallmux_q_0_;
wire FE_RN_1187_0;
wire n_14473;
wire n_40742;
wire newNet_2761;
wire n_5460;
wire n_33014;
wire n_35041;
wire n_26040;
wire n_5512;
wire n_37521;
wire n_20273;
wire n_13024;
wire n_36771;
wire n_2745;
wire n_11203;
wire n_24901;
wire n_22144;
wire n_14891;
wire newNet_57;
wire newNet_1992;
wire newNet_76;
wire n_6143;
wire n_40066;
wire n_32085;
wire FE_RN_109_0;
wire n_13370;
wire n_24548;
wire n_42288;
wire n_29796;
wire delay_add_ln22_unr23_stage9_stallmux_q_25_;
wire n_82;
wire n_14427;
wire n_23653;
wire n_14811;
wire n_23458;
wire n_16626;
wire n_21331;
wire n_34928;
wire newNet_2375;
wire FE_RN_877_0;
wire n_5439;
wire n_39341;
wire FE_OCP_RBN1151_n_13460;
wire n_27139;
wire n_15221;
wire n_24493;
wire n_25748;
wire n_26902;
wire n_18514;
wire n_43562;
wire n_3753;
wire n_2214;
wire n_20735;
wire newNet_1745;
wire n_22993;
wire delay_xor_ln21_unr6_stage3_stallmux_q_20_;
wire n_12469;
wire n_24151;
wire n_38617;
wire n_20291;
wire n_30196;
wire n_22800;
wire n_22934;
wire n_12236;
wire n_8622;
wire n_39625;
wire n_27806;
wire n_20037;
wire FE_OCPN1454_n_18559;
wire n_9721;
wire n_29158;
wire n_43108;
wire n_47002;
wire n_1157;
wire n_5784;
wire n_13691;
wire FE_OCP_DRV_N1571_n_29860;
wire delay_add_ln22_unr2_stage2_stallmux_q_8_;
wire n_19746;
wire n_34100;
wire FE_RN_146_0;
wire n_14703;
wire n_32362;
wire n_17992;
wire n_43095;
wire n_12300;
wire n_40431;
wire n_8605;
wire FE_OCP_RBN2155_n_1602;
wire n_6405;
wire n_31848;
wire n_25405;
wire n_21699;
wire n_24994;
wire FE_OCP_RBN2910_n_26394;
wire n_31612;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_20_;
wire n_28843;
wire n_1371;
wire n_4525;
wire n_41357;
wire FE_OCP_DRV_N1549_n_19053;
wire newNet_2055;
wire n_25023;
wire n_33196;
wire FE_OCPN901_n_44593;
wire n_31468;
wire n_13141;
wire n_301;
wire newNet_785;
wire n_10162;
wire n_39978;
wire n_7821;
wire n_19559;
wire n_36428;
wire n_22739;
wire newNet_275;
wire n_25703;
wire n_23410;
wire n_32205;
wire n_21939;
wire n_30290;
wire n_31353;
wire n_41027;
wire n_16237;
wire n_22964;
wire n_30509;
wire n_35629;
wire n_30674;
wire n_16409;
wire newNet_1503;
wire n_20462;
wire n_34666;
wire FE_OCP_RBN2594_n_25181;
wire n_24502;
wire n_14049;
wire n_31410;
wire n_7687;
wire n_17099;
wire n_10623;
wire FE_RN_445_0;
wire n_23596;
wire n_24404;
wire FE_OCP_RBN3437_n_33750;
wire n_31330;
wire n_39713;
wire n_21266;
wire n_12297;
wire n_5653;
wire n_8208;
wire delay_xor_ln22_unr28_stage10_stallmux_q_3_;
wire n_43891;
wire n_13603;
wire n_26990;
wire n_21173;
wire n_4318;
wire n_11260;
wire n_33257;
wire n_11318;
wire n_32316;
wire n_3001;
wire n_24098;
wire n_38654;
wire newNet_2022;
wire n_18174;
wire n_24397;
wire n_16976;
wire n_34860;
wire FE_RN_169_0;
wire n_42856;
wire n_20059;
wire n_30147;
wire n_34972;
wire n_15309;
wire n_41815;
wire n_25915;
wire newNet_1164;
wire n_28343;
wire n_16460;
wire n_7989;
wire n_41545;
wire n_22406;
wire n_26743;
wire n_31394;
wire n_13312;
wire n_1115;
wire n_38109;
wire n_42148;
wire n_35478;
wire n_15775;
wire n_28881;
wire n_41992;
wire n_37479;
wire n_29808;
wire n_5215;
wire n_18569;
wire n_22450;
wire n_30962;
wire n_11871;
wire FE_RN_1794_0;
wire n_7370;
wire n_29909;
wire FE_OCPN1385_n_470;
wire n_32975;
wire n_24806;
wire n_32222;
wire n_16429;
wire n_31101;
wire n_901;
wire n_40124;
wire n_41578;
wire n_6473;
wire n_43050;
wire n_39520;
wire n_20620;
wire n_32613;
wire n_37539;
wire n_12856;
wire n_7626;
wire n_24606;
wire n_40685;
wire n_40239;
wire n_18781;
wire n_19611;
wire n_10253;
wire n_18757;
wire n_32778;
wire n_11159;
wire n_33275;
wire n_3388;
wire n_6844;
wire n_11091;
wire n_11453;
wire n_30918;
wire n_29226;
wire n_6213;
wire n_29145;
wire n_33893;
wire newNet_114;
wire n_41527;
wire n_35615;
wire n_31322;
wire n_15861;
wire FE_OCPN1034_n_28420;
wire newNet_1553;
wire n_672;
wire n_22694;
wire newNet_2311;
wire n_42874;
wire n_3104;
wire n_4339;
wire n_34065;
wire FE_OCP_RBN2262_n_33691;
wire n_38479;
wire FE_OCP_RBN2365_n_24372;
wire newNet_2878;
wire n_4597;
wire n_860;
wire n_6392;
wire n_564;
wire n_28708;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_21_;
wire n_7220;
wire n_41727;
wire n_740;
wire n_44180;
wire newNet_209;
wire newNet_131;
wire n_37172;
wire n_19735;
wire n_43751;
wire n_31855;
wire n_29371;
wire n_14386;
wire n_12935;
wire n_23547;
wire n_30040;
wire n_30200;
wire n_40549;
wire newNet_3079;
wire n_964;
wire n_614;
wire FE_RN_408_0;
wire n_17741;
wire n_10426;
wire n_42011;
wire n_25982;
wire n_343;
wire n_24971;
wire n_35402;
wire n_44052;
wire newNet_1699;
wire n_39569;
wire n_10855;
wire n_22140;
wire n_10659;
wire n_10742;
wire n_22839;
wire n_26638;
wire n_22295;
wire n_31715;
wire n_42847;
wire n_16095;
wire n_31433;
wire n_26863;
wire n_36941;
wire n_14722;
wire newNet_1100;
wire n_33611;
wire n_10175;
wire n_36878;
wire newNet_3277;
wire n_43461;
wire n_42751;
wire newNet_2966;
wire n_1770;
wire n_10569;
wire n_41580;
wire newNet_2043;
wire n_28196;
wire n_29286;
wire n_33979;
wire n_35737;
wire n_36455;
wire n_39218;
wire n_28468;
wire n_4392;
wire n_28285;
wire newNet_3314;
wire n_25188;
wire FE_OCP_RBN3618_n_14841;
wire n_10732;
wire n_17752;
wire FE_OCPN1406_n_25859;
wire n_25205;
wire n_15240;
wire n_9201;
wire n_43365;
wire n_30703;
wire newNet_218;
wire n_12485;
wire n_30846;
wire n_5992;
wire n_1095;
wire n_2485;
wire n_21001;
wire FE_OCP_RBN3684_FE_RN_770_0;
wire n_21236;
wire n_36674;
wire n_35322;
wire n_26893;
wire n_41614;
wire n_24075;
wire n_2665;
wire n_28847;
wire FE_OCPN935_n_42192;
wire n_18414;
wire n_38565;
wire n_34162;
wire n_13453;
wire FE_OCP_RBN3652_n_10100;
wire n_25562;
wire n_11546;
wire n_11761;
wire n_4557;
wire n_29561;
wire n_36501;
wire n_22464;
wire FE_OCP_RBN3416_n_12739;
wire n_20434;
wire FE_RN_549_0;
wire n_1141;
wire n_23952;
wire n_43186;
wire newNet_38;
wire n_28328;
wire n_15585;
wire n_3128;
wire FE_RN_345_0;
wire n_34353;
wire newNet_2443;
wire newNet_985;
wire n_7035;
wire n_15340;
wire n_19427;
wire n_8445;
wire n_22204;
wire n_2457;
wire n_26612;
wire n_41560;
wire FE_RN_1549_0;
wire n_34891;
wire n_27992;
wire n_34333;
wire n_35240;
wire n_318;
wire n_41251;
wire FE_OCP_RBN2178_n_33022;
wire n_16819;
wire n_808;
wire n_34995;
wire n_26737;
wire n_3100;
wire n_29032;
wire n_38924;
wire n_27319;
wire n_2569;
wire n_25014;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_27_;
wire n_43322;
wire n_557;
wire n_22311;
wire n_10171;
wire n_28218;
wire n_17434;
wire newNet_1109;
wire newNet_3324;
wire n_31201;
wire FE_OCP_RBN3207_n_44365;
wire n_42402;
wire n_34598;
wire n_32734;
wire n_15545;
wire FE_OCP_RBN2939_n_26276;
wire newNet_3557;
wire newNet_2684;
wire n_13291;
wire n_5816;
wire n_35299;
wire n_40939;
wire newNet_801;
wire n_36127;
wire n_13886;
wire n_16490;
wire FE_OCPN1496_n_26528;
wire n_11585;
wire n_24716;
wire n_30482;
wire n_27118;
wire n_13426;
wire n_6204;
wire n_10810;
wire newNet_3672;
wire n_36239;
wire n_38220;
wire n_12465;
wire n_4167;
wire n_34655;
wire n_38184;
wire FE_RN_1866_0;
wire n_42052;
wire n_19511;
wire n_3569;
wire n_32868;
wire FE_OCP_RBN3209_n_44365;
wire n_20468;
wire n_47255;
wire FE_RN_1276_0;
wire n_25344;
wire n_26451;
wire n_37142;
wire n_24998;
wire n_36374;
wire n_10203;
wire n_26360;
wire n_41178;
wire n_21149;
wire n_31290;
wire n_10166;
wire n_26378;
wire n_10192;
wire n_27392;
wire n_22550;
wire n_25124;
wire n_25428;
wire n_24954;
wire FE_OCPN959_n_3951;
wire n_19337;
wire n_36485;
wire n_22968;
wire n_21393;
wire n_20675;
wire n_29754;
wire n_11943;
wire n_8097;
wire n_20753;
wire n_11499;
wire newNet_1676;
wire newNet_714;
wire n_35349;
wire n_29163;
wire delay_add_ln22_unr8_stage4_stallmux_q_0_;
wire n_12709;
wire FE_RN_1532_0;
wire n_8666;
wire n_26815;
wire n_26184;
wire n_43910;
wire n_30791;
wire n_14035;
wire n_44028;
wire n_15898;
wire n_42899;
wire n_36207;
wire n_12593;
wire FE_OCPN3767_n_14439;
wire n_16100;
wire n_37575;
wire newNet_1425;
wire n_10135;
wire n_22363;
wire n_794;
wire n_5718;
wire n_6916;
wire n_1406;
wire n_25393;
wire n_38445;
wire n_20821;
wire n_17607;
wire n_1824;
wire n_41393;
wire n_18254;
wire n_29149;
wire n_35935;
wire n_29913;
wire n_16924;
wire n_4975;
wire n_21150;
wire n_31769;
wire n_41763;
wire n_19607;
wire n_41983;
wire n_30630;
wire n_35503;
wire newNet_2102;
wire n_14294;
wire FE_RN_54_0;
wire n_896;
wire n_18411;
wire newNet_3752;
wire FE_RN_952_0;
wire n_16517;
wire n_21667;
wire n_16124;
wire n_11013;
wire n_41337;
wire n_3210;
wire newNet_1393;
wire n_25950;
wire n_41242;
wire n_8767;
wire n_38387;
wire sin_out_11;
wire n_14115;
wire n_5442;
wire n_16658;
wire n_19689;
wire n_9817;
wire n_9544;
wire n_29818;
wire n_27509;
wire n_44690;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_2_;
wire n_13586;
wire n_26856;
wire n_5355;
wire n_41502;
wire n_8212;
wire n_16013;
wire n_27603;
wire n_35985;
wire n_7976;
wire FE_OCP_RBN3534_n_13765;
wire FE_RN_1793_0;
wire n_2398;
wire n_37072;
wire n_17611;
wire n_31448;
wire n_18538;
wire n_17948;
wire newNet_3609;
wire n_12378;
wire n_36682;
wire n_37833;
wire n_32312;
wire n_6066;
wire n_24323;
wire newNet_1337;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_2_;
wire n_17429;
wire FE_OCP_RBN3663_n_20750;
wire n_24602;
wire FE_OCP_RBN3404_n_28597;
wire n_9516;
wire n_28990;
wire newNet_2211;
wire n_21858;
wire n_9971;
wire n_11773;
wire n_40417;
wire newNet_429;
wire n_7147;
wire n_13417;
wire n_22797;
wire n_36909;
wire newNet_1970;
wire FE_RN_475_0;
wire n_40046;
wire newNet_2915;
wire FE_RN_257_0;
wire newNet_527;
wire newNet_1775;
wire n_7086;
wire n_1199;
wire n_5940;
wire n_13735;
wire n_37821;
wire n_2257;
wire n_8824;
wire n_13663;
wire n_15997;
wire delay_add_ln22_unr14_stage6_stallmux_q_9_;
wire n_23827;
wire n_23529;
wire n_33541;
wire n_10736;
wire n_2729;
wire n_18798;
wire n_31261;
wire n_18018;
wire n_19729;
wire n_28476;
wire n_35474;
wire n_39598;
wire FE_OCP_DRV_N3159_n_31303;
wire n_38315;
wire delay_xor_ln22_unr6_stage3_stallmux_q_1_;
wire FE_OCP_RBN2427_n_19599;
wire newNet_2724;
wire n_43351;
wire n_1854;
wire n_42070;
wire n_24053;
wire newNet_3034;
wire n_38768;
wire n_1687;
wire FE_OCPN1407_n_672;
wire n_2028;
wire n_6676;
wire n_7726;
wire n_4674;
wire n_13286;
wire n_31342;
wire newNet_1792;
wire n_34211;
wire newNet_2476;
wire FE_RN_1813_0;
wire n_13377;
wire n_35833;
wire n_33769;
wire n_10809;
wire n_33667;
wire n_2448;
wire n_709;
wire n_10524;
wire n_24344;
wire n_14738;
wire n_864;
wire newNet_1623;
wire n_38800;
wire n_5343;
wire n_28810;
wire n_18129;
wire n_15156;
wire n_744;
wire n_30572;
wire n_25734;
wire n_27829;
wire n_25753;
wire n_17914;
wire n_6783;
wire FE_RN_1762_0;
wire n_32741;
wire delay_add_ln22_unr14_stage6_stallmux_q_21_;
wire n_6270;
wire FE_OCP_RBN3676_n_21039;
wire delay_add_ln22_unr5_stage3_stallmux_q_30_;
wire n_19780;
wire n_14287;
wire n_39994;
wire FE_OCP_RBN3645_n_44490;
wire n_31326;
wire n_40592;
wire n_42426;
wire n_30899;
wire n_638;
wire n_18737;
wire cos_out_30;
wire n_29281;
wire n_34541;
wire n_22718;
wire n_29343;
wire n_9128;
wire n_2067;
wire n_12193;
wire n_17989;
wire n_25295;
wire n_45311;
wire n_18371;
wire n_26578;
wire n_28569;
wire FE_OFN4_n_43918;
wire n_24857;
wire n_32233;
wire n_3037;
wire n_26637;
wire n_102;
wire n_31859;
wire n_7040;
wire delay_add_ln22_unr27_stage10_stallmux_q_1_;
wire n_42396;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_23_;
wire n_22483;
wire n_39139;
wire n_11784;
wire n_22583;
wire n_32907;
wire FE_RN_74_0;
wire n_2511;
wire n_9591;
wire n_9931;
wire n_26984;
wire FE_OCP_RBN3021_n_39942;
wire FE_RN_1647_0;
wire n_16329;
wire n_39470;
wire n_37489;
wire n_10401;
wire n_13988;
wire n_42152;
wire n_24062;
wire FE_OCP_RBN3454_FE_OCPN1240_n_7721;
wire n_12869;
wire n_26067;
wire n_39060;
wire n_40132;
wire n_22952;
wire n_32786;
wire n_30448;
wire n_38340;
wire n_25983;
wire n_43507;
wire n_42624;
wire n_15800;
wire n_23298;
wire n_29661;
wire n_39386;
wire FE_RN_1248_0;
wire n_15925;
wire n_9289;
wire n_3695;
wire n_12439;
wire n_16489;
wire n_316;
wire n_16063;
wire n_22622;
wire newNet_3098;
wire n_35098;
wire n_30223;
wire newNet_378;
wire n_23848;
wire n_25307;
wire n_15286;
wire n_3850;
wire n_37699;
wire n_20425;
wire newNet_2667;
wire FE_RN_613_0;
wire n_19575;
wire FE_RN_253_0;
wire n_40891;
wire n_28349;
wire n_36732;
wire newNet_3330;
wire newNet_3581;
wire n_3255;
wire n_40465;
wire n_29473;
wire n_39587;
wire n_29742;
wire n_18653;
wire n_37794;
wire n_40674;
wire n_31092;
wire n_30381;
wire n_32336;
wire n_34821;
wire n_12348;
wire FE_RN_1350_0;
wire newNet_373;
wire FE_OCP_RBN3855_n_21224;
wire n_24586;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_25_;
wire n_8332;
wire n_26979;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_27_;
wire n_6556;
wire n_19682;
wire n_5480;
wire newNet_3063;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_15_;
wire newNet_1293;
wire FE_OCP_RBN3064_n_22170;
wire n_40293;
wire n_17403;
wire n_28603;
wire n_33885;
wire n_12725;
wire n_36972;
wire FE_OCP_RBN2839_n_4692;
wire n_41812;
wire n_2874;
wire n_45120;
wire n_2495;
wire n_24769;
wire n_7382;
wire n_35198;
wire n_11523;
wire n_7785;
wire n_36980;
wire n_36694;
wire n_17502;
wire n_28383;
wire FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_32981;
wire FE_RN_912_0;
wire n_24877;
wire n_35679;
wire n_42947;
wire n_4387;
wire n_19309;
wire n_38248;
wire n_44071;
wire newNet_2465;
wire n_11403;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_3_;
wire n_19489;
wire FE_RN_955_0;
wire n_9138;
wire n_35211;
wire n_10329;
wire n_12149;
wire newNet_105;
wire n_21379;
wire FE_RN_1137_0;
wire n_28099;
wire delay_add_ln22_unr20_stage8_stallmux_q_25_;
wire n_38512;
wire n_17765;
wire n_6438;
wire newNet_2171;
wire n_767;
wire n_12647;
wire n_31277;
wire n_13556;
wire n_31999;
wire n_21637;
wire n_21822;
wire n_32506;
wire n_34329;
wire n_12255;
wire n_43630;
wire n_5569;
wire n_11081;
wire n_17964;
wire n_25052;
wire n_11657;
wire n_14491;
wire n_5523;
wire newNet_129;
wire n_33145;
wire n_1945;
wire n_11696;
wire n_27190;
wire n_905;
wire n_45896;
wire n_33194;
wire n_34740;
wire FE_RN_1865_0;
wire n_28827;
wire newNet_1124;
wire n_3546;
wire delay_xor_ln22_unr28_stage10_stallmux_q_2_;
wire n_33631;
wire n_12902;
wire newNet_351;
wire n_37919;
wire n_33299;
wire n_9398;
wire FE_OCPN1800_FE_OFN780_n_17093;
wire n_22608;
wire n_27802;
wire newNet_3590;
wire n_25105;
wire n_7478;
wire n_40438;
wire n_17879;
wire n_31883;
wire n_17692;
wire n_36797;
wire n_12084;
wire n_25856;
wire n_3327;
wire n_7103;
wire n_17042;
wire n_38005;
wire n_15917;
wire n_2991;
wire n_45312;
wire n_26661;
wire n_11033;
wire newNet_1867;
wire n_31881;
wire n_29594;
wire n_23568;
wire n_33268;
wire n_36713;
wire FE_OCPN1389_n_9220;
wire n_29955;
wire n_38041;
wire FE_OCPN3165_n_44267;
wire n_21431;
wire n_10418;
wire n_36038;
wire n_17292;
wire n_41380;
wire n_3452;
wire n_23390;
wire n_9496;
wire n_10264;
wire FE_RN_843_0;
wire FE_OCP_RBN2888_n_46957;
wire n_31546;
wire n_36963;
wire n_19540;
wire n_20914;
wire n_38287;
wire FE_RN_611_0;
wire n_9966;
wire FE_OCP_RBN2199_n_2032;
wire n_23480;
wire newNet_1632;
wire newNet_246;
wire n_23127;
wire n_20796;
wire n_8700;
wire n_11490;
wire n_40600;
wire n_34114;
wire FE_RN_1129_0;
wire n_10650;
wire n_32123;
wire n_32941;
wire n_25385;
wire n_28548;
wire n_6269;
wire n_15757;
wire n_29241;
wire n_33701;
wire n_22659;
wire n_5771;
wire n_18632;
wire n_3314;
wire n_16850;
wire n_11836;
wire n_38129;
wire n_1845;
wire n_38992;
wire n_16113;
wire n_13011;
wire n_33329;
wire n_6152;
wire n_25873;
wire n_41370;
wire n_24081;
wire n_27398;
wire newNet_759;
wire n_23767;
wire n_28667;
wire newNet_3509;
wire n_41953;
wire n_14676;
wire n_40856;
wire newNet_383;
wire n_26461;
wire n_4476;
wire n_18886;
wire n_26947;
wire FE_RN_917_0;
wire n_6326;
wire n_13785;
wire n_9887;
wire n_19861;
wire n_33237;
wire n_38507;
wire n_34263;
wire n_41110;
wire n_46368;
wire n_2303;
wire n_15226;
wire n_836;
wire n_13798;
wire n_2381;
wire n_41929;
wire n_30824;
wire n_37389;
wire newNet_3479;
wire n_27079;
wire n_29485;
wire n_40252;
wire n_9682;
wire FE_OCP_RBN3482_n_13667;
wire n_24801;
wire newNet_2351;
wire newNet_3175;
wire n_576;
wire n_14534;
wire n_16219;
wire n_7701;
wire n_35304;
wire n_27165;
wire n_41752;
wire n_10556;
wire n_32889;
wire n_10449;
wire newNet_3428;
wire newNet_110;
wire FE_OCPN1037_n_28318;
wire n_13365;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_4_;
wire n_41551;
wire n_2194;
wire n_25707;
wire n_18269;
wire n_5660;
wire n_29041;
wire n_35786;
wire n_17539;
wire n_33508;
wire n_41828;
wire n_15481;
wire n_17215;
wire n_36614;
wire n_19771;
wire n_17591;
wire n_823;
wire newNet_1356;
wire n_7266;
wire n_41716;
wire FE_OCP_RBN2346_n_29448;
wire n_1440;
wire n_14575;
wire n_28031;
wire n_29322;
wire n_44144;
wire n_4438;
wire n_7234;
wire n_27934;
wire FE_RN_1050_0;
wire n_41433;
wire n_35317;
wire n_24759;
wire FE_OCP_RBN2461_n_14273;
wire n_22727;
wire n_38353;
wire n_498;
wire n_11552;
wire n_25608;
wire n_19238;
wire n_28311;
wire newNet_3201;
wire n_46426;
wire n_34238;
wire newNet_2646;
wire newNet_634;
wire n_14626;
wire FE_OCPN1450_n_20443;
wire n_44360;
wire n_18766;
wire n_8074;
wire n_13226;
wire n_41891;
wire n_35680;
wire n_4483;
wire n_13503;
wire n_24478;
wire n_7137;
wire n_36788;
wire newNet_46;
wire n_32326;
wire n_15810;
wire FE_OCP_RBN2504_n_13896;
wire newNet_3628;
wire n_5844;
wire n_11342;
wire n_40490;
wire n_1401;
wire n_205;
wire n_38232;
wire n_5835;
wire FE_OCP_RBN3116_n_22710;
wire delay_xor_ln22_unr3_stage2_stallmux_q_23_;
wire newNet_1727;
wire n_11550;
wire n_231;
wire n_13051;
wire n_18046;
wire n_12683;
wire n_19349;
wire n_43414;
wire n_5146;
wire newNet_2959;
wire newNet_2882;
wire n_19194;
wire FE_OCP_RBN2945_FE_RN_1269_0;
wire n_16770;
wire n_40478;
wire n_17279;
wire n_35867;
wire n_11739;
wire n_10908;
wire n_25633;
wire newNet_2953;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_2_;
wire n_11518;
wire n_21913;
wire n_41162;
wire n_41201;
wire FE_OCPN1414_n_19715;
wire FE_OCP_RBN2161_n_40687;
wire newNet_2303;
wire n_35039;
wire n_28576;
wire n_28910;
wire n_29532;
wire FE_OCP_RBN1352_n_19148;
wire n_43902;
wire n_36514;
wire n_31861;
wire n_24182;
wire n_16082;
wire n_18356;
wire n_16274;
wire n_47279;
wire FE_RN_298_0;
wire n_14038;
wire newNet_1654;
wire n_9146;
wire n_8633;
wire n_32540;
wire n_427;
wire n_12043;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_4_;
wire n_32724;
wire n_11269;
wire n_33353;
wire n_26827;
wire n_39258;
wire n_27225;
wire n_31365;
wire n_9841;
wire n_11623;
wire newNet_228;
wire n_14262;
wire n_20050;
wire n_8506;
wire newNet_1857;
wire n_31704;
wire n_3239;
wire n_47266;
wire n_27457;
wire n_27479;
wire n_36075;
wire n_18204;
wire n_18291;
wire n_5880;
wire n_27691;
wire n_19076;
wire n_5679;
wire n_29866;
wire FE_RN_1045_0;
wire n_6183;
wire n_25005;
wire n_30649;
wire n_28588;
wire FE_OCP_RBN3718_n_39913;
wire n_3085;
wire n_21519;
wire n_35593;
wire FE_OCPN1766_n_33447;
wire n_14338;
wire n_22351;
wire n_8659;
wire n_7255;
wire n_18695;
wire n_5632;
wire n_28373;
wire n_23152;
wire n_6225;
wire n_41042;
wire n_13870;
wire n_35150;
wire n_37990;
wire n_20513;
wire n_26916;
wire n_24270;
wire n_31555;
wire newNet_181;
wire n_28728;
wire n_11172;
wire n_46936;
wire n_23088;
wire n_4041;
wire n_29575;
wire FE_RN_90_0;
wire n_41085;
wire n_33937;
wire n_299;
wire FE_RN_320_0;
wire FE_OCP_RBN3635_n_47260;
wire n_16246;
wire n_32484;
wire newNet_1447;
wire n_15064;
wire n_32559;
wire n_15399;
wire n_32260;
wire n_33651;
wire n_27844;
wire n_31163;
wire n_10279;
wire n_22647;
wire FE_OCP_RBN3088_FE_OCPN1052_n_31674;
wire newNet_288;
wire n_19501;
wire n_4617;
wire n_31689;
wire n_42537;
wire n_21802;
wire n_2296;
wire n_20502;
wire n_43703;
wire newNet_2373;
wire n_42794;
wire cos_out_16;
wire FE_OCPN3773_n_15371;
wire n_5079;
wire n_8804;
wire n_43705;
wire n_43672;
wire n_41993;
wire newNet_1894;
wire n_8040;
wire n_34610;
wire n_5336;
wire n_14645;
wire n_41884;
wire n_24728;
wire FE_RN_1193_0;
wire n_37965;
wire n_33452;
wire n_23557;
wire n_16714;
wire n_23096;
wire n_44575;
wire n_2168;
wire delay_xor_ln21_unr15_stage6_stallmux_q_0_;
wire n_885;
wire n_29049;
wire n_7150;
wire n_18168;
wire n_38637;
wire n_39944;
wire n_10285;
wire n_41870;
wire n_14684;
wire n_8111;
wire n_38967;
wire n_10107;
wire n_26989;
wire n_22381;
wire n_19401;
wire n_30623;
wire n_16371;
wire n_40362;
wire n_29059;
wire n_29768;
wire n_1041;
wire n_24819;
wire n_39201;
wire delay_add_ln22_unr8_stage4_stallmux_q_20_;
wire n_33820;
wire n_8846;
wire n_30903;
wire n_40567;
wire n_13682;
wire FE_OCP_RBN3384_n_33108;
wire newNet_1441;
wire n_38897;
wire n_6513;
wire n_42889;
wire newNet_3527;
wire n_12366;
wire newNet_3690;
wire n_40019;
wire FE_OCP_RBN2177_n_1864;
wire n_38485;
wire n_39694;
wire newNet_2937;
wire n_3994;
wire n_9245;
wire n_37717;
wire n_17800;
wire FE_OCPN1405_n_25859;
wire FE_OCP_RBN2531_n_38693;
wire n_20281;
wire FE_OCPUNCON3143_n_19138;
wire n_36134;
wire n_17864;
wire n_36811;
wire n_3439;
wire n_16032;
wire n_34251;
wire FE_OCP_RBN2276_n_24077;
wire n_14540;
wire n_23210;
wire n_33352;
wire FE_RN_1658_0;
wire n_20626;
wire newNet_2113;
wire n_22575;
wire n_32947;
wire n_36801;
wire n_5922;
wire n_7336;
wire n_5508;
wire n_3475;
wire n_28685;
wire delay_xor_ln22_unr3_stage2_stallmux_q_3_;
wire n_6602;
wire n_24930;
wire n_39906;
wire n_6341;
wire n_17414;
wire n_36932;
wire newNet_452;
wire n_40860;
wire delay_add_ln22_unr2_stage2_stallmux_q_27_;
wire n_2967;
wire n_14015;
wire n_12533;
wire n_20194;
wire n_6357;
wire FE_RN_1376_0;
wire n_40724;
wire FE_OCPN1762_n_37877;
wire n_9784;
wire n_40957;
wire n_9833;
wire n_10456;
wire n_23073;
wire newNet_613;
wire n_40324;
wire newNet_2890;
wire n_9737;
wire newNet_2543;
wire n_28264;
wire n_3956;
wire n_38134;
wire n_29501;
wire n_1938;
wire delay_add_ln22_unr2_stage2_stallmux_q_6_;
wire n_16140;
wire n_32832;
wire n_35691;
wire n_32918;
wire newNet_3151;
wire newNet_574;
wire newNet_2733;
wire n_9575;
wire n_16544;
wire n_39447;
wire n_10216;
wire newNet_1688;
wire n_36652;
wire n_3899;
wire n_42738;
wire n_40734;
wire n_25150;
wire n_869;
wire n_6716;
wire n_32495;
wire n_16891;
wire newNet_749;
wire n_35971;
wire FE_OCP_DRV_N1572_n_29860;
wire n_13006;
wire n_3384;
wire n_47240;
wire n_4082;
wire n_15906;
wire newNet_2462;
wire n_42224;
wire newNet_1046;
wire n_6016;
wire n_28800;
wire newNet_2268;
wire n_36141;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_27_;
wire n_40278;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_12_;
wire newNet_1133;
wire n_9639;
wire FE_OCP_RBN2725_n_4219;
wire n_35774;
wire newNet_1707;
wire FE_OCPN1508_n_23414;
wire n_43623;
wire n_36361;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_29_;
wire n_2001;
wire n_40964;
wire n_8172;
wire FE_RN_1760_0;
wire n_12749;
wire FE_OCP_RBN2293_n_2438;
wire n_23294;
wire n_28893;
wire newNet_2409;
wire n_3996;
wire n_33907;
wire n_33426;
wire n_8761;
wire n_31405;
wire n_1735;
wire n_40749;
wire n_45192;
wire n_42797;
wire n_18575;
wire n_36956;
wire newNet_1921;
wire n_31974;
wire delay_xor_ln21_unr21_stage8_stallmux_q_9_;
wire n_40154;
wire n_21867;
wire n_34878;
wire n_41923;
wire n_41325;
wire n_21757;
wire n_23093;
wire n_11313;
wire n_2273;
wire FE_OCPN1029_n_28423;
wire n_23137;
wire n_5938;
wire n_17762;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire n_20785;
wire n_15767;
wire n_31623;
wire n_33972;
wire n_35739;
wire newNet_1909;
wire n_11000;
wire FE_OCPN1495_n_26528;
wire newNet_1605;
wire n_3265;
wire n_5629;
wire n_6171;
wire n_28926;
wire n_31311;
wire newNet_2439;
wire n_515;
wire n_26054;
wire n_10111;
wire n_11106;
wire n_36902;
wire n_40610;
wire n_2631;
wire n_33740;
wire n_19838;
wire n_16396;
wire n_17073;
wire n_24780;
wire n_2265;
wire n_41418;
wire n_38393;
wire n_36409;
wire n_38862;
wire n_3911;
wire n_36849;
wire n_37941;
wire n_30553;
wire FE_OCP_RBN2520_n_8762;
wire n_7929;
wire n_26449;
wire n_30372;
wire n_14117;
wire newNet_3182;
wire n_26319;
wire n_1117;
wire n_25974;
wire n_19381;
wire FE_OCP_RBN2608_n_3807;
wire newNet_1698;
wire newNet_1286;
wire n_1491;
wire newNet_2616;
wire newNet_67;
wire n_14090;
wire n_40540;
wire FE_RN_1304_0;
wire n_2752;
wire newNet_2136;
wire n_3344;
wire n_28629;
wire n_17363;
wire n_17893;
wire n_19994;
wire n_20363;
wire newNet_2579;
wire n_7011;
wire FE_RN_1864_0;
wire n_22786;
wire n_33494;
wire FE_RN_643_0;
wire FE_OCP_RBN2550_n_44944;
wire n_29707;
wire newNet_548;
wire n_12619;
wire n_25651;
wire n_22361;
wire n_40622;
wire n_13048;
wire n_22874;
wire FE_OCP_RBN2891_n_10568;
wire n_15626;
wire n_22671;
wire n_30337;
wire newNet_2422;
wire n_13401;
wire n_27711;
wire n_27988;
wire n_30490;
wire newNet_3560;
wire newNet_3604;
wire n_44223;
wire n_20944;
wire n_32275;
wire n_24290;
wire n_12843;
wire FE_OCP_RBN2526_n_3421;
wire n_18138;
wire n_6504;
wire n_27997;
wire n_39647;
wire n_30295;
wire n_9609;
wire n_32229;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_31_;
wire n_1762;
wire n_17009;
wire n_22988;
wire newNet_2444;
wire n_18862;
wire n_17135;
wire n_12260;
wire n_16748;
wire n_23054;
wire n_37040;
wire newNet_1987;
wire n_26205;
wire n_40926;
wire n_25999;
wire FE_OCPN1011_n_7802;
wire n_3590;
wire FE_RN_205_0;
wire n_33040;
wire n_87;
wire n_3302;
wire newNet_153;
wire n_26527;
wire n_36498;
wire n_2684;
wire n_43799;
wire n_6701;
wire n_28052;
wire n_174;
wire n_7571;
wire n_26518;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_13_;
wire n_5121;
wire n_4191;
wire FE_OCP_RBN2713_n_14982;
wire n_19888;
wire n_28120;
wire n_14755;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_12_;
wire n_39329;
wire n_28141;
wire n_25223;
wire newNet_1756;
wire FE_RN_1116_0;
wire n_28011;
wire n_7170;
wire n_26606;
wire FE_OCP_RBN3680_n_10338;
wire n_19570;
wire n_14852;
wire n_2011;
wire n_11181;
wire n_36854;
wire n_30442;
wire n_8326;
wire n_14131;
wire n_35951;
wire n_15842;
wire n_36740;
wire n_40380;
wire newNet_1942;
wire n_13763;
wire n_46337;
wire FE_RN_1732_0;
wire n_13390;
wire n_23632;
wire n_6094;
wire n_42000;
wire FE_RN_775_0;
wire n_4800;
wire n_5553;
wire n_8348;
wire delay_add_ln22_unr2_stage2_stallmux_q_16_;
wire n_41520;
wire n_8426;
wire n_29833;
wire n_38461;
wire n_40388;
wire n_9640;
wire n_3526;
wire n_28958;
wire n_38731;
wire n_38375;
wire n_13727;
wire n_15774;
wire FE_OCPN1388_n_11041;
wire n_39708;
wire n_40754;
wire n_9648;
wire n_35254;
wire n_5325;
wire n_14757;
wire newNet_1572;
wire FE_OCP_RBN1191_n_14911;
wire n_43192;
wire n_7116;
wire n_30345;
wire n_37858;
wire n_10377;
wire n_15957;
wire n_10979;
wire newNet_2127;
wire n_35423;
wire FE_OCP_RBN2338_n_24325;
wire n_11285;
wire n_33442;
wire n_1733;
wire n_28940;
wire n_2430;
wire n_9360;
wire n_37193;
wire n_7360;
wire n_31149;
wire n_39043;
wire n_36274;
wire n_29895;
wire n_1679;
wire n_5801;
wire n_34042;
wire n_2954;
wire FE_OCP_RBN2893_n_26152;
wire n_908;
wire n_30106;
wire n_10840;
wire n_39652;
wire FE_OCPN911_n_43022;
wire n_17724;
wire n_16730;
wire n_3122;
wire n_3367;
wire n_9856;
wire n_29943;
wire n_7502;
wire n_18483;
wire n_9669;
wire n_20727;
wire n_20687;
wire n_42388;
wire n_42215;
wire n_23498;
wire n_45323;
wire n_39818;
wire n_13815;
wire n_15171;
wire n_28897;
wire n_41039;
wire n_4216;
wire n_37470;
wire n_26191;
wire n_28181;
wire n_7544;
wire n_9415;
wire n_1837;
wire newNet_2988;
wire n_36900;
wire n_11663;
wire n_993;
wire n_11915;
wire n_38382;
wire newNet_1091;
wire n_21192;
wire n_22059;
wire n_41295;
wire n_34275;
wire n_13631;
wire n_9822;
wire FE_RN_805_0;
wire n_39514;
wire n_36258;
wire FE_OCPN1499_n_26125;
wire newNet_3276;
wire n_24383;
wire n_3954;
wire n_32512;
wire n_1800;
wire n_38901;
wire n_15687;
wire n_22922;
wire FE_OCP_RBN3474_n_7886;
wire n_43466;
wire beta_20;
wire n_11532;
wire n_31897;
wire n_21227;
wire n_23865;
wire n_25321;
wire n_28290;
wire n_34581;
wire n_31605;
wire n_25328;
wire FE_RN_1808_0;
wire n_21330;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_24_;
wire n_41448;
wire n_42260;
wire n_7193;
wire n_15734;
wire FE_RN_969_0;
wire n_24687;
wire FE_OCP_RBN2586_n_9009;
wire n_26974;
wire FE_OCP_RBN3129_n_32266;
wire n_20681;
wire n_829;
wire n_33097;
wire n_11129;
wire FE_RN_865_0;
wire n_37507;
wire n_16157;
wire n_44804;
wire n_4685;
wire n_732;
wire n_28585;
wire n_20890;
wire newNet_199;
wire n_21544;
wire newNet_1374;
wire n_41908;
wire n_34840;
wire FE_OCP_RBN3483_n_13667;
wire n_40315;
wire n_13041;
wire n_25259;
wire n_1636;
wire n_20797;
wire newNet_1862;
wire n_7841;
wire n_35078;
wire n_21610;
wire n_39279;
wire n_22601;
wire n_43426;
wire n_34463;
wire n_14809;
wire n_21154;
wire n_16341;
wire n_32367;
wire n_27704;
wire n_5127;
wire n_3877;
wire n_19354;
wire n_37466;
wire n_12374;
wire FE_RN_1683_0;
wire n_5017;
wire n_5971;
wire n_13525;
wire n_33171;
wire n_7303;
wire n_12992;
wire n_19262;
wire n_24831;
wire n_43580;
wire n_36725;
wire newNet_1645;
wire n_12750;
wire n_25604;
wire n_9168;
wire newNet_2069;
wire n_10367;
wire n_32843;
wire FE_OCP_RBN3818_n_44061;
wire newNet_1084;
wire n_8374;
wire n_21529;
wire n_43694;
wire n_12495;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_7_;
wire n_22967;
wire n_33411;
wire n_24535;
wire n_15569;
wire n_11365;
wire n_34293;
wire n_35740;
wire n_23611;
wire n_34907;
wire n_34218;
wire n_16948;
wire n_28331;
wire n_34935;
wire n_43737;
wire n_3338;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_31_;
wire n_15085;
wire n_35274;
wire n_4283;
wire n_41939;
wire n_33104;
wire n_24165;
wire newNet_365;
wire n_372;
wire n_28300;
wire n_37681;
wire n_1673;
wire FE_OCP_RBN3667_n_20812;
wire n_16179;
wire n_28206;
wire n_14101;
wire n_40873;
wire n_26546;
wire n_10571;
wire n_26504;
wire FE_OCP_RBN2491_n_3338;
wire n_43483;
wire n_2181;
wire newNet_2094;
wire FE_OCP_RBN3495_n_19390;
wire FE_RN_1675_0;
wire n_11275;
wire n_26064;
wire n_8944;
wire n_4470;
wire n_2650;
wire FE_OCP_RBN2007_n_45209;
wire n_6009;
wire n_20596;
wire n_6759;
wire n_20988;
wire n_36461;
wire n_18683;
wire newNet_260;
wire n_1107;
wire n_38490;
wire n_29651;
wire FE_RN_434_0;
wire n_24040;
wire FE_RN_881_0;
wire newNet_2006;
wire n_14163;
wire n_20044;
wire FE_OCP_RBN2570_n_29922;
wire n_41598;
wire n_43868;
wire n_26941;
wire n_46150;
wire n_13572;
wire n_10297;
wire n_13343;
wire n_42081;
wire n_18813;
wire n_35035;
wire n_42321;
wire n_42348;
wire n_11893;
wire FE_OCP_RBN3436_n_29163;
wire n_42871;
wire n_383;
wire n_33605;
wire FE_OCP_RBN2308_n_29298;
wire n_45065;
wire n_44309;
wire n_34729;
wire newNet_2458;
wire n_35017;
wire delay_xor_ln21_unr3_stage2_stallmux_q_17_;
wire n_9883;
wire n_34534;
wire n_7960;
wire n_9310;
wire n_14371;
wire n_46358;
wire n_38453;
wire n_6804;
wire n_34641;
wire n_15525;
wire n_19648;
wire n_32255;
wire n_15137;
wire n_32620;
wire n_18890;
wire newNet_790;
wire newNet_3046;
wire n_31375;
wire n_32963;
wire n_11968;
wire FE_OCPN1863_n_26171;
wire FE_RN_654_0;
wire n_11362;
wire n_23753;
wire FE_OCPN1789_n_18119;
wire newNet_3629;
wire n_40794;
wire n_21104;
wire n_19116;
wire n_40905;
wire n_17850;
wire n_37374;
wire n_7165;
wire FE_OCP_RBN2900_n_44853;
wire delay_add_ln22_unr8_stage4_stallmux_q_30_;
wire n_33394;
wire n_30284;
wire n_34791;
wire n_4493;
wire n_34053;
wire n_17718;
wire n_32215;
wire n_24340;
wire newNet_2813;
wire n_41139;
wire FE_RN_1285_0;
wire FE_RN_1417_0;
wire n_19602;
wire n_9987;
wire n_22693;
wire n_39562;
wire n_9080;
wire n_43041;
wire n_33635;
wire n_40877;
wire n_44034;
wire n_17086;
wire n_5021;
wire n_28368;
wire newNet_3399;
wire n_13544;
wire n_23008;
wire newNet_2361;
wire n_13598;
wire n_27310;
wire n_33366;
wire FE_OCP_RBN2720_n_9494;
wire n_11992;
wire n_42781;
wire n_12343;
wire n_17928;
wire n_23929;
wire n_24099;
wire n_11613;
wire n_20517;
wire n_2740;
wire n_13606;
wire n_25216;
wire n_19469;
wire n_22060;
wire n_33847;
wire FE_RN_1318_0;
wire n_1063;
wire n_13261;
wire n_29326;
wire n_17872;
wire n_33128;
wire n_15770;
wire n_23108;
wire n_30920;
wire n_9770;
wire FE_RN_830_0;
wire n_20224;
wire newNet_1222;
wire n_27903;
wire n_36212;
wire n_26076;
wire n_37296;
wire n_39247;
wire n_41634;
wire n_10735;
wire newNet_106;
wire FE_OCP_RBN3677_n_21051;
wire n_24269;
wire n_21384;
wire delay_xor_ln22_unr9_stage4_stallmux_q_3_;
wire n_20375;
wire FE_OCPN3760_n_2466;
wire n_28820;
wire n_16413;
wire n_40894;
wire n_10864;
wire n_3909;
wire n_743;
wire n_10019;
wire n_2922;
wire n_20334;
wire n_18236;
wire FE_OCP_RBN2344_FE_OCPN870_n_2737;
wire n_36477;
wire n_28176;
wire n_43640;
wire FE_OCP_RBN2673_n_14991;
wire n_15929;
wire FE_OCP_RBN2786_n_15079;
wire n_7290;
wire FE_RN_1505_0;
wire n_31043;
wire n_7338;
wire n_2284;
wire n_33274;
wire n_17475;
wire n_10727;
wire n_13468;
wire newNet_3688;
wire n_5574;
wire n_39669;
wire n_30675;
wire n_6870;
wire n_20126;
wire n_36897;
wire FE_OCPN898_n_44776;
wire n_3966;
wire n_24364;
wire n_46383;
wire n_41899;
wire n_11954;
wire n_27415;
wire n_25673;
wire n_10926;
wire n_29227;
wire n_3596;
wire n_11139;
wire n_20312;
wire n_5622;
wire FE_OCP_RBN2281_n_29111;
wire n_30016;
wire n_35872;
wire n_45484;
wire FE_OCP_RBN3644_n_44490;
wire n_24972;
wire n_29872;
wire n_38468;
wire newNet_1190;
wire FE_OCP_RBN2810_n_15433;
wire n_31864;
wire n_24285;
wire n_43377;
wire n_2771;
wire n_28494;
wire FE_OCPN1420_n_14003;
wire newNet_602;
wire n_5605;
wire delay_xor_ln22_unr21_stage8_stallmux_q_7_;
wire newNet_2584;
wire FE_OFN831_n_19807;
wire newNet_3646;
wire delay_add_ln22_unr27_stage10_stallmux_q_18_;
wire newNet_2023;
wire n_13016;
wire newNet_1568;
wire newNet_3544;
wire newNet_1439;
wire n_1959;
wire n_7440;
wire n_8531;
wire n_19142;
wire n_23933;
wire n_22038;
wire n_29596;
wire n_29463;
wire n_4070;
wire n_1081;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_5_;
wire n_925;
wire n_25348;
wire n_17542;
wire n_20290;
wire delay_xor_ln21_unr3_stage2_stallmux_q_22_;
wire n_419;
wire newNet_3305;
wire n_27042;
wire n_34349;
wire n_34368;
wire n_36640;
wire n_6154;
wire n_1878;
wire n_6218;
wire FE_OCP_RBN2267_n_2430;
wire n_38413;
wire n_18074;
wire n_38837;
wire n_20931;
wire n_35550;
wire newNet_3054;
wire newNet_2874;
wire newNet_3662;
wire n_18968;
wire FE_OCP_RBN2806_n_30643;
wire n_2958;
wire n_32612;
wire n_35487;
wire newNet_448;
wire n_32780;
wire n_50;
wire n_37520;
wire newNet_3538;
wire n_27816;
wire n_22301;
wire n_3519;
wire n_16313;
wire n_10821;
wire FE_OCP_RBN3822_n_44061;
wire n_22216;
wire n_40506;
wire n_26970;
wire n_13679;
wire n_21248;
wire FE_OCP_RBN2432_n_14018;
wire n_14030;
wire n_20236;
wire n_5186;
wire n_188;
wire n_18744;
wire n_843;
wire n_31467;
wire n_15967;
wire newNet_162;
wire n_7807;
wire n_4586;
wire n_3103;
wire n_5961;
wire n_38780;
wire n_47205;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_31_;
wire n_2543;
wire n_5919;
wire n_7454;
wire FE_OCP_RBN2354_n_13858;
wire n_8292;
wire FE_OCP_RBN3376_n_6822;
wire n_24300;
wire n_25712;
wire n_3890;
wire FE_RN_1110_0;
wire n_13179;
wire cos_out_4;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_1_;
wire n_31356;
wire n_8056;
wire n_16047;
wire FE_OCP_RBN1906_n_29080;
wire n_7062;
wire n_31819;
wire n_41960;
wire n_20010;
wire n_36340;
wire n_40663;
wire n_33052;
wire n_35898;
wire n_13649;
wire FE_OCP_RBN3369_n_32436;
wire n_37379;
wire n_13761;
wire n_1695;
wire n_4688;
wire FE_OCP_RBN2347_n_29448;
wire n_6832;
wire n_41143;
wire n_30992;
wire n_20734;
wire n_19779;
wire n_38921;
wire n_36739;
wire n_3943;
wire n_26166;
wire n_39950;
wire n_6118;
wire n_4154;
wire n_12419;
wire newNet_3078;
wire n_31385;
wire n_43014;
wire n_11053;
wire n_31236;
wire n_4111;
wire delay_xor_ln21_unr21_stage8_stallmux_q_7_;
wire n_33976;
wire FE_RN_959_0;
wire newNet_2560;
wire FE_OCP_RBN2265_n_29033;
wire n_42583;
wire n_15830;
wire n_30341;
wire FE_RN_110_0;
wire newNet_3746;
wire n_41000;
wire n_11841;
wire n_17583;
wire n_18050;
wire n_19807;
wire n_304;
wire n_38295;
wire n_45873;
wire FE_RN_617_0;
wire newNet_3505;
wire n_27729;
wire n_41409;
wire FE_OCP_RBN3023_n_39942;
wire n_26723;
wire FE_OCPN1464_n_29630;
wire newNet_2568;
wire n_3070;
wire n_1549;
wire n_35072;
wire n_8457;
wire n_35234;
wire n_8369;
wire n_26037;
wire n_12945;
wire newNet_2429;
wire n_17903;
wire n_8933;
wire n_13511;
wire n_16448;
wire n_42557;
wire n_31498;
wire n_33446;
wire n_42474;
wire n_18640;
wire newNet_3376;
wire n_12166;
wire n_28964;
wire n_39601;
wire n_4547;
wire n_15796;
wire n_18549;
wire n_45753;
wire newNet_1096;
wire n_9327;
wire n_14200;
wire n_34738;
wire n_44068;
wire newNet_1248;
wire n_14135;
wire n_42868;
wire newNet_943;
wire n_12060;
wire FE_RN_1568_0;
wire n_12920;
wire n_35250;
wire n_12926;
wire n_25181;
wire n_34487;
wire n_26161;
wire n_32653;
wire n_11412;
wire n_29901;
wire n_17620;
wire n_41061;
wire n_43231;
wire n_39027;
wire FE_RN_202_0;
wire n_44262;
wire newNet_1028;
wire n_3202;
wire n_30776;
wire n_31246;
wire newNet_3061;
wire n_30116;
wire n_37250;
wire n_27193;
wire n_8227;
wire n_891;
wire n_9655;
wire n_20545;
wire n_40695;
wire FE_OCP_DRV_N3743_n_25400;
wire n_37012;
wire n_20124;
wire n_23617;
wire newNet_2252;
wire n_6350;
wire delay_add_ln22_unr20_stage8_stallmux_q_30_;
wire n_15603;
wire n_16026;
wire n_3216;
wire delay_add_ln22_unr17_stage7_stallmux_q_16_;
wire n_5232;
wire n_10411;
wire n_32796;
wire n_37173;
wire FE_RN_1074_0;
wire n_7861;
wire n_43221;
wire n_25902;
wire n_8573;
wire n_13847;
wire n_25025;
wire n_42373;
wire n_17056;
wire n_31522;
wire FE_OCP_RBN3591_n_14704;
wire n_17967;
wire n_5450;
wire FE_RN_1449_0;
wire newNet_3183;
wire n_33762;
wire n_33880;
wire n_1120;
wire n_47016;
wire newNet_516;
wire n_3022;
wire n_7143;
wire FE_OCPN1797_n_20333;
wire n_20420;
wire n_17452;
wire n_32319;
wire newNet_1058;
wire n_17812;
wire n_13088;
wire n_23196;
wire n_6880;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_0_;
wire FE_OCP_DRV_N3168_FE_RN_1789_0;
wire n_16829;
wire n_25931;
wire n_32593;
wire n_18553;
wire FE_OCP_RBN2224_n_12902;
wire n_99;
wire n_10658;
wire n_21041;
wire n_19310;
wire n_37339;
wire n_35186;
wire n_1542;
wire n_27993;
wire n_12879;
wire n_26702;
wire n_27004;
wire n_6040;
wire n_17753;
wire newNet_20;
wire n_15573;
wire n_28356;
wire n_2675;
wire n_30693;
wire n_17804;
wire n_18;
wire n_6631;
wire n_15414;
wire n_16038;
wire n_37773;
wire n_29234;
wire n_21789;
wire FE_OCPN3184_n_22294;
wire newNet_986;
wire newNet_501;
wire n_36672;
wire n_21863;
wire n_40557;
wire n_25535;
wire n_41457;
wire n_29780;
wire n_16905;
wire newNet_2917;
wire n_43822;
wire n_5447;
wire n_19480;
wire n_3030;
wire newNet_3233;
wire n_35164;
wire FE_OCP_RBN2923_n_5130;
wire n_14397;
wire n_11639;
wire n_25034;
wire n_26697;
wire n_22349;
wire n_6925;
wire mux_while_ln12_psv_q_2_;
wire n_31501;
wire n_36690;
wire n_42807;
wire n_37766;
wire FE_OCP_DRV_N1565_n_28654;
wire n_12716;
wire newNet_2654;
wire n_23140;
wire newNet_3494;
wire n_3533;
wire n_17744;
wire n_22926;
wire n_33706;
wire n_32381;
wire n_23963;
wire n_35138;
wire n_31289;
wire n_37411;
wire n_34308;
wire n_9226;
wire n_26777;
wire n_30130;
wire n_21093;
wire n_8132;
wire n_28617;
wire n_34374;
wire newNet_43;
wire n_22331;
wire n_7612;
wire n_33387;
wire delay_xor_ln21_unr3_stage2_stallmux_q_6_;
wire n_45627;
wire n_43135;
wire n_32355;
wire n_2605;
wire newNet_2669;
wire n_25276;
wire n_7654;
wire n_25129;
wire n_41195;
wire n_2450;
wire n_13394;
wire n_38523;
wire FE_OCP_RBN3657_n_15314;
wire n_2444;
wire n_3194;
wire newNet_1150;
wire n_11480;
wire delay_xor_ln22_unr9_stage4_stallmux_q_10_;
wire n_9353;
wire n_19665;
wire newNet_3291;
wire delay_xor_ln21_unr9_stage4_stallmux_q_0_;
wire FE_OCP_RBN2006_n_45209;
wire newNet_2234;
wire n_26597;
wire n_39729;
wire n_15210;
wire newNet_2757;
wire n_2371;
wire n_12388;
wire FE_OCP_RBN3402_n_28597;
wire newNet_3212;
wire n_38168;
wire n_18066;
wire n_42236;
wire n_3112;
wire n_30037;
wire n_29908;
wire n_28268;
wire n_2515;
wire n_16579;
wire n_33204;
wire n_33157;
wire n_6896;
wire n_21080;
wire newNet_1779;
wire n_5308;
wire n_7824;
wire n_18170;
wire n_9369;
wire n_17890;
wire n_30515;
wire n_12967;
wire delay_add_ln22_unr5_stage3_stallmux_q_3_;
wire n_2828;
wire n_29204;
wire n_14653;
wire n_27887;
wire n_28398;
wire n_4820;
wire n_3627;
wire newNet_3618;
wire FE_OCP_RBN1132_n_12827;
wire n_44454;
wire n_37594;
wire n_38983;
wire n_12569;
wire n_28339;
wire n_33474;
wire FE_OCP_RBN2493_n_8508;
wire n_6849;
wire n_28094;
wire n_42756;
wire n_9443;
wire n_24528;
wire n_13995;
wire n_5229;
wire delay_add_ln22_unr14_stage6_stallmux_q_19_;
wire n_28888;
wire n_17997;
wire n_8838;
wire n_3964;
wire FE_RN_1196_0;
wire FE_OCP_RBN1715_n_20734;
wire n_31613;
wire n_18627;
wire n_28370;
wire n_1565;
wire n_15946;
wire n_43037;
wire newNet_2663;
wire n_10442;
wire n_38698;
wire FE_OCP_DRV_N3167_FE_RN_1789_0;
wire n_23489;
wire newNet_1014;
wire n_23114;
wire n_2616;
wire FE_OCP_RBN1355_n_44259;
wire FE_RN_1871_0;
wire n_7366;
wire FE_RN_1789_0;
wire n_11527;
wire n_1718;
wire n_32060;
wire FE_OCP_RBN1136_n_17040;
wire n_26634;
wire n_29064;
wire newNet_201;
wire n_37401;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_9_;
wire n_1152;
wire n_30878;
wire n_31317;
wire n_12106;
wire n_25337;
wire n_27620;
wire n_26514;
wire n_16556;
wire n_18278;
wire n_6302;
wire n_23801;
wire n_29542;
wire n_39621;
wire n_27383;
wire newNet_2710;
wire FE_RN_1280_0;
wire n_38383;
wire n_13537;
wire n_46219;
wire n_20383;
wire n_36976;
wire n_22453;
wire n_15243;
wire n_20634;
wire FE_OCP_RBN3528_n_13765;
wire n_5562;
wire n_19963;
wire n_29703;
wire n_41933;
wire n_7760;
wire FE_RN_1241_0;
wire n_37039;
wire newNet_2348;
wire n_4578;
wire n_35455;
wire n_34697;
wire n_4901;
wire FE_RN_1472_0;
wire n_23652;
wire n_9474;
wire n_30173;
wire n_4453;
wire n_39013;
wire FE_RN_12_0;
wire n_5110;
wire n_41309;
wire n_23455;
wire newNet_2984;
wire n_38721;
wire n_12392;
wire n_40015;
wire n_29995;
wire n_37722;
wire n_36776;
wire n_35960;
wire n_7886;
wire n_21763;
wire n_34830;
wire n_34289;
wire n_46234;
wire newNet_958;
wire n_31826;
wire FE_RN_958_0;
wire n_27669;
wire n_34021;
wire n_35310;
wire n_17035;
wire FE_OCP_RBN3392_n_37557;
wire n_9524;
wire n_11626;
wire n_35439;
wire n_3423;
wire n_24173;
wire n_34688;
wire n_43747;
wire n_41156;
wire n_7052;
wire n_9433;
wire n_10804;
wire n_42932;
wire n_13630;
wire n_23812;
wire n_26381;
wire newNet_3585;
wire n_7582;
wire n_19188;
wire n_7243;
wire n_22390;
wire newNet_856;
wire n_22274;
wire n_13164;
wire n_10778;
wire n_43750;
wire n_18213;
wire n_14341;
wire n_22898;
wire FE_RN_1669_0;
wire n_28426;
wire n_4629;
wire n_38612;
wire n_34478;
wire n_25668;
wire newNet_1613;
wire n_35711;
wire n_41387;
wire n_37922;
wire n_2716;
wire n_14511;
wire n_22708;
wire newNet_1074;
wire n_14551;
wire newNet_3380;
wire n_11259;
wire n_31116;
wire n_15847;
wire n_17596;
wire n_8259;
wire n_17711;
wire n_38503;
wire FE_RN_1067_0;
wire n_21602;
wire n_8541;
wire n_2082;
wire n_11317;
wire n_20406;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_28_;
wire n_36452;
wire n_8305;
wire n_29667;
wire n_16236;
wire n_42076;
wire n_1975;
wire n_27773;
wire FE_OCP_RBN1689_n_18986;
wire n_37868;
wire n_45617;
wire n_28291;
wire newNet_639;
wire n_36946;
wire n_36488;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_1_;
wire n_38496;
wire FE_OCP_RBN3523_n_8242;
wire n_12267;
wire FE_OCP_RBN3568_n_29857;
wire n_12311;
wire n_2913;
wire n_20251;
wire n_235;
wire n_9789;
wire n_31714;
wire n_36994;
wire n_28805;
wire newNet_2053;
wire newNet_2636;
wire n_16158;
wire n_20302;
wire n_751;
wire n_30860;
wire n_42337;
wire n_41912;
wire n_30195;
wire n_36582;
wire n_643;
wire FE_RN_1108_0;
wire n_2867;
wire n_39739;
wire n_85;
wire n_30000;
wire n_12919;
wire n_1398;
wire n_40706;
wire n_7523;
wire n_27278;
wire n_19616;
wire n_9196;
wire n_27432;
wire n_2472;
wire n_39415;
wire n_3540;
wire n_24522;
wire n_27199;
wire n_5951;
wire n_4057;
wire n_10337;
wire delay_xor_ln22_unr3_stage2_stallmux_q_1_;
wire n_22978;
wire n_34661;
wire n_2161;
wire n_32882;
wire FE_OCP_RBN1354_n_33584;
wire n_22554;
wire n_34948;
wire n_40257;
wire n_23150;
wire FE_RN_1263_0;
wire n_20461;
wire n_3502;
wire newNet_3432;
wire n_28058;
wire FE_OCP_RBN3309_n_44722;
wire n_35640;
wire n_4851;
wire n_14816;
wire n_34008;
wire n_10360;
wire n_12932;
wire n_30211;
wire n_42759;
wire n_16604;
wire FE_OCP_RBN2868_n_16088;
wire n_39897;
wire n_9264;
wire n_22699;
wire n_7130;
wire newNet_3228;
wire n_26616;
wire n_7223;
wire n_22632;
wire n_11542;
wire n_6957;
wire n_21029;
wire n_37607;
wire newNet_1748;
wire newNet_2078;
wire newNet_555;
wire n_15563;
wire newNet_54;
wire FE_OCP_RBN1154_n_18375;
wire newNet_1167;
wire FE_RN_1377_0;
wire n_10620;
wire n_26930;
wire n_34348;
wire n_35626;
wire n_38806;
wire n_33891;
wire n_25302;
wire n_15142;
wire newNet_208;
wire newNet_1345;
wire n_16451;
wire n_23608;
wire n_14148;
wire n_39645;
wire n_1255;
wire n_37117;
wire newNet_1692;
wire n_36331;
wire n_1212;
wire n_39281;
wire newNet_2417;
wire n_3148;
wire n_13121;
wire n_20900;
wire n_30915;
wire n_30683;
wire n_43433;
wire n_39872;
wire FE_OCPN1022_n_23195;
wire n_26436;
wire n_29826;
wire n_29805;
wire n_36552;
wire n_37124;
wire n_33642;
wire n_26009;
wire FE_OCPN1240_n_7721;
wire n_20356;
wire FE_OCP_RBN2495_n_8641;
wire n_41822;
wire n_1450;
wire n_39917;
wire n_29608;
wire n_37309;
wire n_37083;
wire n_7209;
wire newNet_1767;
wire n_446;
wire newNet_2283;
wire n_10425;
wire n_23599;
wire n_16938;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_30_;
wire n_24881;
wire n_3586;
wire n_4529;
wire n_39435;
wire n_41906;
wire n_42093;
wire n_27919;
wire n_33376;
wire n_9583;
wire n_41022;
wire n_4000;
wire n_2208;
wire n_23795;
wire sin_out_8;
wire n_26714;
wire n_8106;
wire n_30023;
wire n_20295;
wire n_39844;
wire n_7916;
wire n_4420;
wire FE_OCP_RBN3643_n_44490;
wire n_1662;
wire n_37909;
wire FE_RN_1298_0;
wire n_9686;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_18_;
wire n_36268;
wire n_22424;
wire n_25828;
wire n_5832;
wire newNet_223;
wire n_2563;
wire n_40599;
wire n_19248;
wire n_6103;
wire n_42538;
wire newNet_2940;
wire n_37955;
wire n_32813;
wire n_19597;
wire n_39862;
wire n_26100;
wire FE_OCPN3180_FE_OCP_RBN2744_n_15319;
wire n_18284;
wire n_36065;
wire n_17247;
wire n_25164;
wire n_16255;
wire n_15862;
wire n_47264;
wire n_37958;
wire n_19330;
wire n_6609;
wire n_19952;
wire n_9562;
wire n_7999;
wire n_4962;
wire n_10373;
wire n_38546;
wire n_20565;
wire n_29186;
wire n_31911;
wire n_33723;
wire n_23995;
wire n_13317;
wire n_2929;
wire n_38919;
wire FE_OCP_RBN1912_n_20965;
wire n_42447;
wire n_10984;
wire n_28387;
wire n_21345;
wire n_31108;
wire n_30378;
wire n_4090;
wire FE_OCP_RBN2559_n_44576;
wire n_33733;
wire n_40578;
wire n_4950;
wire n_26411;
wire newNet_2178;
wire newNet_1433;
wire n_9807;
wire n_15360;
wire n_2942;
wire n_18114;
wire FE_RN_1069_0;
wire n_14960;
wire n_25114;
wire n_41818;
wire n_25318;
wire newNet_3522;
wire newNet_1655;
wire n_42293;
wire n_28919;
wire n_5972;
wire n_5636;
wire n_34709;
wire n_1470;
wire n_15988;
wire n_1490;
wire n_38475;
wire delay_sub_ln23_unr25_stage8_stallmux_q_3_;
wire newNet_2118;
wire n_25788;
wire n_25479;
wire n_37546;
wire FE_OCPN1230_n_42201;
wire newNet_3387;
wire n_33216;
wire newNet_154;
wire n_23066;
wire n_36873;
wire n_41997;
wire n_25373;
wire n_23721;
wire n_19019;
wire n_39365;
wire n_4023;
wire n_11888;
wire n_15821;
wire n_32029;
wire n_11191;
wire n_17284;
wire n_25551;
wire n_27461;
wire newNet_3367;
wire FE_OCP_RBN3367_n_44722;
wire n_43111;
wire newNet_1825;
wire newNet_1929;
wire n_35880;
wire n_25199;
wire n_25482;
wire n_35385;
wire n_23850;
wire newNet_2806;
wire FE_RN_1371_0;
wire n_1274;
wire n_36554;
wire n_24432;
wire newNet_1417;
wire n_13755;
wire n_21878;
wire FE_RN_1863_0;
wire n_11226;
wire n_18955;
wire n_6710;
wire n_9674;
wire n_17885;
wire n_19969;
wire newNet_1556;
wire n_20658;
wire n_38254;
wire FE_RN_679_0;
wire n_24093;
wire n_4919;
wire n_39269;
wire FE_OCPN1391_n_7925;
wire newNet_31;
wire n_30061;
wire n_3840;
wire FE_OCPN1468_n_12968;
wire n_10331;
wire n_14343;
wire newNet_1714;
wire n_33482;
wire n_36907;
wire n_37215;
wire n_13651;
wire n_35529;
wire n_26824;
wire newNet_2907;
wire n_41440;
wire n_3670;
wire n_33523;
wire n_39056;
wire n_43292;
wire n_7741;
wire n_14082;
wire n_40537;
wire n_19200;
wire n_35362;
wire beta_29;
wire n_6970;
wire n_30587;
wire newNet_2851;
wire n_27665;
wire newNet_3126;
wire n_8115;
wire FE_OFN761_n_45813;
wire n_2145;
wire n_30629;
wire delay_add_ln22_unr23_stage9_stallmux_q_10_;
wire n_42678;
wire n_36010;
wire n_41361;
wire n_46149;
wire n_5094;
wire n_5871;
wire n_37978;
wire n_36288;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_6_;
wire n_27285;
wire n_19282;
wire n_32536;
wire n_37321;
wire n_13925;
wire FE_OCP_RBN1905_n_29080;
wire n_23772;
wire n_12605;
wire FE_OFN744_n_23604;
wire n_5415;
wire n_7261;
wire FE_RN_951_0;
wire n_30350;
wire n_27366;
wire n_33803;
wire newNet_147;
wire n_3784;
wire n_28278;
wire n_38014;
wire n_21919;
wire n_16262;
wire n_31358;
wire n_34227;
wire n_36307;
wire newNet_1900;
wire n_8144;
wire n_4179;
wire n_14217;
wire n_15726;
wire n_32515;
wire n_36667;
wire n_4947;
wire n_45501;
wire n_38374;
wire FE_OFN755_n_44461;
wire n_41712;
wire n_34925;
wire n_27050;
wire n_24794;
wire n_4796;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_28_;
wire n_18463;
wire newNet_2327;
wire FE_OCPN1491_n_22036;
wire n_45866;
wire n_24032;
wire n_41333;
wire n_37884;
wire n_24982;
wire n_25493;
wire n_6024;
wire FE_RN_201_0;
wire n_9927;
wire FE_OCP_RBN2340_n_29470;
wire n_30971;
wire n_14853;
wire n_24158;
wire n_4720;
wire n_464;
wire n_10500;
wire n_22501;
wire n_28211;
wire n_42956;
wire n_43090;
wire n_19350;
wire n_21834;
wire FE_OCP_RBN2612_n_9075;
wire n_25408;
wire n_3092;
wire n_38705;
wire n_7682;
wire n_41231;
wire n_6884;
wire n_15853;
wire n_33221;
wire n_26801;
wire n_295;
wire newNet_1626;
wire n_40210;
wire n_23437;
wire FE_RN_1465_0;
wire n_416;
wire n_11043;
wire n_6828;
wire n_40128;
wire n_18158;
wire n_36911;
wire n_44954;
wire n_588;
wire n_36233;
wire n_17787;
wire FE_RN_1635_0;
wire n_43657;
wire n_16138;
wire n_17125;
wire n_5664;
wire n_27254;
wire n_17407;
wire n_12528;
wire newNet_3190;
wire newNet_1719;
wire n_43405;
wire n_37570;
wire n_27757;
wire n_3918;
wire n_31534;
wire n_42690;
wire newNet_1451;
wire n_36604;
wire n_38082;
wire n_12526;
wire n_8244;
wire newNet_815;
wire n_34880;
wire n_4286;
wire n_18672;
wire n_703;
wire n_45900;
wire n_39789;
wire n_20154;
wire n_8167;
wire n_15273;
wire n_32793;
wire delay_xor_ln22_unr3_stage2_stallmux_q_17_;
wire n_30217;
wire FE_OCP_RBN2873_n_10477;
wire n_14266;
wire FE_OCP_RBN2846_n_30678;
wire n_14362;
wire n_43073;
wire FE_OCP_RBN3250_delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire n_37391;
wire n_346;
wire FE_OCP_RBN2443_n_42051;
wire n_37271;
wire n_27789;
wire FE_OCP_RBN3475_n_7886;
wire n_8556;
wire n_15259;
wire n_35412;
wire n_26999;
wire n_23739;
wire n_13954;
wire n_28972;
wire n_10882;
wire n_20465;
wire newNet_2768;
wire n_2057;
wire n_8784;
wire n_30210;
wire n_42092;
wire n_35596;
wire n_23837;
wire n_26855;
wire n_29117;
wire n_37289;
wire n_35290;
wire n_39510;
wire n_40346;
wire n_23579;
wire newNet_2114;
wire newNet_2174;
wire newNet_2034;
wire n_32413;
wire n_39095;
wire FE_OCPN996_n_44460;
wire n_16892;
wire n_33380;
wire newNet_193;
wire n_40976;
wire n_30768;
wire n_16889;
wire n_15789;
wire n_37113;
wire n_25074;
wire n_33569;
wire n_4261;
wire n_1842;
wire n_27573;
wire n_28784;
wire n_24959;
wire n_22957;
wire FE_RN_206_0;
wire n_11747;
wire n_19751;
wire n_5982;
wire newNet_3203;
wire n_14089;
wire n_179;
wire n_36745;
wire newNet_3656;
wire n_21295;
wire n_33340;
wire n_14039;
wire FE_RN_1355_0;
wire n_41916;
wire FE_RN_1189_0;
wire n_535;
wire n_34744;
wire n_22499;
wire n_23462;
wire n_6028;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_25_;
wire delay_add_ln22_unr23_stage9_stallmux_q_28_;
wire n_14169;
wire n_19982;
wire n_27035;
wire n_18191;
wire n_15756;
wire n_35535;
wire n_28724;
wire newNet_2269;
wire n_36647;
wire n_4413;
wire delay_add_ln22_unr8_stage4_stallmux_q_26_;
wire newNet_2300;
wire n_3056;
wire n_33456;
wire n_29470;
wire n_36864;
wire newNet_2502;
wire n_42123;
wire n_19904;
wire n_42769;
wire n_8073;
wire n_24137;
wire n_31933;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_17_;
wire FE_OCP_RBN2604_n_39126;
wire n_23776;
wire n_20228;
wire n_20272;
wire FE_RN_377_0;
wire n_33234;
wire n_748;
wire n_2006;
wire n_9853;
wire n_5861;
wire newNet_2278;
wire n_2960;
wire n_4574;
wire n_40194;
wire n_18476;
wire n_20255;
wire n_23221;
wire n_17041;
wire n_42788;
wire n_32170;
wire FE_OCP_RBN2711_n_35075;
wire n_637;
wire n_8185;
wire n_22490;
wire n_5945;
wire n_2890;
wire n_5013;
wire n_19015;
wire newNet_3607;
wire n_25613;
wire n_19027;
wire n_25486;
wire n_36903;
wire n_22900;
wire n_8589;
wire newNet_3683;
wire FE_OCP_RBN1333_n_20249;
wire n_9934;
wire n_43452;
wire n_12054;
wire n_39397;
wire n_27612;
wire n_13280;
wire newNet_3009;
wire n_44038;
wire FE_RN_1346_0;
wire n_23243;
wire newNet_1332;
wire n_11579;
wire n_33698;
wire n_33938;
wire n_32282;
wire n_13960;
wire n_10586;
wire newNet_635;
wire n_32702;
wire FE_RN_81_0;
wire n_40464;
wire n_23341;
wire n_4172;
wire n_17922;
wire n_40597;
wire n_13449;
wire n_30864;
wire FE_RN_1594_0;
wire n_46933;
wire n_16963;
wire n_716;
wire n_46238;
wire n_40224;
wire n_31886;
wire delay_add_ln22_unr8_stage4_stallmux_q_10_;
wire n_16772;
wire n_2808;
wire n_41604;
wire n_31750;
wire n_7723;
wire n_12198;
wire n_13700;
wire FE_OCP_RBN2273_n_2457;
wire n_39004;
wire n_20711;
wire FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_OCP_RBN3440_n_33803;
wire newNet_3516;
wire n_46208;
wire newNet_2386;
wire newNet_3172;
wire n_20419;
wire n_37443;
wire FE_OCP_RBN2992_n_35539;
wire n_5493;
wire newNet_1005;
wire n_37853;
wire n_45181;
wire n_5086;
wire n_7094;
wire n_42173;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_20_;
wire n_23023;
wire n_30289;
wire n_14665;
wire n_19002;
wire n_40771;
wire n_40508;
wire n_37532;
wire FE_RN_1508_0;
wire n_9456;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_25_;
wire n_43226;
wire FE_OCP_RBN2506_n_13896;
wire n_28361;
wire newNet_3194;
wire n_28355;
wire n_34252;
wire n_43327;
wire n_9242;
wire n_23393;
wire n_19801;
wire n_2400;
wire n_34867;
wire n_37692;
wire n_2252;
wire n_19960;
wire n_42141;
wire n_31040;
wire n_19468;
wire n_12111;
wire n_40825;
wire n_20605;
wire n_18721;
wire n_18164;
wire n_10280;
wire n_13157;
wire n_32265;
wire n_41165;
wire n_17155;
wire n_9076;
wire n_13617;
wire n_30558;
wire n_27608;
wire n_982;
wire n_10215;
wire n_21286;
wire n_33163;
wire n_44650;
wire n_30787;
wire n_16060;
wire n_23686;
wire FE_RN_1388_0;
wire n_35747;
wire n_13916;
wire n_15731;
wire n_33512;
wire n_25540;
wire FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__;
wire n_3455;
wire n_9087;
wire n_2380;
wire n_13774;
wire n_36195;
wire n_6344;
wire n_28150;
wire n_30263;
wire n_10848;
wire n_29220;
wire n_14687;
wire n_3054;
wire n_29269;
wire n_13168;
wire n_21084;
wire n_4912;
wire n_29989;
wire n_36279;
wire n_8033;
wire n_31204;
wire n_1345;
wire n_13921;
wire n_2900;
wire n_43735;
wire n_31489;
wire n_29396;
wire n_16880;
wire n_37036;
wire n_43726;
wire n_39504;
wire n_4904;
wire n_4348;
wire n_37750;
wire n_41086;
wire n_27022;
wire n_4754;
wire n_34172;
wire n_13866;
wire n_19440;
wire n_21448;
wire n_4126;
wire n_31990;
wire n_42017;
wire newNet_1489;
wire n_38711;
wire n_25329;
wire n_29482;
wire n_27308;
wire n_24423;
wire n_6645;
wire n_43401;
wire n_9153;
wire n_43608;
wire n_26985;
wire FE_RN_686_0;
wire n_11241;
wire n_1137;
wire n_15584;
wire n_20941;
wire n_37138;
wire newNet_3476;
wire n_32965;
wire n_6365;
wire n_41773;
wire n_43559;
wire n_4760;
wire FE_OCP_RBN3373_n_6745;
wire n_18188;
wire n_39680;
wire n_10326;
wire delay_add_ln22_unr5_stage3_stallmux_q_4_;
wire newNet_2597;
wire n_1026;
wire n_32787;
wire n_15622;
wire n_19514;
wire n_21169;
wire n_41344;
wire n_32569;
wire n_7107;
wire n_13347;
wire newNet_2871;
wire n_34815;
wire n_32466;
wire n_43475;
wire delay_add_ln22_unr14_stage6_stallmux_q_15_;
wire n_10879;
wire n_14564;
wire n_42277;
wire newNet_892;
wire n_540;
wire newNet_2962;
wire n_21844;
wire n_1701;
wire n_40400;
wire n_17507;
wire n_14572;
wire n_38517;
wire n_25292;
wire n_28250;
wire n_2554;
wire n_34546;
wire n_33140;
wire n_17791;
wire n_26961;
wire FE_OCP_RBN3671_FE_RN_470_0;
wire n_14176;
wire n_8788;
wire newNet_871;
wire n_31050;
wire n_762;
wire n_26129;
wire n_21786;
wire n_23920;
wire n_27525;
wire n_8204;
wire n_5098;
wire n_19678;
wire n_10140;
wire n_9135;
wire n_17982;
wire n_23391;
wire n_17677;
wire n_16497;
wire n_7285;
wire n_46244;
wire n_5108;
wire n_21673;
wire n_338;
wire delay_add_ln22_unr17_stage7_stallmux_q_4_;
wire n_13890;
wire n_13050;
wire n_24662;
wire FE_OCP_RBN2150_n_11763;
wire n_5258;
wire FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_10831;
wire n_29789;
wire n_5143;
wire FE_OCP_RBN2544_n_9082;
wire n_28073;
wire n_36828;
wire n_39618;
wire n_37147;
wire newNet_1402;
wire n_5968;
wire n_36093;
wire n_30577;
wire newNet_3713;
wire n_228;
wire n_21612;
wire n_28309;
wire n_4661;
wire newNet_1416;
wire n_18251;
wire n_22312;
wire FE_RN_1800_0;
wire n_40056;
wire n_922;
wire n_14967;
wire n_14747;
wire n_26375;
wire newNet_3731;
wire FE_OCP_RBN2225_n_12729;
wire n_27710;
wire n_41173;
wire n_20899;
wire n_33983;
wire n_34191;
wire n_1625;
wire n_43362;
wire n_8749;
wire n_43776;
wire n_37818;
wire n_6006;
wire newNet_2723;
wire n_37564;
wire n_41054;
wire n_13301;
wire n_38727;
wire n_22201;
wire n_24723;
wire n_6936;
wire n_20976;
wire n_21767;
wire n_31328;
wire n_32696;
wire n_29737;
wire FE_OCP_RBN2761_n_15200;
wire n_21297;
wire n_11978;
wire newNet_1627;
wire n_9602;
wire n_17134;
wire n_5304;
wire n_37590;
wire n_39354;
wire n_39129;
wire FE_RN_1405_0;
wire n_602;
wire n_9861;
wire FE_OCP_RBN2803_n_15706;
wire n_34074;
wire n_36718;
wire n_18799;
wire n_28477;
wire n_38057;
wire n_7311;
wire n_33654;
wire newNet_1734;
wire n_27011;
wire n_32609;
wire n_10446;
wire n_7979;
wire n_40803;
wire n_6131;
wire n_34111;
wire n_32649;
wire n_2573;
wire n_38688;
wire newNet_1915;
wire n_35411;
wire n_30542;
wire n_21994;
wire n_10351;
wire n_37414;
wire n_30829;
wire n_10800;
wire n_7851;
wire n_31285;
wire n_17587;
wire n_9519;
wire n_25529;
wire n_37822;
wire n_22386;
wire FE_OCP_RBN2170_n_32892;
wire n_20432;
wire n_21716;
wire n_27101;
wire newNet_3075;
wire n_32276;
wire n_34914;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_21_;
wire n_26492;
wire n_46178;
wire n_41857;
wire FE_RN_1136_0;
wire n_30595;
wire n_15289;
wire n_14948;
wire n_37048;
wire n_596;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_5_;
wire n_6414;
wire FE_OCPN1532_n_21790;
wire n_1334;
wire n_8015;
wire n_711;
wire n_29035;
wire n_47243;
wire n_20784;
wire n_12384;
wire n_34474;
wire n_38201;
wire n_7322;
wire n_32184;
wire n_21564;
wire n_46423;
wire n_23539;
wire newNet_2208;
wire n_44450;
wire n_401;
wire FE_RN_1251_0;
wire n_41113;
wire n_27301;
wire n_21799;
wire n_20148;
wire n_23251;
wire n_26820;
wire n_12291;
wire FE_OCP_RBN2137_n_11907;
wire n_33059;
wire n_8449;
wire FE_RN_735_0;
wire n_43805;
wire n_40287;
wire newNet_302;
wire n_5703;
wire n_36966;
wire n_39597;
wire n_25466;
wire n_20207;
wire n_41328;
wire n_9838;
wire n_8461;
wire n_23967;
wire n_7027;
wire n_14595;
wire n_8380;
wire FE_RN_960_0;
wire n_29556;
wire n_139;
wire n_24943;
wire n_7759;
wire n_6852;
wire n_10087;
wire FE_OCPN1033_n_28420;
wire n_42829;
wire n_34036;
wire n_12907;
wire n_24712;
wire n_37656;
wire FE_RN_1507_0;
wire newNet_934;
wire n_19451;
wire n_7357;
wire FE_OCP_RBN2798_n_10106;
wire n_24655;
wire n_35175;
wire n_2173;
wire n_38442;
wire n_31584;
wire n_5455;
wire n_42928;
wire n_13947;
wire n_34095;
wire n_41760;
wire FE_OCP_DRV_N1573_n_28869;
wire n_22682;
wire n_39439;
wire n_37511;
wire n_3166;
wire FE_RN_666_0;
wire n_25130;
wire FE_RN_1041_0;
wire n_17918;
wire n_31808;
wire n_34631;
wire n_39235;
wire newNet_4;
wire n_24542;
wire n_31894;
wire n_42522;
wire n_3073;
wire n_33279;
wire newNet_1710;
wire n_14971;
wire n_9188;
wire n_24003;
wire n_12222;
wire n_43711;
wire n_311;
wire FE_OCPN1435_n_19855;
wire n_44711;
wire n_37130;
wire n_42727;
wire n_687;
wire n_36133;
wire n_3125;
wire n_20033;
wire FE_OCP_RBN3515_n_8498;
wire n_32291;
wire n_17431;
wire n_21458;
wire n_5811;
wire n_35486;
wire n_27338;
wire FE_OCP_RBN2794_n_10106;
wire n_12574;
wire n_43526;
wire n_37991;
wire n_1508;
wire n_34594;
wire FE_OCP_RBN3688_n_5130;
wire n_29918;
wire n_35864;
wire n_38787;
wire n_43913;
wire n_24836;
wire n_5586;
wire n_37380;
wire n_20744;
wire newNet_2500;
wire n_43915;
wire newNet_1047;
wire n_23662;
wire FE_RN_763_0;
wire n_38845;
wire n_28971;
wire n_21027;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_1_;
wire n_41398;
wire n_1524;
wire n_33941;
wire n_40147;
wire n_31511;
wire n_41014;
wire n_38531;
wire n_20739;
wire n_24620;
wire FE_RN_776_0;
wire n_1309;
wire n_13610;
wire n_16655;
wire n_41683;
wire n_1979;
wire n_6354;
wire n_33287;
wire n_32863;
wire n_17061;
wire n_42332;
wire FE_OCP_RBN2836_FE_RN_745_0;
wire n_40396;
wire n_7044;
wire n_28666;
wire newNet_2559;
wire n_3529;
wire n_15030;
wire n_16547;
wire n_15700;
wire FE_RN_123_0;
wire n_10952;
wire n_29615;
wire newNet_1680;
wire FE_OCP_RBN3509_n_13860;
wire n_20966;
wire n_11535;
wire n_46974;
wire n_4310;
wire n_25381;
wire FE_OCPN930_n_44083;
wire n_30294;
wire n_38042;
wire newNet_3068;
wire n_8005;
wire n_11495;
wire n_39319;
wire n_5887;
wire newNet_710;
wire n_6109;
wire n_24345;
wire n_8431;
wire n_3018;
wire n_35117;
wire FE_OCP_RBN3451_n_37945;
wire n_29495;
wire n_2476;
wire n_2153;
wire n_13066;
wire n_11350;
wire n_15718;
wire n_9321;
wire n_13229;
wire n_37498;
wire n_10344;
wire n_39134;
wire FE_OCP_RBN2588_n_9492;
wire n_31994;
wire n_27410;
wire n_6163;
wire n_3736;
wire FE_OCP_RBN2690_FE_OCPN843_n_3912;
wire newNet_1784;
wire n_4700;
wire newNet_426;
wire n_2917;
wire n_18141;
wire n_2098;
wire n_2064;
wire n_11797;
wire n_10130;
wire n_41847;
wire FE_OCP_RBN3544_n_44575;
wire n_40612;
wire n_10752;
wire FE_RN_1087_0;
wire n_42138;
wire newNet_120;
wire delay_add_ln22_unr27_stage10_stallmux_q_25_;
wire n_8578;
wire FE_OCP_RBN2738_n_15300;
wire newNet_2679;
wire newNet_24;
wire n_18310;
wire n_38738;
wire n_9286;
wire n_30464;
wire n_40189;
wire n_7739;
wire delay_add_ln22_unr14_stage6_stallmux_q_11_;
wire FE_RN_1728_0;
wire FE_OCPN1051_n_31674;
wire n_31007;
wire newNet_1500;
wire n_44160;
wire n_14918;
wire n_44463;
wire n_18093;
wire newNet_3650;
wire newNet_593;
wire n_23876;
wire n_32298;
wire n_12331;
wire n_18045;
wire newNet_1984;
wire n_45827;
wire n_31387;
wire n_31746;
wire n_27866;
wire n_39676;
wire n_8734;
wire n_24614;
wire n_13292;
wire n_20730;
wire n_44166;
wire n_24380;
wire n_32104;
wire n_37960;
wire FE_RN_1423_0;
wire FE_OCP_RBN1681_n_33491;
wire n_256;
wire n_2963;
wire n_14634;
wire n_26952;
wire n_17845;
wire n_34134;
wire FE_OCP_RBN2911_n_30908;
wire n_24862;
wire n_92;
wire n_7369;
wire n_37501;
wire n_11860;
wire n_36109;
wire n_35847;
wire n_17314;
wire n_33527;
wire n_27291;
wire FE_OCP_RBN1852_n_22556;
wire n_21392;
wire n_2784;
wire n_3592;
wire n_25935;
wire FE_OCPN1409_n_27014;
wire n_18078;
wire newNet_2045;
wire n_12700;
wire n_24629;
wire n_38641;
wire newNet_3086;
wire n_35631;
wire n_37875;
wire n_27876;
wire FE_OCP_RBN3012_n_31117;
wire n_30201;
wire n_30280;
wire n_30871;
wire n_21906;
wire n_40033;
wire FE_RN_367_0;
wire n_5981;
wire n_23168;
wire n_37375;
wire newNet_3467;
wire n_290;
wire n_37183;
wire n_29198;
wire n_27488;
wire n_22397;
wire n_31181;
wire n_4596;
wire FE_RN_1601_0;
wire n_17359;
wire newNet_2950;
wire n_24461;
wire n_36767;
wire n_39637;
wire n_34158;
wire newNet_2202;
wire n_17790;
wire n_6061;
wire FE_RN_1674_0;
wire n_35019;
wire n_38243;
wire n_38816;
wire newNet_645;
wire newNet_2926;
wire n_13906;
wire n_13450;
wire n_8983;
wire n_29157;
wire n_14991;
wire n_8323;
wire newNet_2570;
wire n_19197;
wire n_9983;
wire n_10637;
wire n_434;
wire n_45519;
wire n_26016;
wire delay_xor_ln21_unr3_stage2_stallmux_q_2_;
wire n_32675;
wire beta_25;
wire n_43299;
wire n_35851;
wire n_4433;
wire n_26887;
wire n_15556;
wire n_7246;
wire n_31620;
wire n_40086;
wire n_9664;
wire n_22917;
wire n_27845;
wire n_6486;
wire n_1299;
wire n_847;
wire n_17119;
wire FE_OCPN1483_n_18953;
wire n_2110;
wire n_38894;
wire n_11003;
wire n_37721;
wire FE_RN_999_0;
wire n_28626;
wire n_5036;
wire n_40543;
wire newNet_2820;
wire n_12132;
wire n_45809;
wire n_21920;
wire n_976;
wire n_29801;
wire FE_RN_6_0;
wire newNet_1955;
wire delay_xor_ln22_unr15_stage6_stallmux_q_8_;
wire n_7331;
wire newNet_1258;
wire n_12406;
wire n_12459;
wire n_3373;
wire FE_OCP_RBN3598_FE_OCPN1243_n_44460;
wire FE_RN_1361_0;
wire n_33656;
wire n_5592;
wire n_33025;
wire n_36653;
wire delay_add_ln22_unr17_stage7_stallmux_q_5_;
wire n_30966;
wire n_5693;
wire n_38625;
wire n_14619;
wire n_25924;
wire n_20309;
wire FE_RN_385_0;
wire n_2682;
wire n_37022;
wire n_29811;
wire n_14309;
wire n_44061;
wire FE_RN_1534_0;
wire FE_OCP_RBN2658_n_4101;
wire n_13980;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_26_;
wire newNet_1154;
wire n_25758;
wire n_42992;
wire n_13434;
wire n_34623;
wire n_10885;
wire n_29863;
wire FE_OCP_DRV_N1609_n_20146;
wire n_7087;
wire n_7834;
wire n_19420;
wire n_529;
wire n_9635;
wire n_29385;
wire n_27756;
wire n_5374;
wire n_15247;
wire n_26874;
wire n_35510;
wire n_26524;
wire n_15379;
wire n_44827;
wire n_3190;
wire n_6148;
wire n_6375;
wire n_31472;
wire cos_out_29;
wire n_40561;
wire newNet_1351;
wire n_11029;
wire n_14579;
wire n_18026;
wire newNet_3582;
wire FE_RN_701_0;
wire n_23859;
wire delay_xor_ln22_unr9_stage4_stallmux_q_5_;
wire newNet_768;
wire n_19287;
wire n_14515;
wire FE_RN_1577_0;
wire n_4375;
wire n_26939;
wire n_374;
wire n_29602;
wire FE_RN_813_0;
wire newNet_910;
wire n_29817;
wire n_24764;
wire n_36257;
wire newNet_1722;
wire n_7699;
wire n_7668;
wire n_21279;
wire n_25125;
wire n_26314;
wire n_5164;
wire n_15762;
wire n_32420;
wire n_1433;
wire FE_RN_740_0;
wire n_29574;
wire n_8776;
wire n_19591;
wire n_42026;
wire n_23311;
wire n_26096;
wire n_23414;
wire n_15423;
wire n_36703;
wire n_13033;
wire n_33877;
wire delay_add_ln22_unr20_stage8_stallmux_q_26_;
wire n_23360;
wire n_44027;
wire n_10296;
wire n_23494;
wire n_22880;
wire n_6413;
wire n_13839;
wire newNet_1753;
wire mux_while_ln12_psv_q_5_;
wire n_14779;
wire n_4827;
wire n_36563;
wire newNet_3534;
wire n_40758;
wire n_11600;
wire n_17642;
wire n_34523;
wire n_23718;
wire n_40369;
wire n_45091;
wire n_20319;
wire n_3507;
wire n_30033;
wire n_20167;
wire n_16908;
wire n_2730;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_0_;
wire n_16707;
wire n_21208;
wire n_32110;
wire n_39206;
wire n_15673;
wire n_25647;
wire n_34959;
wire n_168;
wire n_23144;
wire n_40311;
wire FE_RN_1624_0;
wire n_28719;
wire n_20886;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_30_;
wire FE_OCP_RBN1220_n_27835;
wire n_2609;
wire newNet_232;
wire newNet_1772;
wire n_4999;
wire n_23594;
wire n_29364;
wire n_39048;
wire newNet_1840;
wire n_37355;
wire n_1819;
wire n_26194;
wire n_6039;
wire n_14238;
wire n_28124;
wire n_37425;
wire n_22008;
wire n_3722;
wire n_30756;
wire n_28139;
wire n_41928;
wire n_15605;
wire n_27604;
wire FE_OCP_RBN2474_n_8664;
wire n_37923;
wire n_5053;
wire n_35005;
wire n_8523;
wire n_37247;
wire n_6123;
wire n_7891;
wire n_7173;
wire n_9804;
wire n_12751;
wire n_35504;
wire n_3451;
wire n_13726;
wire n_35443;
wire newNet_3457;
wire newNet_520;
wire n_28335;
wire n_41503;
wire n_41419;
wire n_12671;
wire n_29887;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_21_;
wire n_41549;
wire n_20778;
wire newNet_2065;
wire n_7812;
wire n_25821;
wire n_45450;
wire n_31943;
wire n_4068;
wire n_26224;
wire n_35160;
wire FE_OCPN1399_n_8670;
wire n_16456;
wire n_3984;
wire n_31219;
wire n_24828;
wire n_25104;
wire n_12252;
wire n_7574;
wire n_10407;
wire n_21577;
wire n_11086;
wire n_40172;
wire n_41462;
wire n_1188;
wire n_29413;
wire newNet_728;
wire n_26642;
wire n_28225;
wire n_4623;
wire n_14485;
wire n_2646;
wire n_27380;
wire FE_OCP_RBN2984_n_35539;
wire n_28417;
wire FE_OCP_RBN2379_n_3502;
wire newNet_2121;
wire n_30327;
wire delay_xor_ln21_unr3_stage2_stallmux_q_10_;
wire n_4482;
wire n_16835;
wire newNet_1899;
wire newNet_996;
wire n_9578;
wire newNet_472;
wire n_8908;
wire n_11970;
wire n_36530;
wire n_40001;
wire n_28530;
wire n_29127;
wire FE_OCPN1232_n_42201;
wire n_38117;
wire n_17328;
wire n_43552;
wire n_1761;
wire n_47250;
wire n_15008;
wire n_14231;
wire n_25694;
wire n_38362;
wire n_19583;
wire n_26807;
wire n_38562;
wire newNet_88;
wire FE_RN_1387_0;
wire n_4992;
wire n_3334;
wire n_27585;
wire FE_OCP_RBN3053_n_39913;
wire n_34525;
wire n_43413;
wire newNet_1667;
wire n_21773;
wire n_16272;
wire newNet_796;
wire FE_RN_381_0;
wire newNet_2782;
wire n_32900;
wire n_18002;
wire newNet_2865;
wire n_29503;
wire n_20946;
wire n_31979;
wire newNet_2466;
wire n_32664;
wire n_8727;
wire FE_OCP_RBN3582_n_44944;
wire newNet_982;
wire n_32020;
wire FE_RN_874_0;
wire FE_OCP_RBN3429_n_13245;
wire FE_RN_1780_0;
wire n_6334;
wire n_15369;
wire newNet_3113;
wire n_3383;
wire n_11237;
wire FE_OCP_RBN3692_n_10852;
wire n_12208;
wire n_16193;
wire newNet_1264;
wire n_19045;
wire n_34352;
wire n_20048;
wire newNet_1596;
wire n_12688;
wire newNet_2650;
wire newNet_487;
wire newNet_391;
wire n_34558;
wire n_30108;
wire n_33182;
wire n_16737;
wire n_6247;
wire n_16348;
wire n_41785;
wire n_3679;
wire FE_RN_378_0;
wire n_41148;
wire n_43116;
wire n_28903;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_19_;
wire n_605;
wire FE_OCPN1457_n_18426;
wire n_4840;
wire FE_OCP_RBN1915_n_20965;
wire n_7113;
wire newNet_3703;
wire newNet_3019;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_19_;
wire n_26141;
wire n_5187;
wire n_8018;
wire n_30924;
wire n_6739;
wire n_5402;
wire n_25881;
wire newNet_1138;
wire n_26715;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_21_;
wire n_45845;
wire n_40767;
wire n_9058;
wire n_4213;
wire n_7602;
wire n_15542;
wire n_29120;
wire n_2726;
wire n_25175;
wire n_13268;
wire n_12087;
wire n_27214;
wire FE_OCP_RBN3450_n_37945;
wire n_20417;
wire FE_OCP_RBN2590_n_14460;
wire n_1592;
wire n_37475;
wire n_12604;
wire n_4029;
wire n_38556;
wire FE_OCPN1031_n_28448;
wire n_3978;
wire n_23087;
wire n_32821;
wire n_28551;
wire n_35559;
wire newNet_2039;
wire n_11838;
wire n_34381;
wire n_15635;
wire n_40076;
wire n_16277;
wire n_20451;
wire n_31419;
wire n_20187;
wire n_6613;
wire n_10956;
wire n_36866;
wire delay_xor_ln21_unr12_stage5_stallmux_q_3_;
wire n_15396;
wire n_17811;
wire n_24065;
wire n_31089;
wire n_20510;
wire n_14804;
wire n_32541;
wire n_8235;
wire n_37900;
wire n_35754;
wire n_18383;
wire n_18417;
wire n_36852;
wire n_25571;
wire FE_OCP_RBN2863_n_39523;
wire newNet_3130;
wire n_30156;
wire n_27206;
wire n_32995;
wire newNet_2451;
wire newNet_2338;
wire n_17707;
wire n_30575;
wire newNet_1514;
wire n_1242;
wire n_24132;
wire delay_add_ln22_unr5_stage3_stallmux_q_16_;
wire newNet_979;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_18_;
wire n_8047;
wire n_17239;
wire n_10347;
wire n_36404;
wire n_17131;
wire FE_OCP_RBN2611_n_3718;
wire n_19561;
wire n_43677;
wire n_42597;
wire n_13329;
wire n_27242;
wire n_33834;
wire n_24281;
wire n_6711;
wire newNet_3301;
wire newNet_225;
wire n_17632;
wire n_39243;
wire n_37982;
wire n_1261;
wire n_22432;
wire n_6942;
wire newNet_465;
wire n_22686;
wire n_1443;
wire n_27475;
wire n_11123;
wire FE_RN_272_0;
wire n_10530;
wire n_39691;
wire n_35343;
wire newNet_457;
wire newNet_888;
wire FE_OCP_RBN3122_n_32239;
wire n_11517;
wire n_32556;
wire n_153;
wire FE_RN_1827_0;
wire n_2894;
wire n_8678;
wire n_32758;
wire n_11918;
wire newNet_1066;
wire n_5836;
wire n_16393;
wire n_23328;
wire n_35473;
wire newNet_3197;
wire n_10372;
wire n_31443;
wire newNet_3727;
wire n_15265;
wire FE_OCP_RBN2204_n_18242;
wire n_37613;
wire n_13056;
wire n_40583;
wire n_8147;
wire newNet_606;
wire FE_RN_1570_0;
wire n_5276;
wire n_10686;
wire FE_OCP_DRV_N1579_n_35482;
wire n_392;
wire n_36012;
wire n_36365;
wire n_21624;
wire n_43494;
wire newNet_102;
wire FE_OCP_RBN2420_n_24505;
wire n_13408;
wire FE_OCP_RBN2361_n_13818;
wire n_21670;
wire n_21889;
wire n_10610;
wire n_17188;
wire n_6557;
wire n_37219;
wire FE_OCP_RBN3633_n_20568;
wire n_37223;
wire n_28096;
wire n_24327;
wire n_2858;
wire FE_OCP_RBN2929_n_5221;
wire n_2247;
wire n_32001;
wire n_28523;
wire n_3777;
wire FE_OCP_DRV_N1577_n_33904;
wire n_18631;
wire newNet_2887;
wire n_36935;
wire n_43904;
wire n_37285;
wire FE_RN_1421_0;
wire n_9428;
wire n_21801;
wire n_11298;
wire n_21728;
wire FE_OCPN3171_n_34222;
wire FE_OCPN3766_n_14439;
wire n_41167;
wire n_31709;
wire newNet_3392;
wire n_41217;
wire n_4108;
wire n_7593;
wire n_13812;
wire n_11996;
wire FE_OCP_RBN2871_n_39542;
wire n_40846;
wire n_20961;
wire FE_OCP_RBN1211_n_31515;
wire newNet_2640;
wire n_7550;
wire n_32154;
wire n_36328;
wire newNet_306;
wire FE_OCP_RBN3532_n_13765;
wire n_23451;
wire n_31729;
wire n_10906;
wire n_37328;
wire newNet_1396;
wire n_31543;
wire n_8493;
wire n_37350;
wire n_7127;
wire n_27458;
wire n_31636;
wire n_32809;
wire n_21706;
wire n_22413;
wire newNet_64;
wire FE_OCP_RBN3332_n_44962;
wire n_41825;
wire n_39947;
wire n_12800;
wire n_3170;
wire n_15043;
wire n_42902;
wire newNet_2318;
wire n_25716;
wire mux_while_ln12_psv_q_3_;
wire n_10321;
wire delay_sub_ln23_unr21_stage7_stallmux_q_1_;
wire FE_RN_1003_0;
wire n_21360;
wire newNet_865;
wire newNet_2900;
wire newNet_2934;
wire n_24224;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_2_;
wire newNet_332;
wire n_14095;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_14_;
wire n_41090;
wire n_6250;
wire n_17293;
wire n_33269;
wire n_42086;
wire n_33944;
wire FE_OCP_RBN3690_n_16146;
wire newNet_3154;
wire FE_OFN50_n_1045;
wire newNet_2622;
wire n_24218;
wire n_2946;
wire FE_OCP_RBN3693_n_10852;
wire n_37089;
wire FE_OCP_RBN2477_n_8599;
wire newNet_2647;
wire n_6763;
wire n_12559;
wire n_43532;
wire FE_OCP_RBN2499_n_8835;
wire n_14224;
wire n_32148;
wire n_38352;
wire n_35918;
wire n_22789;
wire n_6719;
wire FE_RN_970_0;
wire n_39481;
wire n_997;
wire FE_RN_177_0;
wire newNet_2708;
wire n_36598;
wire FE_RN_1384_0;
wire n_3389;
wire n_23469;
wire newNet_828;
wire FE_RN_810_0;
wire n_16542;
wire n_34023;
wire n_10432;
wire n_12522;
wire n_42444;
wire n_31408;
wire n_6268;
wire n_10287;
wire n_40727;
wire newNet_1689;
wire n_27853;
wire n_2030;
wire n_44713;
wire newNet_862;
wire n_4095;
wire n_26092;
wire n_7205;
wire FE_RN_1167_0;
wire n_33810;
wire n_43901;
wire n_35398;
wire n_46349;
wire n_25894;
wire n_861;
wire n_44722;
wire n_16717;
wire n_36324;
wire n_18419;
wire n_9876;
wire n_9558;
wire n_6500;
wire n_31781;
wire FE_OCPN936_n_42192;
wire FE_OCP_RBN2955_n_26231;
wire n_3959;
wire n_17315;
wire n_28777;
wire n_25389;
wire n_22177;
wire n_44857;
wire n_5666;
wire n_5645;
wire FE_OFN40_n_45813;
wire FE_OCP_RBN3134_n_6567;
wire n_13884;
wire n_43881;
wire n_25000;
wire n_16915;
wire newNet_2296;
wire n_13777;
wire newNet_183;
wire n_12298;
wire n_42008;
wire n_30734;
wire newNet_2403;
wire n_40589;
wire n_22862;
wire FE_RN_1240_0;
wire n_32567;
wire n_37639;
wire n_31153;
wire n_28915;
wire n_6619;
wire n_37668;
wire FE_RN_1467_0;
wire newNet_1855;
wire n_2810;
wire n_10051;
wire n_11586;
wire n_10305;
wire FE_OCP_DRV_N1574_n_28869;
wire newNet_2862;
wire n_18277;
wire n_2980;
wire n_3340;
wire n_9886;
wire n_27550;
wire n_20087;
wire n_958;
wire n_46225;
wire n_14448;
wire n_34983;
wire n_324;
wire n_17737;
wire n_30877;
wire n_800;
wire newNet_1467;
wire n_34132;
wire n_5800;
wire n_13480;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_2_;
wire n_23095;
wire n_17189;
wire n_25624;
wire newNet_2749;
wire n_27437;
wire n_18054;
wire n_18094;
wire FE_OCP_RBN2200_n_13889;
wire n_9594;
wire newNet_1711;
wire n_12762;
wire n_10682;
wire n_42636;
wire newNet_3278;
wire n_15404;
wire FE_RN_765_0;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_12_;
wire n_18165;
wire newNet_3166;
wire n_7553;
wire n_18772;
wire n_8558;
wire n_18638;
wire n_29293;
wire n_27451;
wire n_18523;
wire n_20943;
wire n_2083;
wire n_39981;
wire FE_OCPN978_n_21973;
wire n_40326;
wire n_14484;
wire newNet_335;
wire FE_OCP_RBN2645_n_34980;
wire n_33451;
wire n_2700;
wire n_12213;
wire n_17702;
wire n_33699;
wire n_8101;
wire n_28823;
wire n_8041;
wire n_28214;
wire newNet_3501;
wire n_7017;
wire n_39942;
wire n_2899;
wire n_45060;
wire newNet_2001;
wire n_5671;
wire n_26327;
wire newNet_2645;
wire FE_RN_875_0;
wire n_41871;
wire n_29993;
wire newNet_3402;
wire newNet_2122;
wire newNet_285;
wire n_8786;
wire n_28520;
wire n_3198;
wire delay_add_ln22_unr5_stage3_stallmux_q_0_;
wire n_3799;
wire n_3917;
wire n_8850;
wire n_6286;
wire n_31460;
wire n_18741;
wire n_32825;
wire n_42683;
wire n_27589;
wire n_16270;
wire n_9758;
wire n_38434;
wire n_8482;
wire n_22722;
wire n_33579;
wire n_36632;
wire n_28419;
wire newNet_1004;
wire n_6393;
wire n_44626;
wire n_40325;
wire n_18873;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_27_;
wire n_32725;
wire n_2672;
wire n_33644;
wire n_39376;
wire n_26722;
wire newNet_479;
wire n_17637;
wire n_32658;
wire n_15489;
wire n_13057;
wire n_37178;
wire n_5273;
wire n_39193;
wire n_22801;
wire n_22526;
wire newNet_2888;
wire n_32359;
wire n_33240;
wire n_36411;
wire n_24669;
wire newNet_779;
wire n_24450;
wire newNet_3696;
wire n_32546;
wire n_9898;
wire n_15871;
wire FE_OCP_RBN1167_n_18949;
wire n_34774;
wire n_44256;
wire delay_xor_ln22_unr12_stage5_stallmux_q_12_;
wire newNet_1585;
wire n_23569;
wire FE_OCP_RBN2787_n_15079;
wire n_6071;
wire n_29825;
wire n_24477;
wire n_14823;
wire n_39916;
wire n_38831;
wire n_47257;
wire n_1285;
wire FE_RN_1537_0;
wire n_5818;
wire n_2935;
wire n_22990;
wire n_20906;
wire n_26348;
wire n_33351;
wire n_11008;
wire n_27053;
wire n_21646;
wire newNet_3354;
wire n_38368;
wire FE_OCP_DRV_N1537_n_13646;
wire n_36149;
wire n_13880;
wire n_38541;
wire n_13362;
wire n_3437;
wire n_10757;
wire n_31631;
wire n_9923;
wire n_17048;
wire n_32134;
wire n_37617;
wire n_33264;
wire FE_OCP_RBN1344_n_32520;
wire n_27125;
wire n_27448;
wire n_16561;
wire newNet_3724;
wire n_3396;
wire n_15321;
wire FE_OCP_RBN2780_n_15595;
wire n_2697;
wire n_26917;
wire n_42930;
wire n_20533;
wire n_4432;
wire n_36291;
wire n_10474;
wire n_24706;
wire n_1423;
wire n_3674;
wire n_14139;
wire n_9442;
wire n_7528;
wire n_36901;
wire FE_RN_1344_0;
wire n_8859;
wire delay_add_ln22_unr5_stage3_stallmux_q_26_;
wire n_32835;
wire n_2100;
wire n_34885;
wire n_41345;
wire FE_RN_1277_0;
wire n_19659;
wire n_25056;
wire n_33470;
wire n_16479;
wire n_4083;
wire n_8508;
wire n_22902;
wire n_41273;
wire newNet_240;
wire n_20063;
wire n_43781;
wire n_41092;
wire newNet_2262;
wire newNet_396;
wire n_28416;
wire n_43594;
wire n_42844;
wire newNet_1209;
wire n_18263;
wire n_20241;
wire n_39955;
wire n_9777;
wire n_13948;
wire n_13500;
wire n_28654;
wire n_38922;
wire n_27937;
wire newNet_2018;
wire n_3067;
wire n_16397;
wire n_29414;
wire n_30111;
wire n_31703;
wire newNet_1802;
wire n_11338;
wire n_40717;
wire n_32127;
wire n_36184;
wire n_10513;
wire n_36610;
wire n_41410;
wire newNet_2587;
wire n_37227;
wire n_10872;
wire n_29070;
wire n_23084;
wire n_496;
wire n_7815;
wire n_45843;
wire n_43042;
wire newNet_3112;
wire n_24221;
wire n_17141;
wire n_10093;
wire n_13823;
wire n_40525;
wire newNet_3090;
wire newNet_68;
wire n_42961;
wire n_28110;
wire n_13285;
wire n_32348;
wire FE_OCP_RBN3603_n_8981;
wire n_5286;
wire FE_OCPN1398_n_21973;
wire newNet_1903;
wire newNet_1502;
wire n_18723;
wire n_5511;
wire n_33748;
wire n_15658;
wire FE_OCP_RBN2373_n_8221;
wire FE_OCP_RBN3840_n_19513;
wire n_34250;
wire delay_sub_ln21_unr24_stage9_stallmux_q_5_;
wire n_21929;
wire n_31131;
wire n_7100;
wire n_31896;
wire n_12338;
wire n_27229;
wire n_25360;
wire n_14702;
wire n_27297;
wire newNet_2397;
wire n_37199;
wire n_30757;
wire n_35479;
wire n_25600;
wire n_39902;
wire n_32444;
wire n_8234;
wire n_23500;
wire n_25320;
wire newNet_765;
wire n_7921;
wire n_8138;
wire n_8842;
wire n_28836;
wire n_17018;
wire n_42158;
wire n_46162;
wire n_4762;
wire n_11744;
wire newNet_2658;
wire n_1692;
wire n_43798;
wire FE_RN_631_0;
wire newNet_276;
wire n_19915;
wire n_2323;
wire n_40272;
wire FE_RN_559_0;
wire newNet_805;
wire FE_OCP_RBN1058_n_18267;
wire n_27073;
wire n_43627;
wire n_7592;
wire FE_OCP_RBN3820_n_44061;
wire n_40411;
wire n_12821;
wire n_41546;
wire n_13097;
wire FE_OCP_RBN2684_n_35213;
wire n_43084;
wire n_2390;
wire n_20684;
wire n_32672;
wire n_377;
wire FE_OCP_RBN2519_n_8762;
wire n_39490;
wire n_25061;
wire n_3623;
wire n_4792;
wire n_15803;
wire n_23315;
wire n_14992;
wire n_7789;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_28_;
wire n_3027;
wire delay_add_ln22_unr14_stage6_stallmux_q_0_;
wire n_2864;
wire n_16809;
wire n_25291;
wire FE_OCP_RBN3061_FE_RN_640_0;
wire n_20040;
wire n_35370;
wire n_21838;
wire n_17984;
wire n_7892;
wire newNet_672;
wire n_7579;
wire n_35715;
wire n_26510;
wire n_40739;
wire n_45003;
wire n_34174;
wire n_4411;
wire n_42881;
wire n_31920;
wire n_36944;
wire n_11728;
wire n_23231;
wire n_29797;
wire n_43193;
wire n_5552;
wire n_10363;
wire n_29688;
wire n_34151;
wire n_2640;
wire n_41179;
wire n_19050;
wire n_26463;
wire n_13903;
wire n_1853;
wire n_40863;
wire n_38966;
wire n_14711;
wire n_5858;
wire n_21792;
wire n_37629;
wire n_2556;
wire newNet_3468;
wire newNet_2469;
wire n_11392;
wire n_12739;
wire n_21843;
wire n_6315;
wire n_14462;
wire newNet_1649;
wire n_6732;
wire n_37051;
wire n_18834;
wire FE_OCP_DRV_N3744_FE_OFN737_n_22641;
wire FE_OCP_RBN3379_n_7073;
wire n_27730;
wire n_18622;
wire n_25761;
wire n_31905;
wire newNet_2760;
wire FE_OCP_RBN2807_n_30643;
wire n_33592;
wire n_18513;
wire n_4951;
wire n_37357;
wire newNet_887;
wire newNet_772;
wire n_24421;
wire n_41528;
wire n_10472;
wire n_39097;
wire FE_OCPN3182_FE_OCP_RBN2831_n_10198;
wire n_8413;
wire n_37352;
wire n_12676;
wire n_23821;
wire n_32488;
wire n_30527;
wire n_28609;
wire n_10132;
wire n_14928;
wire n_24178;
wire n_13022;
wire n_6749;
wire n_43561;
wire n_35205;
wire n_38032;
wire n_35171;
wire n_24008;
wire n_20763;
wire FE_OCP_RBN3448_n_37945;
wire n_15372;
wire n_35656;
wire n_9809;
wire n_16607;
wire n_32870;
wire n_11603;
wire n_30409;
wire n_16882;
wire n_36729;
wire n_42540;
wire n_7981;
wire n_10782;
wire n_28995;
wire n_13680;
wire n_17842;
wire n_22615;
wire n_979;
wire FE_OCP_RBN2718_n_9182;
wire FE_OCPN1780_n_24097;
wire newNet_1986;
wire n_563;
wire n_9828;
wire n_7384;
wire n_10972;
wire n_24860;
wire n_41074;
wire newNet_1630;
wire n_22545;
wire n_26206;
wire n_36884;
wire n_14752;
wire n_39300;
wire n_26053;
wire n_3499;
wire n_10142;
wire n_9461;
wire n_31856;
wire FE_RN_1766_0;
wire n_20387;
wire n_10523;
wire n_11010;
wire n_32467;
wire delay_add_ln22_unr14_stage6_stallmux_q_6_;
wire n_38676;
wire n_32853;
wire n_27343;
wire newNet_159;
wire n_11107;
wire n_17057;
wire n_38337;
wire n_40180;
wire n_30245;
wire n_29376;
wire FE_OCP_RBN3842_n_19555;
wire n_24775;
wire n_16050;
wire n_39430;
wire n_34113;
wire n_5054;
wire n_28078;
wire n_9706;
wire n_10174;
wire n_40548;
wire n_29275;
wire n_25579;
wire n_5306;
wire FE_OCP_RBN2337_n_8269;
wire delay_sub_ln22_unr24_stage9_stallmux_q_6_;
wire FE_RN_1523_0;
wire newNet_2151;
wire n_28086;
wire n_8974;
wire delay_xor_ln21_unr3_stage2_stallmux_q_13_;
wire n_4850;
wire FE_RN_698_0;
wire n_1813;
wire FE_RN_1255_0;
wire n_21443;
wire n_28284;
wire n_10881;
wire FE_RN_1233_0;
wire n_12065;
wire n_16931;
wire n_31777;
wire n_42019;
wire n_9101;
wire n_23055;
wire n_42567;
wire n_6761;
wire n_21394;
wire n_28621;
wire n_4894;
wire n_36564;
wire n_37086;
wire n_20480;
wire FE_RN_504_0;
wire n_13545;
wire FE_RN_747_0;
wire n_15519;
wire n_43215;
wire n_24851;
wire n_4236;
wire n_2486;
wire n_28200;
wire n_27717;
wire newNet_3315;
wire newNet_971;
wire n_7830;
wire n_36458;
wire n_37043;
wire n_35832;
wire n_28372;
wire n_25085;
wire n_7948;
wire n_12427;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_25_;
wire n_15125;
wire n_40031;
wire n_31565;
wire n_25595;
wire n_10029;
wire n_14257;
wire n_5103;
wire n_36430;
wire n_39080;
wire n_33908;
wire delay_add_ln22_unr27_stage10_stallmux_q_23_;
wire n_26011;
wire n_33687;
wire n_17599;
wire n_7847;
wire FE_RN_1089_0;
wire n_8325;
wire FE_RN_449_0;
wire n_46989;
wire n_34890;
wire n_24247;
wire n_31579;
wire n_17330;
wire n_37551;
wire n_17749;
wire n_16975;
wire n_28137;
wire n_24674;
wire n_33024;
wire n_3648;
wire n_38829;
wire n_34010;
wire n_33575;
wire FE_RN_526_0;
wire n_39561;
wire FE_RN_1614_0;
wire n_21511;
wire n_33610;
wire FE_RN_1476_0;
wire n_37783;
wire n_32974;
wire n_34625;
wire newNet_3001;
wire newNet_1882;
wire n_4872;
wire n_14508;
wire newNet_58;
wire n_21463;
wire n_18568;
wire n_5681;
wire n_42035;
wire n_11872;
wire n_31975;
wire n_24012;
wire n_33500;
wire n_37451;
wire n_40730;
wire n_18840;
wire n_31766;
wire n_28795;
wire n_21691;
wire n_8173;
wire n_16360;
wire n_5953;
wire n_18756;
wire newNet_3087;
wire n_31225;
wire n_6298;
wire n_6166;
wire n_35445;
wire n_3221;
wire n_3834;
wire n_23774;
wire n_1730;
wire n_46959;
wire n_40751;
wire n_22598;
wire n_27885;
wire n_1983;
wire n_20787;
wire n_24289;
wire n_23791;
wire n_24240;
wire n_17972;
wire FE_OCP_DRV_N1538_n_13646;
wire n_12273;
wire n_38984;
wire delay_xor_ln22_unr18_stage7_stallmux_q_4_;
wire n_8656;
wire n_27012;
wire n_7623;
wire FE_RN_1102_0;
wire n_38751;
wire n_28100;
wire n_2440;
wire n_4353;
wire n_10128;
wire n_15097;
wire n_35133;
wire n_31551;
wire n_28390;
wire n_1658;
wire n_26933;
wire n_1629;
wire n_5284;
wire n_10563;
wire n_41803;
wire n_4671;
wire FE_RN_307_0;
wire FE_RN_1852_0;
wire n_39391;
wire n_16101;
wire n_6642;
wire newNet_2717;
wire n_26580;
wire n_40882;
wire FE_OCP_RBN2157_n_1614;
wire n_6817;
wire delay_xor_ln22_unr3_stage2_stallmux_q_20_;
wire n_12950;
wire n_31646;
wire n_24817;
wire FE_OCPN979_n_21973;
wire n_13743;
wire n_45878;
wire n_8448;
wire FE_OCP_RBN3033_n_43000;
wire n_29710;
wire n_16512;
wire n_29528;
wire n_38284;
wire n_223;
wire n_45488;
wire n_20993;
wire newNet_1186;
wire n_33302;
wire n_4655;
wire n_33311;
wire n_26691;
wire n_43527;
wire n_4974;
wire n_19429;
wire n_17349;
wire n_23970;
wire n_909;
wire n_5266;
wire n_8703;
wire n_36138;
wire n_31382;
wire n_31803;
wire n_43350;
wire n_6019;
wire newNet_722;
wire FE_OCPN1007_n_13962;
wire n_20749;
wire newNet_1920;
wire FE_OCP_RBN3371_n_27970;
wire n_8148;
wire n_28446;
wire delay_xor_ln22_unr3_stage2_stallmux_q_13_;
wire n_7909;
wire newNet_984;
wire newNet_2745;
wire n_42736;
wire newNet_1274;
wire n_43716;
wire n_8739;
wire FE_OCPN1529_n_26090;
wire n_32984;
wire n_23538;
wire n_3165;
wire n_10904;
wire n_17557;
wire FE_RN_179_0;
wire n_32949;
wire n_39244;
wire n_23962;
wire FE_RN_71_0;
wire n_38864;
wire FE_OCP_RBN1147_n_13098;
wire n_32797;
wire n_30506;
wire n_19467;
wire delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_33981;
wire n_41600;
wire newNet_1301;
wire n_13100;
wire n_35348;
wire n_24554;
wire newNet_1686;
wire n_675;
wire n_32086;
wire newNet_423;
wire n_32056;
wire n_28326;
wire n_32928;
wire n_38689;
wire n_23121;
wire n_12110;
wire newNet_2440;
wire n_23991;
wire n_14830;
wire newNet_2214;
wire FE_OCPN1856_n_33341;
wire n_42924;
wire newNet_2607;
wire FE_OCP_RBN1690_n_29491;
wire FE_RN_1612_0;
wire n_3132;
wire n_41089;
wire n_25956;
wire n_2187;
wire n_32235;
wire n_11372;
wire FE_OCP_DRV_N1593_n_34494;
wire FE_RN_892_0;
wire n_36710;
wire n_14212;
wire n_8392;
wire n_6696;
wire n_8008;
wire n_35705;
wire n_8807;
wire n_34458;
wire n_13961;
wire n_14204;
wire n_29603;
wire newNet_3119;
wire n_15019;
wire n_40102;
wire n_23854;
wire n_18539;
wire delay_add_ln22_unr20_stage8_stallmux_q_4_;
wire n_5916;
wire n_1584;
wire FE_RN_1224_0;
wire delay_add_ln22_unr23_stage9_stallmux_q_23_;
wire n_30410;
wire delay_add_ln22_unr11_stage5_stallmux_q_9_;
wire n_35537;
wire n_42177;
wire n_8569;
wire n_24293;
wire n_15951;
wire n_46177;
wire n_43767;
wire n_14877;
wire n_40443;
wire n_27938;
wire n_37576;
wire n_7327;
wire n_39924;
wire n_6931;
wire n_45744;
wire n_20756;
wire n_34166;
wire FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_23_;
wire n_21509;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_22_;
wire n_17582;
wire n_28241;
wire n_32120;
wire n_9306;
wire n_18797;
wire n_38773;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_27_;
wire n_47180;
wire n_35671;
wire n_40241;
wire n_29421;
wire n_46372;
wire FE_OCPN1860_n_35415;
wire n_34964;
wire n_19747;
wire n_3045;
wire FE_RN_1633_0;
wire n_35266;
wire n_8388;
wire delay_add_ln22_unr2_stage2_stallmux_q_26_;
wire n_27086;
wire n_27998;
wire n_29534;
wire n_23783;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_10_;
wire n_10955;
wire n_34814;
wire n_28811;
wire n_38996;
wire n_11692;
wire n_22933;
wire n_37829;
wire n_14584;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_26_;
wire n_12724;
wire n_22243;
wire FE_OCP_RBN1694_n_19052;
wire n_35839;
wire n_28205;
wire n_32931;
wire n_27522;
wire n_26029;
wire n_20702;
wire n_36796;
wire n_21661;
wire n_33141;
wire n_4218;
wire n_37060;
wire n_40159;
wire n_24717;
wire n_34748;
wire n_34197;
wire n_43245;
wire n_7970;
wire FE_OCP_RBN3135_n_6567;
wire n_23254;
wire n_132;
wire n_26945;
wire n_21966;
wire n_14415;
wire n_37855;
wire n_43800;
wire n_22203;
wire n_38906;
wire n_3297;
wire n_36476;
wire n_8663;
wire n_22409;
wire n_19880;
wire n_26767;
wire n_41369;
wire FE_RN_663_0;
wire newNet_1976;
wire n_26563;
wire n_20712;
wire n_26962;
wire newNet_2350;
wire n_10412;
wire n_6137;
wire n_38527;
wire n_17309;
wire n_12088;
wire FE_OCP_RBN2181_n_1916;
wire n_37381;
wire n_18366;
wire n_19827;
wire n_12404;
wire n_42139;
wire n_4227;
wire n_12395;
wire n_7345;
wire n_176;
wire n_25688;
wire n_26283;
wire n_12227;
wire n_20647;
wire n_24330;
wire n_46256;
wire n_14742;
wire n_41059;
wire n_46240;
wire n_39542;
wire n_15159;
wire n_32698;
wire n_27682;
wire n_11927;
wire FE_OCPN1864_n_26171;
wire newNet_389;
wire n_5543;
wire n_8766;
wire FE_OCPN1523_n_45072;
wire FE_RN_1093_0;
wire newNet_1179;
wire n_1179;
wire n_28308;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_4_;
wire n_37141;
wire n_39590;
wire delay_add_ln22_unr17_stage7_stallmux_q_12_;
wire FE_RN_694_0;
wire n_1335;
wire n_37614;
wire n_10124;
wire n_4176;
wire delay_sub_ln22_unr24_stage9_stallmux_q_5_;
wire n_38709;
wire n_32691;
wire n_40074;
wire n_16503;
wire n_31216;
wire n_17402;
wire n_41094;
wire n_38976;
wire n_15079;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_8_;
wire n_27188;
wire n_29104;
wire n_16190;
wire n_9514;
wire n_46285;
wire FE_RN_447_0;
wire n_26133;
wire n_42057;
wire n_3738;
wire n_25354;
wire n_24941;
wire n_3069;
wire n_39755;
wire n_31594;
wire n_19458;
wire FE_RN_1825_0;
wire n_31530;
wire n_32687;
wire n_29854;
wire n_25906;
wire n_1555;
wire n_7832;
wire n_45472;
wire n_39706;
wire n_36047;
wire n_21233;
wire n_34438;
wire n_37719;
wire n_16300;
wire n_23143;
wire n_15730;
wire n_2251;
wire n_20603;
wire n_37797;
wire n_35219;
wire n_35499;
wire FE_OCP_RBN3637_n_44490;
wire n_29848;
wire n_41471;
wire newNet_1771;
wire n_30543;
wire newNet_80;
wire n_42708;
wire n_12733;
wire n_782;
wire n_12646;
wire n_19975;
wire n_10366;
wire n_26156;
wire n_13150;
wire newNet_1364;
wire FE_OCP_RBN3708_n_31396;
wire newNet_3580;
wire n_3254;
wire delay_xor_ln21_unr21_stage8_stallmux_q_10_;
wire n_9235;
wire n_23020;
wire n_42251;
wire n_40009;
wire n_12190;
wire n_15943;
wire n_37139;
wire n_37462;
wire n_15629;
wire n_11581;
wire n_34999;
wire n_34445;
wire n_32384;
wire n_40359;
wire n_3821;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_29_;
wire n_21291;
wire FE_RN_608_0;
wire n_41941;
wire n_33356;
wire n_13799;
wire n_2306;
wire n_4209;
wire n_9356;
wire n_31212;
wire n_7993;
wire newNet_2066;
wire n_19785;
wire n_40645;
wire n_32453;
wire n_6325;
wire n_39137;
wire n_31024;
wire n_34615;
wire n_27659;
wire n_23750;
wire n_34401;
wire FE_OCP_RBN2971_n_31239;
wire n_11279;
wire FE_RN_321_0;
wire n_39099;
wire n_34494;
wire FE_OCPN1515_n_35367;
wire n_18220;
wire n_41427;
wire n_36096;
wire n_40897;
wire n_43601;
wire n_35379;
wire n_33328;
wire n_989;
wire n_35148;
wire n_16204;
wire n_23175;
wire newNet_1000;
wire n_19640;
wire n_30821;
wire n_29720;
wire n_31306;
wire n_15237;
wire FE_OCP_RBN3501_n_8187;
wire FE_OCP_RBN2133_n_45508;
wire n_10259;
wire n_2263;
wire n_17157;
wire newNet_2674;
wire n_3418;
wire newNet_1806;
wire n_7247;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_22_;
wire n_41264;
wire n_28155;
wire n_17766;
wire n_42852;
wire delay_add_ln22_unr5_stage3_stallmux_q_8_;
wire n_14744;
wire n_35122;
wire n_30859;
wire FE_OCP_RBN3396_n_28651;
wire n_3127;
wire n_28117;
wire n_28333;
wire n_41386;
wire n_7677;
wire n_2990;
wire n_36272;
wire FE_OCPN1451_n_27518;
wire n_28568;
wire n_41665;
wire n_31397;
wire n_25138;
wire n_20918;
wire n_19815;
wire n_7715;
wire n_36517;
wire n_4274;
wire FE_OCP_RBN3843_n_24972;
wire n_5799;
wire n_291;
wire n_39538;
wire n_11183;
wire n_33136;
wire FE_OCPN843_n_3912;
wire n_36245;
wire n_16557;
wire n_10263;
wire newNet_3473;
wire n_43206;
wire n_35877;
wire n_8180;
wire n_36728;
wire n_22812;
wire n_5490;
wire n_21629;
wire n_3566;
wire n_2407;
wire newNet_2613;
wire n_16215;
wire n_1075;
wire n_39835;
wire n_32707;
wire delay_xor_ln21_unr12_stage5_stallmux_q_10_;
wire n_19948;
wire n_3326;
wire n_18817;
wire n_399;
wire n_13307;
wire n_806;
wire n_4907;
wire n_46421;
wire n_28676;
wire n_1892;
wire newNet_3209;
wire n_21285;
wire n_10692;
wire n_15808;
wire n_7786;
wire n_1742;
wire n_22972;
wire n_32982;
wire newNet_2505;
wire n_16011;
wire n_10816;
wire n_40989;
wire n_14949;
wire n_41751;
wire n_41918;
wire n_39223;
wire FE_RN_1672_0;
wire n_1571;
wire n_11557;
wire n_42656;
wire n_3856;
wire newNet_640;
wire n_6777;
wire FE_OCP_RBN3037_n_47269;
wire n_26469;
wire newNet_2701;
wire FE_RN_1360_0;
wire n_9724;
wire n_456;
wire FE_RN_518_0;
wire n_1348;
wire n_6415;
wire FE_OCP_RBN2110_n_6616;
wire n_15698;
wire n_39176;
wire n_4535;
wire FE_RN_1533_0;
wire n_44031;
wire n_27099;
wire n_33458;
wire n_32856;
wire n_9334;
wire n_7429;
wire n_19622;
wire n_20209;
wire n_34820;
wire newNet_3667;
wire n_21062;
wire FE_OCPN1425_n_18099;
wire n_23357;
wire n_38049;
wire newNet_2108;
wire n_12199;
wire n_40498;
wire n_19988;
wire n_2219;
wire n_20948;
wire n_6230;
wire n_11280;
wire n_32472;
wire n_41390;
wire n_32906;
wire n_26379;
wire n_25723;
wire n_38181;
wire n_31916;
wire n_32766;
wire n_32101;
wire delay_xor_ln22_unr18_stage7_stallmux_q_6_;
wire n_36588;
wire delay_add_ln22_unr14_stage6_stallmux_q_1_;
wire newNet_2385;
wire n_15295;
wire n_18009;
wire n_25874;
wire FE_RN_352_0;
wire n_37654;
wire n_5375;
wire n_35988;
wire FE_RN_343_0;
wire n_34569;
wire n_35633;
wire newNet_1873;
wire n_23930;
wire n_2704;
wire n_29193;
wire n_16811;
wire n_13116;
wire n_39063;
wire n_29395;
wire n_22950;
wire n_19488;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_12_;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_27_;
wire delay_add_ln22_unr5_stage3_stallmux_q_10_;
wire n_46935;
wire n_35090;
wire n_17988;
wire n_2802;
wire FE_RN_1456_0;
wire n_23326;
wire n_25839;
wire n_32505;
wire n_38554;
wire n_5779;
wire n_14407;
wire n_39380;
wire n_8562;
wire n_32285;
wire n_24419;
wire n_16742;
wire n_654;
wire n_31829;
wire n_27792;
wire n_41073;
wire n_26687;
wire FE_RN_1544_0;
wire n_38428;
wire n_30488;
wire n_20330;
wire n_40060;
wire n_3696;
wire n_28173;
wire FE_OCP_DRV_N1583_n_30917;
wire newNet_3620;
wire n_23396;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_16_;
wire n_30707;
wire FE_OCP_RBN3125_n_27578;
wire newNet_1225;
wire FE_OFN811_n_29140;
wire n_40377;
wire n_36742;
wire n_16961;
wire n_14004;
wire n_14662;
wire newNet_1059;
wire n_38667;
wire n_15811;
wire n_46387;
wire n_33774;
wire n_24834;
wire n_3405;
wire delay_xor_ln21_unr6_stage3_stallmux_q_2_;
wire n_36761;
wire newNet_2036;
wire n_31482;
wire n_28727;
wire n_16372;
wire n_33433;
wire n_4571;
wire n_23600;
wire n_3145;
wire FE_OCP_RBN3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_22183;
wire newNet_1730;
wire delay_add_ln22_unr23_stage9_stallmux_q_5_;
wire n_42206;
wire n_20819;
wire n_22434;
wire n_42099;
wire delay_add_ln22_unr8_stage4_stallmux_q_1_;
wire newNet_1670;
wire n_17442;
wire n_20277;
wire n_39165;
wire n_13952;
wire n_22382;
wire n_43854;
wire n_3020;
wire n_22823;
wire n_28575;
wire n_27960;
wire newNet_930;
wire n_36015;
wire n_16801;
wire n_232;
wire n_20157;
wire n_7204;
wire n_12204;
wire n_694;
wire n_1602;
wire delay_xor_ln21_unr6_stage3_stallmux_q_12_;
wire n_24905;
wire n_26764;
wire n_21761;
wire newNet_2659;
wire n_10988;
wire n_34317;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_24_;
wire n_815;
wire n_3684;
wire n_5561;
wire delay_add_ln22_unr5_stage3_stallmux_q_13_;
wire n_32356;
wire n_18996;
wire FE_RN_1212_0;
wire n_11477;
wire FE_OCP_RBN1717_n_20734;
wire n_30616;
wire n_35454;
wire FE_OCPN1429_n_23792;
wire n_17102;
wire newNet_1653;
wire n_25907;
wire n_1578;
wire n_26531;
wire n_23291;
wire n_38063;
wire n_7378;
wire n_9507;
wire newNet_2155;
wire n_18210;
wire n_11151;
wire n_42515;
wire n_17100;
wire newNet_2254;
wire n_1921;
wire n_4841;
wire n_1771;
wire n_5078;
wire n_18460;
wire n_426;
wire n_28271;
wire n_19295;
wire n_23649;
wire n_8540;
wire n_41101;
wire n_40138;
wire newNet_2767;
wire delay_add_ln22_unr11_stage5_stallmux_q_31_;
wire n_14899;
wire n_41475;
wire n_32919;
wire n_6973;
wire n_1173;
wire n_32138;
wire n_43005;
wire n_34512;
wire n_16133;
wire n_19241;
wire n_22890;
wire n_12602;
wire n_45507;
wire n_29381;
wire n_2843;
wire n_33801;
wire n_24156;
wire n_29000;
wire FE_OCP_RBN2799_n_15434;
wire n_38781;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_0_;
wire n_8697;
wire n_37844;
wire n_7073;
wire n_39488;
wire newNet_1848;
wire n_9532;
wire n_43890;
wire FE_RN_1179_0;
wire n_34441;
wire FE_RN_590_0;
wire n_18705;
wire n_12083;
wire n_37067;
wire FE_RN_1254_0;
wire n_35796;
wire FE_RN_1433_0;
wire newNet_3699;
wire n_5640;
wire FE_OCP_RBN2670_n_20249;
wire n_33132;
wire n_28907;
wire n_15285;
wire n_2314;
wire n_35318;
wire n_9035;
wire n_26881;
wire n_126;
wire n_32719;
wire n_8464;
wire n_22703;
wire n_35799;
wire n_30407;
wire n_12139;
wire n_34537;
wire n_20159;
wire n_26948;
wire n_15981;
wire n_3601;
wire newNet_47;
wire n_42187;
wire delay_add_ln22_unr14_stage6_stallmux_q_14_;
wire n_14382;
wire FE_RN_473_0;
wire n_33247;
wire newNet_3310;
wire n_38392;
wire n_3653;
wire n_11710;
wire FE_RN_1769_0;
wire n_28832;
wire n_15893;
wire FE_OCP_RBN2983_n_26767;
wire n_18765;
wire n_32684;
wire n_21857;
wire newNet_2876;
wire n_30624;
wire n_34239;
wire n_30650;
wire FE_OCP_RBN3473_n_7886;
wire n_30024;
wire n_4602;
wire n_17659;
wire n_36068;
wire newNet_3022;
wire n_6331;
wire n_14087;
wire newNet_2635;
wire n_9584;
wire n_2814;
wire n_32089;
wire n_4264;
wire n_11026;
wire FE_OCP_RBN3529_n_13765;
wire n_5015;
wire n_19770;
wire n_31462;
wire n_35868;
wire n_41715;
wire n_40707;
wire n_8207;
wire n_29311;
wire newNet_2965;
wire n_21733;
wire n_4925;
wire n_43051;
wire n_32295;
wire n_10106;
wire n_28882;
wire FE_OCP_RBN3459_n_7886;
wire n_29589;
wire n_11192;
wire n_31454;
wire n_6564;
wire n_25397;
wire n_22535;
wire n_37270;
wire n_23000;
wire n_30723;
wire n_41452;
wire n_37002;
wire n_24235;
wire n_23518;
wire n_27824;
wire n_812;
wire n_25134;
wire n_35332;
wire n_38272;
wire FE_OCP_RBN2745_n_47011;
wire n_15233;
wire n_34807;
wire n_3259;
wire n_31437;
wire n_27643;
wire n_7337;
wire n_29691;
wire n_41994;
wire n_10286;
wire n_19900;
wire n_8597;
wire FE_RN_938_0;
wire n_38916;
wire n_6277;
wire FE_OCP_RBN2879_n_15553;
wire n_19180;
wire n_22521;
wire n_7586;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_1_;
wire n_37768;
wire n_15723;
wire n_6245;
wire n_20051;
wire n_33962;
wire n_22736;
wire n_5198;
wire n_5309;
wire n_560;
wire FE_OCP_RBN2681_n_15048;
wire n_4484;
wire FE_RN_1121_0;
wire n_24898;
wire n_12532;
wire FE_OCP_RBN2229_n_7598;
wire n_6439;
wire n_39800;
wire n_29265;
wire n_8057;
wire newNet_75;
wire newNet_3128;
wire newNet_1717;
wire n_24251;
wire n_16170;
wire n_35346;
wire n_46365;
wire n_40215;
wire n_38550;
wire n_30298;
wire n_14021;
wire n_42218;
wire n_33437;
wire n_2968;
wire n_42151;
wire n_23183;
wire n_38259;
wire FE_RN_1047_0;
wire n_32228;
wire n_27814;
wire n_15477;
wire n_1273;
wire n_17568;
wire n_5139;
wire n_14228;
wire FE_OCP_DRV_N1601_n_21639;
wire newNet_3347;
wire n_4626;
wire n_36435;
wire n_39446;
wire n_11738;
wire n_35901;
wire n_36875;
wire n_24573;
wire FE_OCP_DRV_N1599_n_21493;
wire n_2289;
wire n_18268;
wire n_35699;
wire n_38333;
wire n_31152;
wire n_24684;
wire n_44847;
wire n_26695;
wire FE_OCP_RBN2217_FE_OCPN950_n_28595;
wire n_3549;
wire n_15865;
wire n_23151;
wire n_2949;
wire n_21110;
wire FE_RN_734_0;
wire n_14400;
wire n_47269;
wire n_24200;
wire newNet_1437;
wire n_46340;
wire n_13972;
wire n_24228;
wire n_24505;
wire n_39123;
wire n_23951;
wire n_286;
wire FE_OCP_RBN3849_n_20290;
wire n_10506;
wire n_29970;
wire n_36302;
wire FE_RN_1617_0;
wire n_41431;
wire n_33378;
wire n_2927;
wire n_35897;
wire n_38303;
wire n_7276;
wire n_47239;
wire newNet_854;
wire newNet_128;
wire n_43521;
wire n_25582;
wire n_4356;
wire n_15065;
wire n_8089;
wire FE_RN_1151_0;
wire n_41813;
wire newNet_2229;
wire n_37951;
wire n_14981;
wire n_38011;
wire n_12013;
wire n_23558;
wire n_44259;
wire newNet_295;
wire n_4965;
wire n_20000;
wire FE_OCPN957_n_39096;
wire n_4424;
wire n_21426;
wire n_37740;
wire n_31508;
wire n_4285;
wire n_36362;
wire n_17446;
wire n_32055;
wire n_6715;
wire n_28965;
wire n_24092;
wire newNet_1824;
wire FE_OCP_DRV_N1589_n_21343;
wire FE_RN_1511_0;
wire n_33013;
wire n_18995;
wire n_25986;
wire n_28789;
wire n_10315;
wire newNet_2141;
wire newNet_3099;
wire n_13375;
wire n_29426;
wire n_42536;
wire n_27556;
wire n_2228;
wire newNet_2525;
wire n_1049;
wire FE_OCP_RBN2523_n_8951;
wire n_33487;
wire n_38144;
wire n_11112;
wire n_39973;
wire FE_RN_1264_0;
wire n_5316;
wire n_10689;
wire n_41864;
wire newNet_468;
wire n_42888;
wire n_17801;
wire n_19368;
wire n_26906;
wire n_25476;
wire n_11895;
wire n_17387;
wire n_32553;
wire FE_OCPN1415_FE_OCP_RBN1362_n_20504;
wire n_26146;
wire n_36334;
wire n_28996;
wire n_19736;
wire n_30910;
wire n_19835;
wire newNet_3660;
wire n_2799;
wire FE_RN_651_0;
wire n_1216;
wire n_39777;
wire n_20657;
wire n_25650;
wire newNet_840;
wire newNet_2578;
wire newNet_3462;
wire n_29706;
wire n_23029;
wire n_5371;
wire n_14444;
wire n_613;
wire n_22087;
wire n_30253;
wire n_42752;
wire n_38478;
wire sin_out_30;
wire n_8667;
wire FE_OCP_RBN2231_n_13141;
wire n_29189;
wire n_19437;
wire n_40972;
wire FE_OCP_RBN2897_n_45484;
wire n_40256;
wire n_34382;
wire FE_OCP_RBN1346_n_19270;
wire n_30338;
wire n_36999;
wire n_27039;
wire n_8927;
wire n_37302;
wire newNet_454;
wire n_2201;
wire FE_OCP_RBN3334_n_44962;
wire FE_OCP_RBN2941_FE_RN_473_0;
wire n_2973;
wire n_22755;
wire newNet_1142;
wire newNet_813;
wire n_6049;
wire n_36770;
wire n_12261;
wire newNet_3647;
wire FE_OCPN1502_n_20723;
wire n_16231;
wire n_44920;
wire n_18847;
wire FE_OCP_RBN3104_n_40561;
wire n_40081;
wire n_29927;
wire n_17083;
wire n_42149;
wire n_33671;
wire FE_OCP_RBN3065_n_22170;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_6_;
wire n_29330;
wire n_88;
wire FE_OCP_RBN3700_n_43015;
wire n_10567;
wire n_28263;
wire n_36422;
wire n_19730;
wire FE_RN_270_0;
wire n_2130;
wire n_4948;
wire n_28435;
wire n_41304;
wire FE_RN_845_0;
wire n_25239;
wire n_30681;
wire n_25914;
wire newNet_1924;
wire n_3245;
wire FE_RN_124_0;
wire n_11454;
wire n_37670;
wire newNet_1118;
wire n_2274;
wire n_27170;
wire n_12315;
wire n_3385;
wire n_34858;
wire n_23771;
wire n_10383;
wire n_5939;
wire n_28770;
wire n_5218;
wire n_34941;
wire n_5175;
wire n_21143;
wire n_25111;
wire n_28423;
wire n_30443;
wire beta_17;
wire n_33276;
wire n_21127;
wire n_18146;
wire n_12322;
wire n_3003;
wire FE_OCP_RBN3723_n_16975;
wire newNet_90;
wire n_2479;
wire newNet_1253;
wire n_8403;
wire n_42935;
wire n_33741;
wire n_28043;
wire n_27044;
wire newNet_1132;
wire n_43832;
wire n_36838;
wire n_33556;
wire newNet_1697;
wire n_21177;
wire n_23092;
wire n_10900;
wire n_40418;
wire FE_OCP_RBN2885_n_35517;
wire n_30374;
wire n_4528;
wire FE_OCP_RBN1850_n_22639;
wire n_2266;
wire n_12217;
wire delay_add_ln22_unr11_stage5_stallmux_q_14_;
wire n_23330;
wire n_17004;
wire FE_OFN735_n_22641;
wire n_17578;
wire n_3848;
wire n_4331;
wire n_46982;
wire n_4054;
wire n_35088;
wire newNet_1571;
wire n_11632;
wire n_19534;
wire n_16762;
wire n_22695;
wire n_18933;
wire n_43742;
wire n_9949;
wire n_28209;
wire n_40477;
wire n_5029;
wire n_19855;
wire n_42318;
wire n_962;
wire n_18117;
wire n_18444;
wire n_15867;
wire n_26318;
wire n_15965;
wire n_1060;
wire n_11200;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_17_;
wire FE_RN_1325_0;
wire n_38381;
wire newNet_3169;
wire n_30001;
wire n_17190;
wire n_17123;
wire n_36375;
wire n_12713;
wire n_46963;
wire n_24398;
wire FE_RN_887_0;
wire n_13142;
wire n_11256;
wire n_4315;
wire n_41447;
wire n_12850;
wire n_17231;
wire FE_RN_1016_0;
wire n_32498;
wire n_39655;
wire n_43545;
wire n_41186;
wire n_14639;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_18_;
wire n_671;
wire n_28911;
wire n_31814;
wire FE_OCPN1731_n_34369;
wire n_14819;
wire n_40454;
wire n_37620;
wire n_31611;
wire n_25306;
wire n_43467;
wire n_35623;
wire n_13632;
wire n_9262;
wire n_4916;
wire n_22921;
wire n_40155;
wire n_8197;
wire n_16408;
wire n_12447;
wire n_6034;
wire n_2052;
wire n_39307;
wire n_21696;
wire n_27766;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_24_;
wire n_15270;
wire n_15170;
wire FE_OCP_DRV_N3745_FE_OFN737_n_22641;
wire n_33197;
wire sin_out_5;
wire n_42023;
wire delay_add_ln22_unr8_stage4_stallmux_q_4_;
wire n_42225;
wire n_5380;
wire n_37154;
wire n_34452;
wire FE_OCP_RBN2924_n_5130;
wire n_42261;
wire FE_RN_1757_0;
wire n_28053;
wire n_36000;
wire n_23132;
wire n_1006;
wire n_1486;
wire newNet_3700;
wire n_35641;
wire n_41658;
wire n_2769;
wire n_9900;
wire n_14328;
wire newNet_1746;
wire n_35785;
wire n_8420;
wire n_12125;
wire n_35195;
wire n_34108;
wire n_1151;
wire n_16426;
wire n_7361;
wire n_1580;
wire n_28142;
wire n_13391;
wire n_11909;
wire n_27623;
wire n_1866;
wire FE_OCPN3756_n_13889;
wire n_12482;
wire n_26785;
wire n_13245;
wire n_1256;
wire n_33167;
wire n_7765;
wire n_36990;
wire n_37610;
wire n_14276;
wire n_4441;
wire n_4465;
wire n_28130;
wire n_31120;
wire n_4801;
wire n_20728;
wire newNet_173;
wire n_20568;
wire n_302;
wire n_18584;
wire n_10941;
wire FE_RN_809_0;
wire n_31312;
wire n_18448;
wire FE_OCP_RBN2317_n_41420;
wire cos_out_21;
wire n_14124;
wire newNet_2786;
wire newNet_3411;
wire n_1297;
wire n_42001;
wire n_17915;
wire n_20105;
wire n_18218;
wire n_39716;
wire n_26808;
wire newNet_1336;
wire n_23216;
wire FE_RN_1774_0;
wire n_40577;
wire n_14558;
wire n_40776;
wire n_2073;
wire n_36992;
wire FE_OCP_RBN2454_n_14157;
wire n_16681;
wire newNet_1113;
wire n_15427;
wire n_41292;
wire n_34405;
wire n_10603;
wire n_40604;
wire n_19950;
wire newNet_3442;
wire n_10402;
wire n_34043;
wire n_12329;
wire n_28330;
wire n_14903;
wire n_42316;
wire n_27256;
wire n_17417;
wire n_1699;
wire n_7888;
wire n_23679;
wire n_28187;
wire n_2748;
wire n_33441;
wire n_41678;
wire n_4556;
wire n_11823;
wire n_10356;
wire n_4202;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_8_;
wire n_10293;
wire n_1368;
wire n_8684;
wire n_15433;
wire n_42360;
wire n_1397;
wire n_37709;
wire n_28091;
wire n_46;
wire n_31280;
wire n_26797;
wire n_40152;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_8_;
wire newNet_1069;
wire n_15924;
wire n_5393;
wire n_3353;
wire newNet_3325;
wire n_19326;
wire FE_RN_1394_0;
wire n_19317;
wire n_43760;
wire n_39734;
wire newNet_1181;
wire delay_xor_ln21_unr3_stage2_stallmux_q_20_;
wire newNet_2683;
wire n_32940;
wire newNet_247;
wire n_21859;
wire FE_OFN825_n_5067;
wire n_40808;
wire n_17146;
wire newNet_3736;
wire n_6745;
wire newNet_2916;
wire n_2327;
wire newNet_1712;
wire n_13388;
wire n_22960;
wire n_18237;
wire n_19706;
wire n_17742;
wire n_13644;
wire n_4365;
wire n_41198;
wire n_24990;
wire n_28473;
wire n_32598;
wire n_7282;
wire n_42053;
wire n_5431;
wire n_25245;
wire n_28950;
wire n_43235;
wire n_2447;
wire FE_OCP_RBN2784_n_9859;
wire n_21719;
wire newNet_3290;
wire FE_RN_491_0;
wire n_20699;
wire n_1540;
wire n_22870;
wire n_17437;
wire n_43134;
wire n_32511;
wire n_27944;
wire n_10193;
wire n_31042;
wire newNet_502;
wire n_42965;
wire n_2176;
wire n_8396;
wire newNet_2477;
wire n_1021;
wire n_32869;
wire n_17171;
wire n_3632;
wire n_25032;
wire n_14286;
wire n_15575;
wire n_6950;
wire n_40833;
wire n_35239;
wire n_42831;
wire newNet_3224;
wire n_40264;
wire n_9200;
wire delay_xor_ln22_unr3_stage2_stallmux_q_21_;
wire n_12295;
wire n_19178;
wire n_10624;
wire n_42638;
wire n_33919;
wire n_4587;
wire n_7968;
wire FE_RN_1265_0;
wire n_29905;
wire n_18185;
wire n_10748;
wire n_11396;
wire n_40515;
wire n_26427;
wire n_11169;
wire delay_xor_ln21_unr3_stage2_stallmux_q_14_;
wire newNet_1510;
wire n_11848;
wire n_16982;
wire n_42170;
wire n_27725;
wire n_8900;
wire n_28351;
wire n_13764;
wire n_24792;
wire n_10319;
wire n_19829;
wire n_37609;
wire n_21072;
wire n_5692;
wire n_31862;
wire n_14872;
wire n_5249;
wire n_20903;
wire n_43075;
wire n_22667;
wire FE_OCP_RBN2353_n_13858;
wire delay_add_ln22_unr27_stage10_stallmux_q_19_;
wire n_39494;
wire n_21191;
wire n_17304;
wire n_25358;
wire n_35825;
wire n_3119;
wire n_8619;
wire n_40639;
wire n_24192;
wire n_18608;
wire n_1951;
wire n_7036;
wire n_38036;
wire n_14855;
wire n_5702;
wire n_26844;
wire n_38438;
wire n_19663;
wire n_35210;
wire n_14114;
wire n_6675;
wire newNet_1052;
wire n_5741;
wire n_30948;
wire n_24485;
wire n_2458;
wire delay_xor_ln21_unr9_stage4_stallmux_q_12_;
wire n_273;
wire n_10499;
wire n_12414;
wire n_34377;
wire FE_RN_1680_0;
wire n_14186;
wire n_16197;
wire n_8546;
wire n_14393;
wire n_10033;
wire delay_add_ln22_unr23_stage9_stallmux_q_3_;
wire FE_OCPN1734_n_16143;
wire n_21312;
wire n_1653;
wire n_10935;
wire cos_out_12;
wire FE_RN_297_0;
wire n_6887;
wire n_4722;
wire n_6923;
wire FE_OCP_RBN3728_FE_RN_1787_0;
wire n_25410;
wire n_8632;
wire n_1494;
wire n_33640;
wire n_8642;
wire n_16312;
wire n_39084;
wire newNet_1029;
wire FE_OCPN971_n_14716;
wire n_26542;
wire n_14775;
wire n_15791;
wire n_15546;
wire n_37106;
wire n_24434;
wire n_35576;
wire n_13924;
wire newNet_39;
wire n_15216;
wire n_33794;
wire newNet_1624;
wire n_9173;
wire n_1616;
wire FE_RN_287_0;
wire n_34687;
wire n_3773;
wire FE_OCPN1747_n_23354;
wire n_1289;
wire delay_xor_ln22_unr9_stage4_stallmux_q_9_;
wire n_20717;
wire newNet_3405;
wire n_35128;
wire FE_OCP_RBN2462_n_3076;
wire n_28991;
wire FE_OCP_RBN1200_n_25763;
wire n_31878;
wire n_27272;
wire n_11410;
wire n_43907;
wire n_17822;
wire n_10146;
wire n_3131;
wire FE_RN_1239_0;
wire n_13427;
wire newNet_2293;
wire newNet_2563;
wire n_41976;
wire n_40045;
wire n_20120;
wire n_778;
wire n_2776;
wire n_34844;
wire FE_RN_1022_0;
wire newNet_1781;
wire n_41836;
wire n_23981;
wire n_22511;
wire newNet_1412;
wire n_8628;
wire n_34804;
wire n_39471;
wire n_18427;
wire n_21099;
wire n_37995;
wire n_1196;
wire newNet_1032;
wire n_29717;
wire n_42343;
wire n_182;
wire n_5607;
wire n_26000;
wire n_17282;
wire n_610;
wire n_16357;
wire n_225;
wire sin_out_21;
wire delay_add_ln22_unr2_stage2_stallmux_q_30_;
wire n_47011;
wire FE_RN_1366_0;
wire n_24343;
wire n_22336;
wire n_22016;
wire n_42660;
wire n_44862;
wire FE_OCP_DRV_N1563_n_19665;
wire n_42309;
wire newNet_3603;
wire n_9611;
wire n_12104;
wire n_15070;
wire n_11014;
wire newNet_515;
wire n_4073;
wire n_35678;
wire n_41566;
wire n_39230;
wire n_18453;
wire n_33155;
wire FE_OCP_RBN3720_n_39913;
wire n_9437;
wire delay_xor_ln22_unr12_stage5_stallmux_q_17_;
wire newNet_3484;
wire n_39616;
wire n_21328;
wire n_36502;
wire n_3731;
wire n_33536;
wire n_42549;
wire FE_OCP_RBN2889_n_46957;
wire n_10239;
wire n_42376;
wire n_32341;
wire n_38704;
wire n_708;
wire FE_RN_1109_0;
wire n_7456;
wire n_16638;
wire newNet_2555;
wire n_16135;
wire newNet_384;
wire n_22465;
wire n_34461;
wire FE_OCP_RBN3406_n_28597;
wire n_37832;
wire n_19553;
wire FE_OCPN988_n_28353;
wire n_21478;
wire n_4696;
wire FE_RN_1616_0;
wire n_28123;
wire FE_OCPN1047_n_24819;
wire n_3711;
wire n_6956;
wire n_9692;
wire n_41860;
wire n_16919;
wire n_40099;
wire n_21183;
wire n_23663;
wire n_18561;
wire n_13532;
wire n_21796;
wire n_11148;
wire n_37297;
wire n_8594;
wire n_9613;
wire n_4294;
wire n_31492;
wire n_17426;
wire n_16125;
wire n_34098;
wire n_41557;
wire n_38767;
wire n_5444;
wire newNet_1463;
wire n_4184;
wire n_11483;
wire n_12;
wire n_7354;
wire n_36216;
wire n_20237;
wire n_1015;
wire n_6116;
wire n_4689;
wire n_1370;
wire n_36439;
wire n_6172;
wire n_13252;
wire delay_xor_ln21_unr3_stage2_stallmux_q_11_;
wire newNet_2668;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_10700;
wire n_567;
wire n_2422;
wire n_11677;
wire n_17289;
wire n_36211;
wire n_25765;
wire n_18351;
wire newNet_734;
wire FE_OCPN3755_n_1451;
wire n_13585;
wire newNet_3297;
wire n_2630;
wire n_35223;
wire n_42526;
wire n_23260;
wire FE_OCP_RBN1687_n_18986;
wire n_17932;
wire n_19479;
wire n_22248;
wire n_27008;
wire n_15883;
wire FE_RN_1097_0;
wire n_26013;
wire n_29554;
wire n_2115;
wire n_28927;
wire n_26884;
wire n_26265;
wire n_43664;
wire n_29946;
wire newNet_1795;
wire n_6476;
wire n_34201;
wire FE_OCP_RBN3802_n_44721;
wire FE_OCP_RBN3541_n_34487;
wire FE_OFN84_n_46137;
wire n_23465;
wire n_42417;
wire n_12885;
wire n_36575;
wire n_30384;
wire n_7445;
wire FE_OCP_RBN2405_n_24638;
wire n_4303;
wire n_26869;
wire n_20750;
wire n_25097;
wire FE_OCP_RBN3854_n_20848;
wire n_766;
wire n_7164;
wire n_16161;
wire newNet_3162;
wire n_36344;
wire n_7935;
wire n_43262;
wire n_40673;
wire n_10925;
wire n_36751;
wire n_11988;
wire n_39188;
wire n_2654;
wire n_38932;
wire n_10669;
wire newNet_1868;
wire n_29591;
wire n_38403;
wire n_41969;
wire n_35334;
wire n_21505;
wire n_29653;
wire n_23546;
wire n_19174;
wire n_15611;
wire newNet_589;
wire n_28602;
wire n_35073;
wire newNet_2025;
wire n_14422;
wire n_5213;
wire n_9435;
wire n_45024;
wire n_1382;
wire n_23873;
wire n_39723;
wire n_13521;
wire n_35704;
wire n_31578;
wire n_38452;
wire n_12470;
wire n_36569;
wire n_28632;
wire newNet_1812;
wire n_21668;
wire n_43223;
wire n_40579;
wire n_28863;
wire n_11611;
wire n_28499;
wire n_25512;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_13_;
wire n_19089;
wire FE_OCP_RBN3856_FE_RN_779_0;
wire n_16543;
wire n_14796;
wire n_5757;
wire n_12423;
wire n_42440;
wire n_2634;
wire n_23429;
wire n_40956;
wire n_12148;
wire n_56;
wire newNet_3176;
wire n_7383;
wire n_2774;
wire n_39869;
wire n_31569;
wire n_28114;
wire n_37220;
wire n_3926;
wire n_35755;
wire n_46221;
wire delay_add_ln22_unr5_stage3_stallmux_q_22_;
wire n_41267;
wire n_18106;
wire n_40723;
wire n_33260;
wire FE_OCP_RBN2463_n_3076;
wire delay_add_ln22_unr8_stage4_stallmux_q_5_;
wire n_37645;
wire n_15306;
wire newNet_3649;
wire n_11293;
wire n_29484;
wire n_42065;
wire n_39257;
wire n_22819;
wire FE_RN_1502_0;
wire n_41743;
wire n_16840;
wire newNet_1372;
wire n_9397;
wire n_34542;
wire n_24465;
wire n_25830;
wire newNet_480;
wire n_12194;
wire n_3525;
wire n_32785;
wire n_13463;
wire n_6590;
wire n_32753;
wire n_7938;
wire n_10138;
wire n_13236;
wire n_15139;
wire delay_xor_ln21_unr9_stage4_stallmux_q_8_;
wire n_1899;
wire n_11307;
wire n_16777;
wire n_13548;
wire newNet_2592;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_5_;
wire n_41282;
wire newNet_1280;
wire n_30160;
wire newNet_1561;
wire n_39775;
wire n_22953;
wire n_7493;
wire n_19363;
wire n_38808;
wire n_29727;
wire newNet_1194;
wire n_19193;
wire n_5206;
wire n_36112;
wire n_32418;
wire n_31737;
wire n_1149;
wire n_18396;
wire n_29747;
wire n_14452;
wire n_42146;
wire FE_OCP_RBN2132_n_40629;
wire n_4549;
wire FE_RN_1435_0;
wire n_2369;
wire n_25628;
wire n_40363;
wire n_39766;
wire FE_RN_163_0;
wire n_6758;
wire n_12320;
wire n_32679;
wire n_30449;
wire n_24043;
wire n_17512;
wire n_29015;
wire n_11962;
wire n_19115;
wire FE_OCP_RBN2647_n_47014;
wire n_23040;
wire n_20424;
wire n_17481;
wire n_28380;
wire n_18774;
wire n_32108;
wire newNet_436;
wire FE_OCP_RBN3584_n_14681;
wire n_40199;
wire n_16818;
wire n_3746;
wire n_43399;
wire n_16851;
wire n_38784;
wire FE_RN_1075_0;
wire n_7484;
wire FE_RN_1569_0;
wire n_43373;
wire n_385;
wire n_29325;
wire n_16261;
wire n_11833;
wire newNet_686;
wire newNet_1490;
wire n_7565;
wire n_43012;
wire n_29165;
wire n_11134;
wire n_36639;
wire n_32174;
wire n_7751;
wire n_27411;
wire n_36989;
wire n_42625;
wire n_4477;
wire n_24194;
wire n_20456;
wire n_23209;
wire FE_RN_1670_0;
wire n_34930;
wire newNet_3358;
wire n_8266;
wire n_15325;
wire FE_RN_1258_0;
wire n_9084;
wire n_16999;
wire n_33753;
wire FE_OCP_RBN2292_n_2438;
wire n_17470;
wire n_7700;
wire n_24023;
wire newNet_250;
wire n_4381;
wire n_15568;
wire n_22658;
wire n_20340;
wire n_46367;
wire n_5478;
wire n_32061;
wire n_16452;
wire n_16301;
wire n_13512;
wire n_39501;
wire n_45118;
wire n_39606;
wire n_22111;
wire n_32968;
wire n_15448;
wire FE_OCPN1493_n_23398;
wire n_15523;
wire FE_OFN737_n_22641;
wire n_5790;
wire n_19860;
wire n_11598;
wire FE_RN_519_0;
wire n_12755;
wire delay_xor_ln21_unr15_stage6_stallmux_q_10_;
wire n_43732;
wire n_7915;
wire newNet_3707;
wire n_6550;
wire n_28301;
wire n_41946;
wire n_22912;
wire FE_OCPN1403_n_21007;
wire n_38298;
wire n_25446;
wire n_18807;
wire n_34170;
wire n_2666;
wire n_42208;
wire n_23473;
wire n_21415;
wire n_8895;
wire n_9124;
wire FE_OCP_RBN3024_n_39942;
wire n_40872;
wire newNet_3591;
wire n_42357;
wire delay_xor_ln21_unr3_stage2_stallmux_q_9_;
wire n_35742;
wire FE_OCP_RBN3092_n_11475;
wire n_15688;
wire n_8612;
wire n_31657;
wire n_11361;
wire newNet_1965;
wire n_9773;
wire n_42934;
wire n_36206;
wire n_6151;
wire n_8570;
wire n_43812;
wire n_9005;
wire n_12256;
wire n_30099;
wire newNet_2176;
wire n_12327;
wire n_21389;
wire n_39545;
wire n_36673;
wire n_26072;
wire n_4867;
wire n_36218;
wire n_545;
wire n_8373;
wire newNet_416;
wire n_24799;
wire n_33630;
wire n_12692;
wire n_27708;
wire n_1303;
wire n_36964;
wire n_20701;
wire n_35541;
wire n_5524;
wire n_21914;
wire FE_OCPN981_n_31961;
wire n_39274;
wire n_31067;
wire n_5610;
wire n_40133;
wire n_23287;
wire n_41701;
wire n_13829;
wire n_5578;
wire n_37136;
wire n_33418;
wire n_6184;
wire n_19153;
wire newNet_2989;
wire n_18820;
wire newNet_989;
wire n_38595;
wire n_11547;
wire n_34674;
wire n_32846;
wire n_30018;
wire n_12698;
wire n_24125;
wire n_21432;
wire n_20859;
wire n_20030;
wire n_11136;
wire n_42481;
wire n_47254;
wire n_40822;
wire FE_RN_266_0;
wire n_20841;
wire n_23925;
wire n_8969;
wire newNet_1912;
wire n_24367;
wire n_2183;
wire n_30869;
wire n_14171;
wire n_14376;
wire newNet_3010;
wire n_27268;
wire FE_OCP_RBN2241_n_44881;
wire n_39457;
wire n_20795;
wire n_41621;
wire n_20896;
wire n_8291;
wire FE_OCP_RBN3085_n_31819;
wire n_43723;
wire n_26202;
wire n_35554;
wire n_27191;
wire n_37580;
wire n_9370;
wire n_43113;
wire n_42801;
wire n_5158;
wire n_36714;
wire n_6526;
wire n_41858;
wire n_27561;
wire FE_OCP_RBN1698_n_19353;
wire n_990;
wire n_25971;
wire newNet_2938;
wire n_28336;
wire n_11144;
wire delay_xor_ln21_unr9_stage4_stallmux_q_18_;
wire n_14426;
wire n_9607;
wire n_33657;
wire FE_OCPN1518_n_26752;
wire n_3315;
wire n_27064;
wire n_39817;
wire n_37897;
wire n_15242;
wire delay_add_ln22_unr20_stage8_stallmux_q_22_;
wire n_35440;
wire n_23160;
wire newNet_2918;
wire FE_RN_458_0;
wire n_13202;
wire FE_OCP_RBN2692_FE_OCPN843_n_3912;
wire n_30077;
wire delay_xor_ln21_unr15_stage6_stallmux_q_14_;
wire n_37723;
wire n_750;
wire n_21643;
wire n_3345;
wire FE_RN_1114_0;
wire n_10213;
wire FE_RN_1853_0;
wire n_11381;
wire FE_OCPN1055_n_14098;
wire n_35690;
wire n_14239;
wire n_18887;
wire FE_OCP_RBN3655_n_15097;
wire n_16661;
wire n_38760;
wire n_35045;
wire n_6376;
wire n_32111;
wire n_1963;
wire n_37410;
wire n_25544;
wire FE_OCPN3794_FE_RN_1789_0;
wire n_7828;
wire n_373;
wire n_25678;
wire n_26311;
wire newNet_727;
wire newNet_19;
wire n_41922;
wire n_5357;
wire n_32588;
wire newNet_2542;
wire n_12630;
wire n_17954;
wire n_43190;
wire n_39644;
wire FE_RN_1152_0;
wire FE_RN_1754_0;
wire n_41789;
wire n_16909;
wire newNet_995;
wire n_36521;
wire n_40169;
wire newNet_2492;
wire n_19159;
wire n_41905;
wire n_41045;
wire newNet_3149;
wire n_25103;
wire n_29860;
wire newNet_1940;
wire n_28192;
wire n_40383;
wire FE_RN_405_0;
wire n_33499;
wire n_22423;
wire FE_OCPN1001_n_45660;
wire n_13725;
wire n_26193;
wire newNet_339;
wire n_39847;
wire n_3735;
wire n_22083;
wire n_31245;
wire n_9078;
wire n_6384;
wire n_2681;
wire n_14132;
wire n_12975;
wire n_7691;
wire n_14527;
wire n_45754;
wire n_21224;
wire n_34087;
wire n_8812;
wire n_20927;
wire n_9546;
wire n_45826;
wire n_33787;
wire n_2529;
wire n_38788;
wire n_12798;
wire newNet_1983;
wire newNet_1778;
wire n_17369;
wire n_8498;
wire n_23639;
wire n_24918;
wire n_40827;
wire FE_OCP_RBN3072_n_43230;
wire n_11108;
wire n_2276;
wire n_26444;
wire newNet_2059;
wire n_25179;
wire n_23448;
wire n_21599;
wire n_22286;
wire newNet_2606;
wire newNet_2437;
wire n_30062;
wire n_1790;
wire n_14908;
wire newNet_2131;
wire n_43903;
wire n_44133;
wire n_3474;
wire newNet_1327;
wire n_37038;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_16_;
wire n_29763;
wire FE_RN_1651_0;
wire n_35429;
wire n_5322;
wire n_46955;
wire n_31838;
wire n_27399;
wire n_9921;
wire n_25576;
wire n_16622;
wire newNet_2396;
wire n_6704;
wire newNet_2883;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_3_;
wire FE_RN_1076_0;
wire n_36959;
wire n_6813;
wire n_4065;
wire n_42955;
wire n_36787;
wire n_34226;
wire n_29838;
wire n_2010;
wire FE_RN_1554_0;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_11_;
wire n_296;
wire n_40243;
wire n_36705;
wire n_12568;
wire FE_RN_1720_0;
wire n_1809;
wire n_2361;
wire n_19377;
wire FE_OCP_RBN2881_n_21272;
wire n_16079;
wire n_35950;
wire n_3723;
wire newNet_312;
wire n_19726;
wire n_28790;
wire n_25843;
wire n_29702;
wire n_27571;
wire n_37274;
wire n_16732;
wire n_6570;
wire n_33420;
wire n_8140;
wire newNet_2677;
wire n_13904;
wire n_23113;
wire FE_OCPN874_n_44672;
wire n_26513;
wire n_11101;
wire n_15976;
wire delay_add_ln22_unr20_stage8_stallmux_q_16_;
wire n_22676;
wire n_15564;
wire n_621;
wire n_12759;
wire n_31318;
wire n_19573;
wire n_972;
wire n_4056;
wire FE_OCP_RBN2205_n_18242;
wire n_1933;
wire n_21006;
wire n_18786;
wire n_4194;
wire n_15462;
wire n_5583;
wire n_1596;
wire n_24960;
wire n_25891;
wire n_27653;
wire n_44165;
wire n_15748;
wire n_42274;
wire newNet_1750;
wire n_15852;
wire n_1298;
wire newNet_1691;
wire n_6624;
wire n_18824;
wire n_29977;
wire n_13222;
wire n_28698;
wire n_47242;
wire n_31893;
wire n_17308;
wire n_19976;
wire n_31032;
wire n_33041;
wire n_3349;
wire n_10725;
wire delay_xor_ln21_unr15_stage6_stallmux_q_1_;
wire n_35778;
wire n_14530;
wire n_15591;
wire n_33521;
wire n_31628;
wire n_42919;
wire n_8322;
wire n_10458;
wire n_4848;
wire newNet_2416;
wire n_9263;
wire n_42473;
wire newNet_797;
wire n_39517;
wire n_15143;
wire n_38524;
wire n_45758;
wire n_31563;
wire n_29154;
wire n_2393;
wire n_42792;
wire n_36167;
wire newNet_2735;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_25_;
wire n_43748;
wire n_41724;
wire n_30494;
wire FE_OFN773_n_46137;
wire newNet_3220;
wire n_38613;
wire n_32411;
wire newNet_3157;
wire n_27202;
wire n_39280;
wire n_13875;
wire n_23299;
wire n_20133;
wire n_236;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_9_;
wire FE_OCP_RBN3444_n_37945;
wire n_7835;
wire n_41509;
wire n_11164;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_6_;
wire n_587;
wire n_27471;
wire n_29568;
wire n_3038;
wire n_33375;
wire n_3272;
wire n_15744;
wire n_3667;
wire n_37524;
wire n_11096;
wire n_28752;
wire FE_OCP_RBN1680_n_33491;
wire newNet_1538;
wire n_1861;
wire n_3306;
wire FE_OCP_RBN3513_n_13960;
wire n_19101;
wire n_2542;
wire n_15670;
wire n_2240;
wire newNet_1287;
wire n_1974;
wire FE_OCP_RBN2357_n_13818;
wire n_4614;
wire n_33186;
wire n_26525;
wire n_41911;
wire n_24613;
wire FE_OFN77_n_4117;
wire n_34335;
wire n_29896;
wire n_29804;
wire n_36250;
wire n_22484;
wire n_43432;
wire n_13044;
wire n_27294;
wire n_7012;
wire newNet_3433;
wire n_1307;
wire n_34347;
wire n_21249;
wire n_21459;
wire n_39002;
wire n_39697;
wire n_930;
wire newNet_1708;
wire n_41791;
wire n_15907;
wire n_5403;
wire newNet_3003;
wire n_1110;
wire n_45309;
wire n_24880;
wire FE_OCP_RBN3090_FE_OCPN1052_n_31674;
wire n_8410;
wire n_39209;
wire n_12710;
wire n_36451;
wire n_86;
wire n_11924;
wire n_17071;
wire n_36945;
wire n_34520;
wire n_42077;
wire n_26410;
wire n_34137;
wire n_1070;
wire newNet_2314;
wire n_19615;
wire n_10043;
wire n_20945;
wire n_18868;
wire FE_RN_318_0;
wire n_21860;
wire n_12119;
wire n_13406;
wire n_31141;
wire newNet_3198;
wire n_17763;
wire newNet_3691;
wire n_11608;
wire n_41353;
wire FE_OCPN1791_n_25044;
wire FE_RN_1625_0;
wire n_3093;
wire n_30562;
wire n_24778;
wire newNet_3689;
wire n_42240;
wire n_43886;
wire n_32028;
wire newNet_2119;
wire FE_OCP_RBN2291_n_2438;
wire FE_RN_1190_0;
wire n_8796;
wire n_2008;
wire n_31542;
wire n_29342;
wire n_41998;
wire n_13215;
wire n_12578;
wire n_27244;
wire n_40586;
wire newNet_61;
wire FE_RN_1414_0;
wire n_28038;
wire n_43404;
wire n_32720;
wire n_42294;
wire newNet_155;
wire n_25469;
wire n_8772;
wire n_43536;
wire n_28158;
wire n_30891;
wire n_43704;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_25_;
wire newNet_1398;
wire n_941;
wire n_34602;
wire n_35307;
wire n_32830;
wire n_16273;
wire n_41362;
wire n_27971;
wire FE_RN_1684_0;
wire n_27467;
wire FE_OCP_RBN3689_n_16146;
wire n_35890;
wire newNet_577;
wire n_74;
wire n_23078;
wire newNet_2143;
wire n_41036;
wire n_15358;
wire n_39268;
wire n_7941;
wire n_43884;
wire n_9368;
wire n_8553;
wire n_28493;
wire n_24624;
wire n_35351;
wire n_29511;
wire n_22172;
wire n_38728;
wire n_1745;
wire n_4322;
wire newNet_459;
wire n_6202;
wire n_24223;
wire n_17397;
wire n_9421;
wire FE_RN_1634_0;
wire n_42165;
wire n_5250;
wire n_10098;
wire n_40761;
wire newNet_1444;
wire n_14016;
wire n_14267;
wire n_33798;
wire n_5063;
wire n_31747;
wire n_18921;
wire FE_OCP_RBN2174_n_37559;
wire n_26929;
wire delay_add_ln22_unr2_stage2_stallmux_q_12_;
wire n_28384;
wire n_11682;
wire n_9687;
wire n_20874;
wire n_32865;
wire n_14230;
wire n_12268;
wire FE_RN_604_0;
wire n_21581;
wire n_40143;
wire n_38545;
wire newNet_70;
wire n_4437;
wire n_17320;
wire FE_RN_306_0;
wire n_5833;
wire n_19997;
wire n_21800;
wire n_5670;
wire n_11516;
wire n_29351;
wire n_719;
wire n_4504;
wire FE_OCP_RBN1326_n_36489;
wire n_15128;
wire n_21588;
wire n_40770;
wire n_16394;
wire n_18496;
wire n_22549;
wire n_43685;
wire n_31003;
wire newNet_1837;
wire n_42562;
wire n_2246;
wire n_20199;
wire n_3636;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_14_;
wire n_30733;
wire n_13032;
wire newNet_2275;
wire n_9808;
wire n_40322;
wire n_10616;
wire newNet_1518;
wire n_39695;
wire n_37481;
wire n_1241;
wire delay_xor_ln22_unr18_stage7_stallmux_q_9_;
wire n_8503;
wire newNet_184;
wire n_11648;
wire n_14699;
wire n_17383;
wire n_35311;
wire n_642;
wire FE_RN_1873_0;
wire n_14621;
wire n_24551;
wire n_28946;
wire n_36308;
wire n_28931;
wire n_13975;
wire newNet_2499;
wire n_11877;
wire n_38710;
wire n_47272;
wire n_7239;
wire n_38926;
wire n_2579;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_3_;
wire FE_RN_1458_0;
wire n_13501;
wire n_37937;
wire FE_OFN757_n_45813;
wire n_10789;
wire n_2880;
wire n_6829;
wire FE_RN_605_0;
wire n_15154;
wire n_1143;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_15_;
wire n_39672;
wire n_1632;
wire FE_OCP_RBN2907_n_16230;
wire n_35001;
wire n_36232;
wire n_22714;
wire n_28557;
wire n_14801;
wire n_34779;
wire n_40580;
wire n_8044;
wire n_2736;
wire n_3232;
wire delay_add_ln22_unr5_stage3_stallmux_q_2_;
wire n_4373;
wire n_17788;
wire n_31416;
wire n_31784;
wire n_371;
wire n_1104;
wire n_7924;
wire FE_OCP_RBN3682_n_26171;
wire n_44798;
wire n_7770;
wire n_43303;
wire n_32905;
wire n_16241;
wire n_40077;
wire n_12175;
wire n_36927;
wire n_4328;
wire n_10397;
wire n_38137;
wire n_22447;
wire n_38557;
wire n_23584;
wire n_16139;
wire n_171;
wire n_36508;
wire n_36635;
wire newNet_2364;
wire FE_RN_1815_0;
wire n_39475;
wire n_5506;
wire n_24742;
wire n_495;
wire n_20414;
wire n_41411;
wire n_43766;
wire n_11437;
wire newNet_2037;
wire n_2586;
wire n_6503;
wire n_29828;
wire n_1880;
wire n_14258;
wire n_32142;
wire n_36263;
wire n_28224;
wire n_21533;
wire newNet_2042;
wire n_27674;
wire n_35397;
wire n_29419;
wire n_3841;
wire newNet_1852;
wire n_39966;
wire n_8243;
wire n_3881;
wire n_21605;
wire n_19214;
wire newNet_1726;
wire n_33934;
wire n_12723;
wire n_32131;
wire n_981;
wire n_31599;
wire n_8118;
wire n_37849;
wire n_824;
wire n_40536;
wire n_4136;
wire n_41470;
wire n_37320;
wire n_28839;
wire n_26991;
wire n_1385;
wire n_18161;
wire n_2692;
wire n_32374;
wire n_23083;
wire n_19275;
wire n_12968;
wire n_5827;
wire n_21938;
wire n_9668;
wire n_9579;
wire n_33601;
wire n_21514;
wire n_12606;
wire n_3082;
wire n_42990;
wire n_42028;
wire n_30786;
wire n_5906;
wire n_38462;
wire n_6419;
wire n_23120;
wire FE_RN_421_0;
wire n_30586;
wire n_5789;
wire n_36259;
wire n_45221;
wire n_31156;
wire n_18099;
wire n_23031;
wire n_20922;
wire n_4171;
wire n_591;
wire FE_OCP_RBN1171_n_13858;
wire n_7897;
wire n_6988;
wire n_23614;
wire n_17029;
wire n_27131;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_16_;
wire n_2690;
wire n_1262;
wire n_7324;
wire n_6025;
wire n_1404;
wire n_4254;
wire n_30321;
wire newNet_3017;
wire FE_OCP_RBN1150_n_17239;
wire newNet_2126;
wire newNet_148;
wire n_17210;
wire n_41233;
wire newNet_3136;
wire FE_RN_474_0;
wire n_9957;
wire n_30923;
wire n_28912;
wire n_21061;
wire n_39894;
wire n_24649;
wire n_4028;
wire n_7471;
wire n_38167;
wire n_31388;
wire n_16035;
wire n_21260;
wire n_29067;
wire n_41711;
wire n_3339;
wire n_32516;
wire n_12363;
wire n_23667;
wire n_13659;
wire n_2658;
wire n_7556;
wire FE_OCPN1505_n_17680;
wire n_17646;
wire FE_OCP_RBN2521_n_8951;
wire FE_OCPN958_n_3951;
wire n_21700;
wire n_17353;
wire newNet_2263;
wire newNet_916;
wire n_15348;
wire n_15987;
wire newNet_2258;
wire n_129;
wire n_32547;
wire n_241;
wire newNet_2301;
wire n_27782;
wire n_40713;
wire FE_RN_980_0;
wire delay_xor_ln21_unr3_stage2_stallmux_q_4_;
wire n_4833;
wire n_24086;
wire n_41944;
wire n_26503;
wire n_25214;
wire n_19676;
wire n_30813;
wire n_34652;
wire n_15928;
wire newNet_79;
wire n_35034;
wire n_8192;
wire n_24787;
wire n_33771;
wire n_40644;
wire n_40406;
wire n_20597;
wire FE_OCPN1000_n_45660;
wire n_34649;
wire n_43482;
wire n_17695;
wire n_5499;
wire n_16118;
wire n_31548;
wire n_30954;
wire n_41776;
wire n_25612;
wire n_10121;
wire n_29965;
wire newNet_2380;
wire n_353;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_27_;
wire n_26573;
wire n_13736;
wire newNet_2007;
wire n_19510;
wire FE_RN_1131_0;
wire FE_RN_1638_0;
wire n_29999;
wire n_20135;
wire n_14161;
wire n_21433;
wire n_2429;
wire n_11440;
wire n_34486;
wire n_28673;
wire n_41599;
wire n_27758;
wire n_26328;
wire FE_OFN754_n_44461;
wire FE_OCPN1445_n_31473;
wire n_41426;
wire n_28404;
wire n_28872;
wire n_3059;
wire n_40857;
wire n_30532;
wire n_6191;
wire newNet_2244;
wire n_23885;
wire n_34264;
wire n_42080;
wire FE_OCPN1794_n_30612;
wire n_15919;
wire n_27805;
wire n_29387;
wire n_12736;
wire n_17941;
wire newNet_2621;
wire n_6153;
wire n_35373;
wire n_42705;
wire n_22262;
wire n_13701;
wire n_34052;
wire n_28665;
wire n_15839;
wire n_23295;
wire n_21103;
wire newNet_1361;
wire n_12078;
wire n_16212;
wire n_24372;
wire n_23363;
wire n_40202;
wire n_16888;
wire n_31090;
wire n_6003;
wire FE_OCP_RBN1350_n_19148;
wire n_5841;
wire n_8912;
wire n_19008;
wire newNet_2812;
wire n_13780;
wire n_46241;
wire n_33388;
wire n_17794;
wire n_44365;
wire newNet_2946;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_18_;
wire n_28543;
wire n_20082;
wire n_40991;
wire n_19252;
wire n_5628;
wire n_18637;
wire n_43283;
wire newNet_3470;
wire n_16335;
wire n_37319;
wire n_2517;
wire FE_OCPN940_n_7712;
wire n_35413;
wire n_37659;
wire n_26128;
wire n_20447;
wire FE_RN_656_0;
wire n_28723;
wire n_809;
wire n_42410;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_3_;
wire newNet_582;
wire n_12655;
wire n_170;
wire n_31297;
wire n_28992;
wire n_43680;
wire n_14050;
wire n_26942;
wire n_6965;
wire n_3944;
wire n_5709;
wire n_40726;
wire n_40316;
wire FE_RN_1782_0;
wire n_26495;
wire n_6318;
wire n_39381;
wire n_29735;
wire n_2686;
wire n_41486;
wire n_15755;
wire n_13915;
wire n_3417;
wire n_40414;
wire n_19728;
wire n_19364;
wire newNet_1757;
wire n_43600;
wire n_27367;
wire n_5644;
wire n_38111;
wire n_17227;
wire n_21404;
wire n_16832;
wire n_39146;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_9_;
wire n_24166;
wire delay_add_ln22_unr8_stage4_stallmux_q_13_;
wire n_38006;
wire n_32903;
wire n_12955;
wire n_31442;
wire n_30557;
wire n_36200;
wire n_15497;
wire n_13930;
wire n_6919;
wire n_22326;
wire FE_RN_780_0;
wire n_14321;
wire n_38965;
wire n_29302;
wire newNet_3333;
wire FE_RN_1013_0;
wire newNet_364;
wire FE_OCP_RBN2509_n_13896;
wire n_29954;
wire n_15664;
wire n_28439;
wire FE_RN_351_0;
wire n_8407;
wire n_34171;
wire n_15750;
wire n_29888;
wire n_43447;
wire n_43055;
wire n_42904;
wire n_34908;
wire n_23897;
wire n_40115;
wire n_30356;
wire n_20223;
wire n_40795;
wire n_27307;
wire n_41819;
wire n_37232;
wire newNet_42;
wire newNet_903;
wire n_30226;
wire FE_RN_1586_0;
wire n_10653;
wire n_631;
wire n_1217;
wire newNet_3236;
wire n_42823;
wire n_28221;
wire n_3406;
wire n_34595;
wire n_11889;
wire n_44566;
wire n_27388;
wire n_12909;
wire n_39313;
wire n_39051;
wire n_13039;
wire FE_OCP_RBN2202_n_12808;
wire n_3595;
wire FE_OCP_RBN2388_n_13860;
wire n_32603;
wire n_42462;
wire n_31415;
wire FE_RN_902_0;
wire n_10352;
wire n_219;
wire n_12115;
wire n_13573;
wire FE_RN_1429_0;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_1_;
wire n_18791;
wire n_4560;
wire n_42655;
wire n_43815;
wire n_1446;
wire n_8539;
wire n_32338;
wire n_20678;
wire newNet_3562;
wire n_46384;
wire n_35805;
wire n_46202;
wire n_4532;
wire n_42201;
wire n_35519;
wire newNet_192;
wire n_42765;
wire n_31197;
wire n_11780;
wire n_2056;
wire newNet_829;
wire n_23973;
wire n_38579;
wire n_34030;
wire n_7181;
wire n_30483;
wire n_9190;
wire n_37388;
wire newNet_3055;
wire n_2950;
wire n_34447;
wire n_23796;
wire n_15274;
wire n_31514;
wire n_42500;
wire FE_OCPN3778_n_36126;
wire n_6857;
wire n_34642;
wire n_15036;
wire n_41356;
wire n_32747;
wire n_24999;
wire FE_OCP_RBN1693_n_19052;
wire n_28059;
wire n_19822;
wire n_13124;
wire n_14272;
wire n_2106;
wire n_20740;
wire FE_OCP_RBN3103_n_32163;
wire n_3329;
wire n_34277;
wire n_21292;
wire n_29409;
wire n_23202;
wire n_4534;
wire n_40593;
wire n_38563;
wire delay_sub_ln23_unr25_stage8_stallmux_q_1_;
wire delay_add_ln22_unr23_stage9_stallmux_q_2_;
wire n_38877;
wire n_13591;
wire n_37449;
wire delay_sub_ln21_unr24_stage9_stallmux_q_4_;
wire n_42421;
wire n_24878;
wire newNet_925;
wire newNet_2382;
wire FE_OCPN1855_n_33341;
wire n_12729;
wire n_33606;
wire n_4445;
wire FE_RN_1090_0;
wire newNet_100;
wire FE_RN_1031_0;
wire n_30972;
wire delay_xor_ln22_unr28_stage10_stallmux_q_0_;
wire n_11323;
wire n_37467;
wire n_8039;
wire n_20489;
wire delay_add_ln22_unr5_stage3_stallmux_q_15_;
wire n_35143;
wire newNet_3421;
wire n_9868;
wire n_23478;
wire n_801;
wire n_35006;
wire n_35187;
wire n_1064;
wire n_3493;
wire n_13248;
wire newNet_3080;
wire newNet_473;
wire n_31706;
wire n_19388;
wire n_23431;
wire newNet_3318;
wire n_32286;
wire n_40049;
wire n_7296;
wire n_9859;
wire n_12640;
wire n_5020;
wire n_34876;
wire n_43395;
wire n_41684;
wire n_42780;
wire n_7424;
wire n_29857;
wire n_19750;
wire n_16437;
wire FE_OCPN1761_n_37877;
wire n_43390;
wire n_32490;
wire n_3494;
wire n_27904;
wire n_8661;
wire n_28050;
wire n_2720;
wire n_40277;
wire n_572;
wire n_20518;
wire n_40500;
wire newNet_3273;
wire newNet_1224;
wire n_29116;
wire n_30088;
wire n_19216;
wire n_7534;
wire n_5293;
wire n_33265;
wire n_35532;
wire n_22872;
wire n_41374;
wire newNet_1735;
wire n_23422;
wire n_18180;
wire n_10324;
wire n_20376;
wire n_20919;
wire newNet_3206;
wire n_3294;
wire newNet_3506;
wire delay_add_ln22_unr2_stage2_stallmux_q_9_;
wire n_38980;
wire n_41408;
wire delay_add_ln22_unr23_stage9_stallmux_q_22_;
wire n_18654;
wire n_17904;
wire n_15715;
wire n_30304;
wire n_17621;
wire n_13824;
wire n_13668;
wire cos_out_11;
wire n_27071;
wire n_9344;
wire n_3605;
wire newNet_1644;
wire n_15316;
wire n_40344;
wire n_39293;
wire n_28748;
wire n_37356;
wire FE_RN_1475_0;
wire n_43409;
wire n_10406;
wire FE_RN_1415_0;
wire newNet_1081;
wire n_9862;
wire n_18536;
wire n_28979;
wire n_29509;
wire newNet_1973;
wire n_39604;
wire n_18913;
wire n_7727;
wire n_10338;
wire n_19806;
wire n_34206;
wire n_10131;
wire n_15537;
wire n_7875;
wire n_35296;
wire n_41091;
wire n_43072;
wire n_39025;
wire n_15415;
wire n_18300;
wire n_37504;
wire n_19338;
wire n_37429;
wire n_37911;
wire FE_RN_1436_0;
wire n_30059;
wire n_2451;
wire n_24713;
wire n_7081;
wire FE_OCP_RBN2234_n_33648;
wire n_39399;
wire n_10255;
wire n_23378;
wire n_9026;
wire n_9785;
wire n_32794;
wire n_28463;
wire n_1686;
wire n_39728;
wire n_30843;
wire n_10141;
wire newNet_3545;
wire newNet_2897;
wire n_8042;
wire n_11689;
wire n_33069;
wire n_27617;
wire n_41573;
wire n_34313;
wire newNet_1247;
wire n_33203;
wire n_32202;
wire n_14864;
wire n_1827;
wire n_4360;
wire n_38216;
wire FE_OCP_RBN2561_n_29819;
wire n_43847;
wire newNet_942;
wire n_5030;
wire FE_OCP_RBN3555_n_44575;
wire beta_4;
wire n_1859;
wire n_17734;
wire n_19422;
wire FE_OCP_RBN3133_n_27736;
wire FE_OCP_RBN3394_n_12504;
wire n_9716;
wire FE_OCP_RBN3265_n_45224;
wire n_34014;
wire n_6963;
wire n_37693;
wire delay_add_ln22_unr14_stage6_stallmux_q_8_;
wire n_34733;
wire n_15298;
wire newNet_1700;
wire n_21137;
wire n_43150;
wire n_30057;
wire n_40059;
wire n_34702;
wire n_44287;
wire n_7793;
wire n_37878;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_30_;
wire n_21473;
wire FE_OCP_RBN2970_n_42896;
wire n_40294;
wire n_34911;
wire n_63;
wire FE_OCP_RBN3493_n_19390;
wire n_20757;
wire n_29023;
wire n_9511;
wire FE_OCPN887_n_42367;
wire FE_RN_527_0;
wire n_6774;
wire n_8822;
wire n_10820;
wire n_42851;
wire n_31189;
wire n_7406;
wire n_40103;
wire n_35432;
wire cos_out_3;
wire n_16449;
wire FE_OCP_RBN1091_n_45224;
wire FE_RN_1084_0;
wire n_37984;
wire newNet_2921;
wire n_24729;
wire FE_OCP_RBN2514_n_8739;
wire newNet_3573;
wire FE_OCP_RBN2837_FE_RN_745_0;
wire n_33462;
wire n_19322;
wire n_41537;
wire n_14153;
wire n_16580;
wire newNet_420;
wire n_2782;
wire n_8881;
wire n_36030;
wire n_15012;
wire n_3905;
wire n_22220;
wire n_22046;
wire newNet_3184;
wire newNet_2830;
wire n_13762;
wire n_40664;
wire n_19524;
wire n_31947;
wire n_21397;
wire n_31519;
wire n_23321;
wire n_35460;
wire newNet_2189;
wire n_12456;
wire FE_OCP_RBN3113_n_32254;
wire n_39398;
wire newNet_165;
wire newNet_1671;
wire n_11498;
wire n_15269;
wire n_35419;
wire newNet_2591;
wire n_14942;
wire n_13335;
wire n_1747;
wire FE_OCP_RBN1188_n_14823;
wire n_34007;
wire n_28016;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_20_;
wire n_36103;
wire n_25035;
wire delay_xor_ln21_unr3_stage2_stallmux_q_0_;
wire n_37264;
wire n_31969;
wire n_18135;
wire n_20039;
wire n_8856;
wire n_26187;
wire n_4402;
wire n_10719;
wire n_23681;
wire n_23957;
wire n_13611;
wire n_12836;
wire n_2374;
wire delay_xor_ln22_unr15_stage6_stallmux_q_6_;
wire n_36671;
wire n_38229;
wire n_41962;
wire n_12890;
wire n_32073;
wire n_28982;
wire n_22886;
wire n_43015;
wire n_19887;
wire newNet_2249;
wire FE_OCPN1428_n_13510;
wire n_22925;
wire n_37417;
wire n_17375;
wire n_34574;
wire n_33427;
wire n_22858;
wire n_29235;
wire n_26227;
wire FE_OFN771_n_46337;
wire FE_OCP_DRV_N1542_n_26125;
wire FE_RN_856_0;
wire FE_OCP_RBN3660_n_15233;
wire n_22901;
wire n_8923;
wire n_16671;
wire n_13883;
wire newNet_1498;
wire n_5886;
wire n_39351;
wire n_21092;
wire FE_RN_48_0;
wire n_35494;
wire n_26566;
wire n_36755;
wire n_19461;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_14_;
wire newNet_3636;
wire n_12580;
wire n_22275;
wire n_41240;
wire n_38314;
wire n_13384;
wire n_12276;
wire newNet_566;
wire n_42556;
wire FE_OCP_RBN2122_n_45224;
wire n_39094;
wire n_2443;
wire n_14932;
wire n_15441;
wire n_5153;
wire n_19637;
wire n_33017;
wire n_16061;
wire newNet_2992;
wire n_5347;
wire n_5358;
wire n_7098;
wire FE_OCP_RBN3648_n_15281;
wire n_33156;
wire n_15211;
wire n_46992;
wire n_32311;
wire newNet_700;
wire n_25231;
wire n_403;
wire n_25687;
wire n_2856;
wire FE_OCPN1792_n_25044;
wire n_6014;
wire n_34924;
wire newNet_1297;
wire n_21054;
wire n_25901;
wire n_9309;
wire n_39377;
wire n_2524;
wire n_18779;
wire n_35324;
wire n_33473;
wire n_46972;
wire n_2404;
wire n_16500;
wire n_29622;
wire delay_xor_ln22_unr9_stage4_stallmux_q_22_;
wire n_17770;
wire n_319;
wire n_40786;
wire n_39736;
wire n_22035;
wire newNet_2446;
wire n_44327;
wire n_9557;
wire n_31521;
wire n_24942;
wire n_26376;
wire n_13994;
wire n_31776;
wire n_15680;
wire n_27834;
wire FE_OCP_RBN3478_n_13756;
wire n_8275;
wire n_33047;
wire n_27120;
wire newNet_2506;
wire cos_out_31;
wire n_38662;
wire n_29272;
wire n_21130;
wire n_25750;
wire n_579;
wire n_23244;
wire n_11659;
wire FE_RN_1078_0;
wire n_33114;
wire n_2410;
wire n_16485;
wire n_1322;
wire n_3124;
wire n_28023;
wire newNet_2198;
wire FE_OCP_RBN2460_n_2818;
wire n_43216;
wire n_17813;
wire n_7640;
wire n_19417;
wire FE_OCP_RBN2815_n_25986;
wire delay_add_ln22_unr5_stage3_stallmux_q_6_;
wire n_40801;
wire n_39925;
wire FE_RN_1828_0;
wire newNet_1422;
wire n_17856;
wire n_8839;
wire n_20421;
wire FE_OCP_RBN1677_n_44847;
wire n_2619;
wire n_36791;
wire n_16863;
wire n_4143;
wire n_37202;
wire n_28321;
wire newNet_3033;
wire n_17882;
wire n_33033;
wire n_8014;
wire n_39156;
wire n_6136;
wire n_45517;
wire n_18197;
wire FE_OCPN1738_n_19052;
wire n_33620;
wire n_18965;
wire n_22525;
wire n_21959;
wire n_11011;
wire FE_OCP_RBN1325_n_29056;
wire n_18682;
wire n_17537;
wire newNet_3559;
wire n_15588;
wire n_41898;
wire n_9605;
wire n_31471;
wire n_5009;
wire FE_RN_966_0;
wire n_5332;
wire n_36775;
wire newNet_1749;
wire n_20400;
wire n_39636;
wire n_7887;
wire n_14102;
wire n_35620;
wire n_8224;
wire n_2135;
wire newNet_3533;
wire n_1978;
wire newNet_2678;
wire n_26615;
wire n_41492;
wire n_20429;
wire FE_RN_1810_0;
wire n_24805;
wire n_10641;
wire n_4782;
wire n_12129;
wire n_42392;
wire n_15029;
wire n_34103;
wire n_9048;
wire n_22696;
wire n_37542;
wire n_10420;
wire n_23405;
wire n_4595;
wire n_23699;
wire n_29800;
wire n_29054;
wire FE_OCPN1245_n_43120;
wire n_6353;
wire FE_OCP_DRV_N1611_n_21706;
wire n_305;
wire n_33572;
wire newNet_113;
wire n_23374;
wire n_9960;
wire n_7262;
wire n_22674;
wire n_19073;
wire n_7025;
wire n_41979;
wire n_32499;
wire newNet_1690;
wire FE_OCPN873_n_44672;
wire delay_xor_ln21_unr6_stage3_stallmux_q_14_;
wire n_37800;
wire n_27568;
wire n_3380;
wire n_4334;
wire n_7332;
wire n_789;
wire n_9206;
wire n_35646;
wire n_32615;
wire n_30102;
wire n_3191;
wire FE_OCP_RBN2468_n_8767;
wire n_918;
wire n_26323;
wire FE_OCPN879_n_31944;
wire n_20902;
wire n_25667;
wire FE_OCP_RBN1987_delay_xor_ln23_unr6_stage3_stallmux_q;
wire n_15625;
wire n_17896;
wire n_41675;
wire n_38931;
wire newNet_1115;
wire n_12938;
wire n_31616;
wire FE_RN_1188_0;
wire n_11004;
wire newNet_331;
wire FE_RN_171_0;
wire n_27591;
wire n_31393;
wire n_16784;
wire n_154;
wire n_10767;
wire n_41957;
wire n_41638;
wire FE_OCP_RBN3678_n_21051;
wire n_17508;
wire FE_OCPN1785_n_30134;
wire n_30917;
wire n_12330;
wire n_30467;
wire n_20337;
wire n_40781;
wire n_29285;
wire n_36551;
wire FE_RN_1751_0;
wire n_24543;
wire n_3901;
wire n_7711;
wire newNet_3059;
wire n_42879;
wire n_2346;
wire n_36004;
wire n_20492;
wire FE_RN_1432_0;
wire FE_OCP_RBN1366_n_20879;
wire n_6700;
wire n_18775;
wire n_528;
wire n_2939;
wire n_447;
wire n_42385;
wire newNet_23;
wire FE_RN_730_0;
wire n_41657;
wire n_40542;
wire n_35388;
wire n_28736;
wire n_37454;
wire n_23549;
wire n_24771;
wire FE_OFN835_n_4333;
wire n_5934;
wire FE_OCP_RBN2203_n_18242;
wire n_1229;
wire n_19318;
wire n_3006;
wire n_12641;
wire n_34202;
wire n_31793;
wire newNet_207;
wire n_2964;
wire n_28113;
wire n_2783;
wire n_16098;
wire n_6487;
wire n_17919;
wire n_6841;
wire n_35464;
wire n_19685;
wire n_38803;
wire n_37555;
wire n_26951;
wire FE_OCP_RBN2679_n_14768;
wire n_12264;
wire n_33890;
wire newNet_204;
wire n_34429;
wire n_9820;
wire n_253;
wire n_4728;
wire n_26231;
wire n_40234;
wire n_9905;
wire n_21172;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_20_;
wire n_13470;
wire n_32023;
wire n_28513;
wire n_35848;
wire n_14488;
wire n_8300;
wire n_20825;
wire n_4452;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_28_;
wire n_21011;
wire n_5388;
wire n_18810;
wire n_18407;
wire newNet_2549;
wire n_25776;
wire n_43146;
wire n_2087;
wire n_32068;
wire n_3756;
wire n_40680;
wire n_9182;
wire n_18554;
wire n_16475;
wire n_39047;
wire FE_RN_1653_0;
wire n_27877;
wire n_15103;
wire FE_RN_1473_0;
wire n_32365;
wire n_4446;
wire n_25565;
wire n_30340;
wire n_23060;
wire n_31350;
wire n_23474;
wire newNet_2925;
wire n_6140;
wire n_167;
wire newNet_1997;
wire n_25201;
wire n_22419;
wire n_23628;
wire FE_OCP_DRV_N1564_n_19665;
wire n_21493;
wire n_42757;
wire n_15604;
wire n_14381;
wire FE_RN_786_0;
wire n_15246;
wire n_369;
wire n_30434;
wire n_28885;
wire n_46968;
wire n_41446;
wire n_691;
wire n_31125;
wire n_23131;
wire FE_OCP_RBN3575_n_4528;
wire n_26089;
wire newNet_3456;
wire n_36080;
wire n_26313;
wire n_24829;
wire FE_RN_1817_0;
wire n_22731;
wire n_24637;
wire n_21578;
wire n_36967;
wire n_28754;
wire n_15215;
wire n_19152;
wire n_8579;
wire n_44346;
wire n_23813;
wire n_2414;
wire n_11208;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_1_;
wire beta_0;
wire n_18092;
wire n_14618;
wire n_6251;
wire FE_OCP_RBN2050_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire n_26354;
wire n_5568;
wire n_44464;
wire n_11047;
wire FE_OCP_RBN3123_n_6557;
wire n_3421;
wire n_19850;
wire n_11882;
wire FE_OCP_RBN1686_n_18986;
wire n_15389;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_13_;
wire n_11389;
wire n_22356;
wire n_42991;
wire n_42074;
wire n_27491;
wire n_6301;
wire newNet_2135;
wire n_17889;
wire n_18445;
wire n_21255;
wire n_43842;
wire delay_xor_ln21_unr18_stage7_stallmux_q_13_;
wire FE_OCPN1743_n_24962;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_4_;
wire n_6180;
wire n_10200;
wire n_26734;
wire n_40067;
wire n_1373;
wire FE_RN_664_0;
wire n_5812;
wire n_8968;
wire n_40187;
wire n_8161;
wire n_17712;
wire n_43033;
wire n_17590;
wire n_36898;
wire n_34784;
wire n_41677;
wire n_36609;
wire n_29431;
wire n_24756;
wire n_7119;
wire delay_xor_ln22_unr3_stage2_stallmux_q_22_;
wire n_30830;
wire n_20118;
wire FE_OCPN1027_n_4182;
wire n_39554;
wire n_38203;
wire n_36601;
wire n_21752;
wire n_9432;
wire newNet_2372;
wire n_6007;
wire newNet_2526;
wire n_43486;
wire n_37890;
wire n_17727;
wire n_3424;
wire n_10388;
wire n_31475;
wire n_14843;
wire n_7644;
wire n_31841;
wire n_30766;
wire FE_RN_650_0;
wire n_32643;
wire n_6295;
wire n_28184;
wire n_22251;
wire newNet_2841;
wire n_1434;
wire delay_xor_ln22_unr6_stage3_stallmux_q_14_;
wire n_34850;
wire n_34460;
wire n_12679;
wire n_8343;
wire n_33878;
wire n_12794;
wire n_42015;
wire newNet_2556;
wire newNet_786;
wire n_26516;
wire newNet_3144;
wire newNet_215;
wire n_36482;
wire n_42308;
wire n_11474;
wire n_39497;
wire n_34290;
wire n_30216;
wire n_35797;
wire n_33061;
wire n_415;
wire n_33991;
wire n_24275;
wire n_34572;
wire FE_RN_1750_0;
wire n_604;
wire n_21597;
wire n_32211;
wire n_39893;
wire FE_RN_1551_0;
wire newNet_1104;
wire FE_RN_1048_0;
wire n_4031;
wire n_40766;
wire FE_OCPN1246_n_43120;
wire newNet_1640;
wire n_29607;
wire n_26903;
wire n_24000;
wire newNet_1215;
wire n_40999;
wire n_7685;
wire FE_OCP_RBN2627_n_14590;
wire n_17654;
wire n_3330;
wire n_39788;
wire n_38474;
wire n_32829;
wire n_32750;
wire n_24578;
wire n_27373;
wire n_21982;
wire n_23438;
wire FE_RN_1127_0;
wire newNet_2158;
wire n_10415;
wire n_17550;
wire n_26559;
wire n_21875;
wire newNet_1172;
wire n_4125;
wire n_13190;
wire n_38969;
wire n_37305;
wire n_13957;
wire newNet_3368;
wire FE_OCPN3747_n_29439;
wire n_9502;
wire n_35909;
wire newNet_2713;
wire n_12720;
wire n_39034;
wire n_21474;
wire n_9170;
wire n_23043;
wire n_2957;
wire n_21449;
wire n_30691;
wire n_12623;
wire FE_RN_817_0;
wire n_39824;
wire n_40173;
wire n_35247;
wire n_29126;
wire newNet_2533;
wire n_17374;
wire n_38953;
wire delay_xor_ln21_unr3_stage2_stallmux_q_27_;
wire n_8692;
wire FE_RN_910_0;
wire n_23366;
wire n_30431;
wire n_463;
wire n_30421;
wire n_33806;
wire n_24646;
wire newNet_2461;
wire n_27678;
wire n_23691;
wire n_32676;
wire n_21641;
wire n_37598;
wire n_9453;
wire n_24627;
wire n_2861;
wire n_38491;
wire FE_RN_1654_0;
wire delay_xor_ln21_unr12_stage5_stallmux_q_9_;
wire n_40702;
wire n_32812;
wire n_25333;
wire n_22064;
wire n_32082;
wire n_11399;
wire FE_OCP_RBN2624_n_3848;
wire newNet_3029;
wire n_23014;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_21_;
wire n_38364;
wire n_20815;
wire n_20027;
wire n_10946;
wire n_38013;
wire n_36531;
wire n_15668;
wire FE_RN_3_0;
wire n_29442;
wire n_23003;
wire n_36022;
wire n_26260;
wire n_41505;
wire n_14300;
wire n_8852;
wire n_6577;
wire n_18992;
wire n_11649;
wire n_37959;
wire n_26836;
wire FE_RN_166_0;
wire n_14598;
wire FE_OCP_RBN2547_n_44944;
wire n_40986;
wire n_15044;
wire n_36917;
wire n_27420;
wire newNet_1828;
wire n_7228;
wire delay_xor_ln22_unr6_stage3_stallmux_q_16_;
wire n_22963;
wire n_26507;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_15_;
wire n_14686;
wire n_12597;
wire newNet_233;
wire n_31279;
wire n_10013;
wire n_9075;
wire n_3228;
wire newNet_1149;
wire n_14896;
wire n_16105;
wire n_37221;
wire n_10209;
wire n_31642;
wire newNet_3013;
wire n_19201;
wire n_32105;
wire newNet_2077;
wire n_26922;
wire newNet_1845;
wire n_29778;
wire n_28718;
wire n_22082;
wire n_40772;
wire n_16349;
wire n_46948;
wire n_39057;
wire n_4806;
wire newNet_3680;
wire n_37956;
wire n_41430;
wire n_29988;
wire n_30186;
wire n_18942;
wire n_13836;
wire n_28344;
wire n_32151;
wire newNet_3391;
wire n_27360;
wire n_9448;
wire FE_RN_1154_0;
wire n_21212;
wire n_9429;
wire n_9568;
wire n_2713;
wire FE_OCP_RBN2554_n_44576;
wire n_14693;
wire FE_OCP_RBN3681_n_26171;
wire n_19556;
wire n_10948;
wire n_28902;
wire n_5696;
wire n_39799;
wire n_29697;
wire n_25822;
wire n_6724;
wire FE_OCP_RBN3342_delay_add_ln22_unr23_stage9_stallmux_q_24_;
wire n_27469;
wire n_32582;
wire newNet_825;
wire n_35431;
wire n_11152;
wire n_39346;
wire n_17178;
wire n_31515;
wire n_41136;
wire n_31097;
wire n_10939;
wire n_13093;
wire n_510;
wire n_3096;
wire n_13623;
wire n_24911;
wire FE_OCP_RBN3388_n_33108;
wire FE_RN_45_0;
wire n_30458;
wire n_41622;
wire newNet_573;
wire n_41104;
wire n_12801;
wire n_16433;
wire n_41216;
wire n_43349;
wire FE_OCP_RBN1159_n_18517;
wire n_26591;
wire n_40335;
wire n_4938;
wire n_4735;
wire n_34888;
wire n_31510;
wire n_31411;
wire n_42815;
wire n_37327;
wire newNet_523;
wire n_28168;
wire n_34015;
wire n_2887;
wire n_12667;
wire n_35405;
wire n_34124;
wire n_36337;
wire n_34077;
wire newNet_664;
wire n_7079;
wire n_5975;
wire n_7583;
wire n_41138;
wire n_40042;
wire n_28592;
wire n_8990;
wire FE_OCP_RBN1186_n_14823;
wire n_42087;
wire n_17283;
wire n_13279;
wire n_3260;
wire n_5472;
wire n_22094;
wire delay_xor_ln21_unr12_stage5_stallmux_q_4_;
wire newNet_855;
wire FE_OCP_RBN2414_n_2922;
wire n_30939;
wire n_20049;
wire n_19560;
wire n_1472;
wire n_8621;
wire n_7048;
wire n_6612;
wire n_36870;
wire n_25471;
wire n_11225;
wire n_2647;
wire n_33213;
wire n_7132;
wire n_3376;
wire FE_OCP_RBN3389_n_33108;
wire n_33318;
wire n_1251;
wire n_29095;
wire n_1664;
wire n_35361;
wire n_34841;
wire n_36043;
wire n_33465;
wire n_27348;
wire n_27576;
wire n_40273;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_28_;
wire n_35226;
wire n_6637;
wire n_12023;
wire n_18617;
wire n_30960;
wire n_6937;
wire n_33849;
wire n_23206;
wire n_27745;
wire n_12046;
wire FE_RN_949_0;
wire n_7252;
wire n_10077;
wire n_6022;
wire n_6943;
wire n_28930;
wire newNet_2449;
wire newNet_3125;
wire n_289;
wire n_4632;
wire n_20621;
wire n_2622;
wire n_23996;
wire n_7377;
wire newNet_1491;
wire FE_OCP_RBN2165_n_28249;
wire n_31718;
wire n_2832;
wire n_6086;
wire n_12182;
wire n_15884;
wire n_8679;
wire n_18708;
wire n_384;
wire n_24734;
wire newNet_3726;
wire n_46166;
wire n_18593;
wire FE_RN_154_0;
wire n_27548;
wire n_21671;
wire n_42132;
wire n_16960;
wire n_28217;
wire newNet_2856;
wire n_17327;
wire n_15266;
wire n_43315;
wire n_21625;
wire n_36929;
wire newNet_673;
wire newNet_328;
wire n_14535;
wire n_6551;
wire newNet_532;
wire FE_OCP_RBN2617_n_44561;
wire n_13887;
wire n_35070;
wire n_5837;
wire newNet_626;
wire n_2823;
wire n_32119;
wire n_14044;
wire n_29337;
wire n_26496;
wire n_11727;
wire n_9165;
wire n_18669;
wire n_17187;
wire newNet_1436;
wire n_36936;
wire n_26967;
wire n_42559;
wire n_31909;
wire FE_RN_1208_0;
wire n_30126;
wire n_28484;
wire FE_OCPN855_n_20367;
wire FE_RN_635_0;
wire n_19166;
wire n_16633;
wire n_33233;
wire newNet_2517;
wire n_5860;
wire n_9852;
wire n_17260;
wire n_210;
wire n_35386;
wire n_18706;
wire n_7053;
wire newNet_739;
wire n_2354;
wire FE_OCP_RBN2811_n_15433;
wire n_44995;
wire n_29397;
wire n_35110;
wire FE_RN_1234_0;
wire delay_xor_ln22_unr9_stage4_stallmux_q_17_;
wire n_36719;
wire FE_OCP_RBN3098_n_17315;
wire n_32996;
wire n_24033;
wire n_32759;
wire FE_OCP_RBN2575_n_34822;
wire n_8930;
wire n_31272;
wire newNet_3066;
wire n_34062;
wire n_33707;
wire n_9882;
wire n_37630;
wire newNet_2226;
wire n_13460;
wire n_37258;
wire n_16728;
wire n_40813;
wire n_13359;
wire FE_OCP_RBN2685_n_38870;
wire n_25630;
wire newNet_375;
wire n_25975;
wire n_43648;
wire n_534;
wire n_15972;
wire n_40225;
wire newNet_1261;
wire n_35059;
wire n_39227;
wire FE_OCP_RBN2835_n_39586;
wire newNet_272;
wire n_46239;
wire n_22877;
wire FE_RN_1643_0;
wire n_17137;
wire newNet_1331;
wire n_14571;
wire n_14059;
wire n_53;
wire n_3248;
wire n_23222;
wire n_7794;
wire n_107;
wire n_7446;
wire newNet_3008;
wire n_25949;
wire n_13402;
wire newNet_2024;
wire n_20227;
wire delay_xor_ln22_unr12_stage5_stallmux_q_4_;
wire newNet_1548;
wire FE_RN_310_0;
wire FE_RN_846_0;
wire n_31329;
wire n_33778;
wire n_16154;
wire n_24992;
wire n_32740;
wire n_4928;
wire n_13448;
wire n_35962;
wire n_37689;
wire n_32387;
wire n_43052;
wire n_35016;
wire n_31743;
wire n_11845;
wire n_32680;
wire n_38573;
wire n_23714;
wire FE_OFN86_n_46137;
wire FE_OCP_RBN2253_n_13017;
wire n_6436;
wire n_43440;
wire n_4076;
wire n_24230;
wire n_37016;
wire n_21816;
wire n_11762;
wire n_26626;
wire n_24219;
wire n_15903;
wire n_43665;
wire n_43517;
wire n_40698;
wire n_18564;
wire delay_add_ln22_unr2_stage2_stallmux_q_24_;
wire n_29476;
wire n_36345;
wire n_26794;
wire n_5852;
wire n_9988;
wire n_773;
wire n_19647;
wire n_43202;
wire n_39291;
wire n_21244;
wire n_27510;
wire FE_OCP_RBN3600_FE_OCPN1243_n_44460;
wire n_22982;
wire FE_OFN823_n_15791;
wire n_24697;
wire n_42091;
wire n_7811;
wire n_23939;
wire n_17920;
wire n_37288;
wire n_33895;
wire n_43495;
wire n_24906;
wire FE_OCP_RBN3087_n_36535;
wire n_12941;
wire newNet_2308;
wire n_7480;
wire n_44139;
wire newNet_74;
wire n_34511;
wire newNet_610;
wire n_5983;
wire n_39640;
wire n_43366;
wire newNet_3677;
wire n_22958;
wire n_41582;
wire n_43251;
wire n_36746;
wire n_23978;
wire n_35560;
wire n_41900;
wire n_13209;
wire n_29939;
wire n_34357;
wire n_33120;
wire FE_OCP_RBN3730_n_31819;
wire n_32460;
wire n_27404;
wire n_30769;
wire n_38746;
wire delay_xor_ln21_unr3_stage2_stallmux_q_8_;
wire n_10461;
wire n_37751;
wire n_38669;
wire n_17873;
wire n_22498;
wire n_42730;
wire n_39634;
wire n_30083;
wire newNet_681;
wire n_23834;
wire n_35724;
wire n_25966;
wire n_33800;
wire n_5891;
wire newNet_2050;
wire n_40975;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_7_;
wire n_41867;
wire n_8261;
wire n_37583;
wire n_7168;
wire n_5275;
wire n_43256;
wire n_24157;
wire n_10928;
wire n_41633;
wire n_20090;
wire delay_add_ln22_unr8_stage4_stallmux_q_17_;
wire delay_xor_ln21_unr15_stage6_stallmux_q_8_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_24_;
wire n_10987;
wire n_19903;
wire n_9491;
wire FE_OCPN972_n_15900;
wire n_20937;
wire n_7803;
wire n_16686;
wire n_21334;
wire n_18309;
wire n_40267;
wire n_8354;
wire n_41015;
wire n_393;
wire n_4913;
wire n_18393;
wire n_25090;
wire newNet_411;
wire n_31610;
wire n_11054;
wire n_38302;
wire n_2047;
wire newNet_1877;
wire n_3213;
wire n_40070;
wire n_1061;
wire n_29650;
wire n_18289;
wire n_2385;
wire n_902;
wire n_23881;
wire n_12191;
wire n_42118;
wire cordic_combinational_sub_ln23_0_unr16_z_0_;
wire n_21736;
wire n_43697;
wire newNet_937;
wire n_29046;
wire n_15288;
wire newNet_2097;
wire newNet_3630;
wire n_38714;
wire newNet_2482;
wire newNet_1529;
wire newNet_1968;
wire n_11894;
wire n_5969;
wire n_11133;
wire delay_xor_ln21_unr12_stage5_stallmux_q_6_;
wire n_28369;
wire n_1903;
wire n_30034;
wire n_10250;
wire n_34212;
wire newNet_3712;
wire n_6080;
wire FE_OCP_RBN3853_n_20848;
wire n_41389;
wire n_16930;
wire n_1928;
wire n_22266;
wire n_18896;
wire n_5107;
wire FE_RN_337_0;
wire n_7958;
wire n_34006;
wire FE_OCP_DRV_N1555_n_19384;
wire n_8128;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_0_;
wire FE_OCP_RBN2465_n_4336;
wire n_11253;
wire n_23551;
wire n_17720;
wire n_20667;
wire n_8182;
wire n_2528;
wire n_36758;
wire n_39062;
wire n_28253;
wire n_9598;
wire newNet_2459;
wire n_37442;
wire n_9723;
wire n_32884;
wire n_6480;
wire n_9152;
wire newNet_956;
wire n_9651;
wire n_18253;
wire n_17855;
wire n_8402;
wire FE_OCP_RBN2392_n_19434;
wire FE_OCP_RBN2322_n_2638;
wire n_21156;
wire n_15834;
wire n_20100;
wire newNet_1377;
wire n_4980;
wire n_9167;
wire n_44219;
wire n_40631;
wire newNet_1531;
wire n_42804;
wire n_46214;
wire n_29834;
wire n_29496;
wire n_43656;
wire n_14666;
wire n_27978;
wire n_9311;
wire n_38126;
wire n_30566;
wire n_34466;
wire n_8350;
wire n_12504;
wire n_19342;
wire FE_RN_939_0;
wire n_43749;
wire n_2040;
wire n_9134;
wire n_37404;
wire n_8098;
wire FE_OCP_RBN2598_n_34388;
wire newNet_484;
wire n_12984;
wire n_34285;
wire n_17379;
wire FE_OCP_DRV_N1575_n_28829;
wire n_42552;
wire n_28611;
wire n_43762;
wire n_18067;
wire FE_OFN5_n_43918;
wire delay_xor_ln22_unr12_stage5_stallmux_q_8_;
wire n_595;
wire n_47236;
wire n_35938;
wire n_12145;
wire n_19171;
wire delay_xor_ln21_unr6_stage3_stallmux_q_8_;
wire n_21502;
wire n_23845;
wire n_35278;
wire newNet_3040;
wire n_1898;
wire n_11308;
wire newNet_1145;
wire n_12098;
wire n_3484;
wire n_43449;
wire newNet_3455;
wire newNet_1597;
wire n_33087;
wire n_23764;
wire n_46419;
wire n_4369;
wire n_10845;
wire n_15612;
wire n_27541;
wire n_25135;
wire n_11699;
wire n_27701;
wire n_8741;
wire newNet_2091;
wire n_5902;
wire n_41117;
wire newNet_1635;
wire n_13167;
wire n_16339;
wire n_22518;
wire n_34992;
wire n_1622;
wire n_35822;
wire newNet_499;
wire n_21563;
wire n_7328;
wire n_15886;
wire newNet_2329;
wire n_35513;
wire n_18385;
wire FE_OCP_RBN2732_n_4219;
wire FE_RN_1364_0;
wire n_1408;
wire n_17745;
wire n_5353;
wire n_24122;
wire n_16230;
wire n_20883;
wire n_19710;
wire newNet_2231;
wire n_39535;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_6_;
wire newNet_2754;
wire n_11288;
wire n_7487;
wire n_27484;
wire n_34682;
wire n_31284;
wire FE_OCP_RBN3047_n_6013;
wire n_38530;
wire newNet_3552;
wire FE_OCP_RBN2476_n_8599;
wire n_28601;
wire n_19038;
wire n_33977;
wire n_31178;
wire n_45216;
wire newNet_911;
wire n_4693;
wire n_41153;
wire n_39997;
wire n_37819;
wire n_33674;
wire n_28630;
wire n_34440;
wire n_21917;
wire n_18883;
wire n_3279;
wire n_18910;
wire n_662;
wire FE_OCP_RBN3520_n_19663;
wire n_43165;
wire FE_OCP_RBN3480_n_13664;
wire n_10564;
wire FE_OCP_RBN3220_n_21358;
wire n_29907;
wire n_43712;
wire n_14916;
wire n_7737;
wire n_21257;
wire n_31320;
wire n_25536;
wire n_25390;
wire newNet_1292;
wire n_25364;
wire n_8006;
wire n_35243;
wire newNet_2538;
wire n_23290;
wire n_1993;
wire n_20123;
wire FE_OCP_RBN3006_n_11087;
wire FE_OCPN1516_n_35367;
wire n_4575;
wire n_43347;
wire n_37847;
wire n_9049;
wire n_40286;
wire n_6362;
wire n_26091;
wire n_18422;
wire n_11582;
wire n_1463;
wire n_39087;
wire n_27041;
wire n_16708;
wire n_39363;
wire n_38942;
wire n_24580;
wire n_10240;
wire n_36157;
wire newNet_441;
wire n_35027;
wire n_3102;
wire n_2097;
wire n_3360;
wire FE_RN_1250_0;
wire n_27830;
wire n_43385;
wire n_21613;
wire newNet_1020;
wire FE_OCP_RBN2886_n_10570;
wire n_8050;
wire n_43474;
wire n_26422;
wire FE_OCP_RBN2163_n_12312;
wire n_14968;
wire n_25452;
wire n_27721;
wire FE_OCP_RBN3642_n_44490;
wire n_15119;
wire n_20960;
wire n_7963;
wire n_14285;
wire n_15572;
wire newNet_843;
wire n_36469;
wire newNet_248;
wire n_7955;
wire n_27917;
wire n_16000;
wire FE_OCP_RBN1177_n_18981;
wire n_27005;
wire n_25018;
wire newNet_3253;
wire n_39617;
wire n_6132;
wire n_18426;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_15_;
wire n_16678;
wire n_6928;
wire n_20975;
wire FE_RN_1874_0;
wire n_28478;
wire n_16386;
wire n_46999;
wire n_45479;
wire newNet_644;
wire n_3868;
wire n_13437;
wire n_3539;
wire n_39731;
wire n_10734;
wire n_9542;
wire n_41854;
wire n_19495;
wire n_7318;
wire n_4376;
wire n_35782;
wire n_39920;
wire n_33223;
wire newNet_760;
wire n_6117;
wire n_16090;
wire n_24348;
wire n_17484;
wire n_17220;
wire n_11327;
wire n_38202;
wire n_17382;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_7_;
wire n_38173;
wire n_25485;
wire n_2192;
wire n_22474;
wire n_3478;
wire n_8932;
wire n_34870;
wire n_6308;
wire n_20208;
wire n_29904;
wire n_1292;
wire n_23719;
wire n_19577;
wire n_33409;
wire n_10932;
wire n_22966;
wire n_34901;
wire n_35161;
wire FE_OCP_RBN2469_n_19806;
wire n_40232;
wire n_13104;
wire n_4300;
wire n_899;
wire n_29616;
wire n_25169;
wire n_2070;
wire n_2419;
wire FE_OCP_RBN2666_n_35207;
wire n_36975;
wire n_113;
wire n_41460;
wire n_42352;
wire n_29571;
wire FE_OCP_RBN2482_n_14326;
wire n_35116;
wire n_33116;
wire n_31499;
wire n_26696;
wire n_33584;
wire newNet_2869;
wire n_41733;
wire n_31180;
wire n_41260;
wire n_38520;
wire n_36984;
wire n_27956;
wire n_19537;
wire n_27418;
wire n_7538;
wire n_31583;
wire n_4087;
wire n_43230;
wire n_8215;
wire n_33965;
wire n_24618;
wire n_846;
wire n_39133;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_9_;
wire n_31242;
wire n_15816;
wire n_11353;
wire n_32955;
wire n_37499;
wire n_11796;
wire n_11425;
wire newNet_706;
wire newNet_2222;
wire n_10894;
wire n_46194;
wire n_10343;
wire n_12923;
wire newNet_1153;
wire n_6471;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_22_;
wire n_7359;
wire n_6802;
wire n_34752;
wire n_33539;
wire n_43024;
wire n_1314;
wire n_13740;
wire n_31691;
wire FE_OCPN888_n_42367;
wire n_1543;
wire n_7217;
wire n_16417;
wire newNet_329;
wire n_17891;
wire n_27090;
wire n_49;
wire n_5195;
wire n_20245;
wire n_41247;
wire newNet_561;
wire n_2764;
wire FE_RN_1531_0;
wire n_23213;
wire FE_RN_1104_0;
wire n_23261;
wire n_5599;
wire n_23197;
wire n_18646;
wire FE_OCP_RBN3205_n_44365;
wire FE_RN_904_0;
wire FE_OCP_RBN2263_n_29033;
wire FE_OCP_RBN2120_n_45224;
wire n_18060;
wire n_26771;
wire n_2603;
wire n_17430;
wire n_24071;
wire n_24628;
wire n_6835;
wire n_12714;
wire n_24462;
wire n_36479;
wire n_123;
wire newNet_1925;
wire n_27942;
wire n_30657;
wire newNet_3625;
wire n_9801;
wire n_33371;
wire n_30013;
wire n_25739;
wire n_17249;
wire n_14437;
wire n_14625;
wire n_945;
wire newNet_1534;
wire n_37153;
wire newNet_3103;
wire n_21548;
wire n_15877;
wire n_91;
wire n_43458;
wire n_14379;
wire FE_OCP_RBN1696_n_19206;
wire n_39213;
wire n_2121;
wire n_25439;
wire n_1820;
wire n_10762;
wire FE_RN_1107_0;
wire n_31936;
wire n_38886;
wire n_42653;
wire n_41640;
wire n_9814;
wire n_34659;
wire n_16044;
wire n_34721;
wire n_9375;
wire FE_OCP_RBN2568_n_8904;
wire n_25379;
wire n_42591;
wire n_18149;
wire n_36395;
wire n_27339;
wire n_18922;
wire n_41619;
wire n_28970;
wire n_798;
wire FE_RN_370_0;
wire n_17230;
wire n_9870;
wire newNet_3106;
wire n_5163;
wire FE_RN_406_0;
wire FE_OCP_RBN2377_n_29480;
wire n_12355;
wire n_2478;
wire FE_OCP_RBN2410_n_13960;
wire FE_OCP_RBN2102_n_44962;
wire n_31835;
wire n_13589;
wire n_12224;
wire n_39592;
wire n_5443;
wire n_7314;
wire n_37347;
wire n_21491;
wire n_42133;
wire n_23522;
wire newNet_2995;
wire n_8382;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_6_;
wire n_4165;
wire newNet_3124;
wire FE_RN_375_0;
wire n_18377;
wire FE_RN_764_0;
wire n_13174;
wire n_89;
wire n_21184;
wire n_13069;
wire n_18015;
wire n_6691;
wire n_32789;
wire newNet_3569;
wire n_17601;
wire n_18519;
wire delay_xor_ln22_unr6_stage3_stallmux_q_11_;
wire n_39605;
wire n_6944;
wire n_5580;
wire n_9803;
wire n_23215;
wire n_5341;
wire n_40797;
wire n_3450;
wire n_41048;
wire n_20201;
wire n_682;
wire newNet_546;
wire n_5901;
wire n_14902;
wire n_4660;
wire n_7421;
wire n_23926;
wire n_23524;
wire n_37518;
wire n_37899;
wire n_25532;
wire n_36700;
wire n_25413;
wire n_37694;
wire n_42650;
wire n_10034;
wire n_37496;
wire newNet_2217;
wire n_8926;
wire n_27283;
wire n_10160;
wire n_41391;
wire n_13615;
wire n_2116;
wire n_45525;
wire n_34554;
wire n_26014;
wire n_16653;
wire n_2821;
wire n_20700;
wire n_10181;
wire n_36974;
wire n_13923;
wire FE_OCP_RBN2117_n_45224;
wire n_17294;
wire n_25242;
wire n_31206;
wire FE_OCP_RBN3695_n_5284;
wire n_36851;
wire FE_OCP_RBN3027_n_39942;
wire n_35407;
wire n_9340;
wire FE_RN_729_0;
wire newNet_627;
wire n_9304;
wire newNet_319;
wire n_32957;
wire n_40341;
wire FE_OCP_RBN3499_n_8187;
wire n_21194;
wire n_4407;
wire n_29555;
wire delay_xor_ln21_unr21_stage8_stallmux_q_2_;
wire newNet_3737;
wire n_40218;
wire n_23985;
wire n_19167;
wire newNet_1773;
wire n_3015;
wire newNet_2494;
wire n_6367;
wire n_2423;
wire n_38044;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_0_;
wire n_41629;
wire n_21098;
wire newNet_3036;
wire n_1674;
wire n_20998;
wire n_25732;
wire n_43320;
wire n_2628;
wire FE_RN_1230_0;
wire n_13599;
wire n_10251;
wire n_1160;
wire n_9819;
wire newNet_3379;
wire n_31324;
wire n_33670;
wire n_26784;
wire newNet_521;
wire n_43013;
wire FE_RN_137_0;
wire n_13379;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_26_;
wire n_33239;
wire newNet_2474;
wire n_10738;
wire n_20192;
wire FE_RN_1120_0;
wire n_23011;
wire n_43275;
wire n_7330;
wire n_19774;
wire n_28664;
wire n_6895;
wire n_41837;
wire n_40978;
wire n_1485;
wire delay_xor_ln21_unr15_stage6_stallmux_q_16_;
wire n_22047;
wire n_34592;
wire FE_OCP_RBN1157_n_18375;
wire FE_OCPN3750_n_44222;
wire n_24346;
wire FE_RN_1676_0;
wire n_16951;
wire n_32231;
wire n_41406;
wire n_39075;
wire n_606;
wire n_21037;
wire n_45879;
wire newNet_2913;
wire n_920;
wire n_158;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_9_;
wire n_6108;
wire n_39308;
wire n_11377;
wire n_21456;
wire newNet_138;
wire n_33424;
wire n_36757;
wire n_13661;
wire n_38416;
wire n_39340;
wire n_2092;
wire n_4680;
wire n_43205;
wire n_19721;
wire n_6272;
wire n_33537;
wire newNet_2843;
wire FE_RN_582_0;
wire n_31347;
wire newNet_607;
wire n_11834;
wire n_35416;
wire n_27346;
wire FE_RN_1425_0;
wire n_6951;
wire n_30335;
wire n_24373;
wire n_16430;
wire n_38963;
wire n_10188;
wire n_45518;
wire newNet_1102;
wire n_2789;
wire n_10791;
wire n_15995;
wire n_7667;
wire n_44610;
wire n_8870;
wire n_8440;
wire FE_OCP_RBN2865_n_39640;
wire n_43441;
wire FE_OCP_RBN3059_n_36515;
wire n_33989;
wire n_20171;
wire n_27728;
wire n_24077;
wire n_43468;
wire n_21327;
wire FE_RN_178_0;
wire n_8272;
wire newNet_1732;
wire newNet_1275;
wire n_12505;
wire n_37949;
wire n_31992;
wire delay_xor_ln22_unr9_stage4_stallmux_q_6_;
wire n_43554;
wire FE_OCP_DRV_N1536_n_12633;
wire n_39899;
wire n_26182;
wire n_513;
wire n_43808;
wire n_5994;
wire n_12309;
wire n_37720;
wire n_8641;
wire FE_OCP_RBN2240_n_44881;
wire n_2175;
wire n_18177;
wire newNet_3446;
wire n_9671;
wire n_20823;
wire n_38127;
wire n_25359;
wire n_23704;
wire n_44275;
wire n_22314;
wire n_11436;
wire n_30535;
wire n_28223;
wire n_31941;
wire n_7368;
wire n_11306;
wire delay_add_ln22_unr27_stage10_stallmux_q_16_;
wire n_2084;
wire FE_OCP_RBN1914_n_20965;
wire n_9172;
wire FE_OCP_RBN3034_n_26842;
wire n_28306;
wire n_14390;
wire newNet_588;
wire n_7033;
wire FE_OCP_RBN3626_n_38870;
wire FE_RN_984_0;
wire n_34765;
wire n_5496;
wire n_38199;
wire n_5149;
wire FE_RN_1455_0;
wire newNet_1954;
wire n_41771;
wire newNet_2377;
wire n_20070;
wire n_27387;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_4_;
wire n_38785;
wire n_5437;
wire FE_RN_1413_0;
wire n_3365;
wire FE_OCP_RBN1356_n_44259;
wire n_35061;
wire n_590;
wire newNet_941;
wire n_20436;
wire n_29115;
wire n_25436;
wire n_17463;
wire n_37888;
wire n_20897;
wire n_24024;
wire n_2386;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_5_;
wire n_29037;
wire n_38510;
wire n_36171;
wire n_12050;
wire n_16496;
wire n_11803;
wire n_22834;
wire n_40809;
wire FE_RN_248_0;
wire n_1415;
wire n_33608;
wire n_35650;
wire n_35297;
wire n_28022;
wire n_36790;
wire n_10652;
wire n_19749;
wire n_25016;
wire n_14539;
wire n_848;
wire n_36676;
wire n_9051;
wire newNet_1423;
wire n_17097;
wire n_17341;
wire FE_OCP_RBN3704_n_26231;
wire n_17436;
wire delay_add_ln22_unr17_stage7_stallmux_q_6_;
wire n_6074;
wire n_23368;
wire n_8023;
wire n_27394;
wire n_27103;
wire n_25680;
wire n_2321;
wire newNet_2064;
wire n_19246;
wire FE_OCP_RBN3533_n_13765;
wire newNet_2970;
wire newNet_2245;
wire n_36483;
wire n_15311;
wire n_20741;
wire n_713;
wire n_6854;
wire n_16531;
wire newNet_3065;
wire n_10793;
wire n_43184;
wire n_37149;
wire newNet_3225;
wire n_9979;
wire n_3640;
wire n_17301;
wire n_16782;
wire newNet_1811;
wire n_9994;
wire n_36503;
wire n_11946;
wire n_13435;
wire n_11763;
wire n_24996;
wire n_35029;
wire n_11976;
wire n_30360;
wire n_21680;
wire n_46246;
wire n_14158;
wire n_39615;
wire FE_OCP_RBN1841_n_20505;
wire n_24966;
wire n_14947;
wire delay_add_ln22_unr17_stage7_stallmux_q_17_;
wire n_2540;
wire n_9140;
wire n_33149;
wire n_20052;
wire n_4323;
wire n_2318;
wire FE_RN_1040_0;
wire n_2166;
wire newNet_752;
wire newNet_2977;
wire n_13083;
wire n_10261;
wire n_23664;
wire n_29483;
wire n_26245;
wire n_41579;
wire n_34079;
wire newNet_1634;
wire n_9396;
wire n_12498;
wire n_21277;
wire n_16174;
wire n_41886;
wire n_37930;
wire n_36205;
wire n_15633;
wire n_20591;
wire n_5587;
wire newNet_3451;
wire newNet_145;
wire n_5291;
wire n_43141;
wire n_17427;
wire n_26870;
wire n_20794;
wire n_7974;
wire n_10847;
wire n_1784;
wire n_5716;
wire FE_OCP_RBN2581_n_3734;
wire n_17585;
wire n_10049;
wire n_7546;
wire n_36715;
wire newNet_1065;
wire n_6241;
wire n_9968;
wire n_33498;
wire n_26663;
wire n_18252;
wire FE_OFN786_n_25834;
wire n_43607;
wire FE_RN_1397_0;
wire n_44842;
wire n_30658;
wire n_17626;
wire n_45073;
wire n_29962;
wire n_36720;
wire n_41910;
wire n_13918;
wire n_33297;
wire newNet_95;
wire n_2906;
wire n_7092;
wire n_12905;
wire n_32943;
wire n_12658;
wire newNet_1865;
wire delay_xor_ln21_unr9_stage4_stallmux_q_9_;
wire n_6239;
wire n_31035;
wire n_8092;
wire newNet_3670;
wire n_5251;
wire n_38328;
wire n_26075;
wire n_31370;
wire n_32247;
wire delay_xor_ln22_unr6_stage3_stallmux_q_2_;
wire n_25615;
wire n_14667;
wire n_29728;
wire n_38627;
wire n_27800;
wire FE_OCP_RBN3405_n_28597;
wire n_45010;
wire n_33703;
wire n_4749;
wire n_6535;
wire n_19810;
wire n_43843;
wire n_40360;
wire n_23037;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_15_;
wire n_35937;
wire n_29957;
wire n_16324;
wire newNet_1195;
wire delay_xor_ln21_unr9_stage4_stallmux_q_16_;
wire FE_OCP_RBN2574_n_34822;
wire n_1847;
wire n_2259;
wire n_45023;
wire delay_xor_ln21_unr18_stage7_stallmux_q_7_;
wire FE_OCP_RBN2210_n_37694;
wire n_39961;
wire n_35511;
wire n_40409;
wire n_28438;
wire n_20138;
wire n_14696;
wire newNet_3719;
wire n_39782;
wire FE_RN_1555_0;
wire n_44828;
wire n_3982;
wire n_38172;
wire n_24600;
wire n_23129;
wire newNet_1754;
wire n_22657;
wire n_37426;
wire n_9271;
wire n_27528;
wire n_15161;
wire newNet_3057;
wire n_6097;
wire n_20618;
wire FE_RN_1832_0;
wire n_39722;
wire n_42717;
wire n_21479;
wire n_4825;
wire FE_OCP_DRV_N1556_n_19384;
wire n_4706;
wire n_46976;
wire n_30067;
wire n_19679;
wire n_22268;
wire n_30866;
wire n_37100;
wire n_41212;
wire n_34753;
wire n_19545;
wire n_10122;
wire n_34646;
wire n_29592;
wire newNet_1948;
wire n_39996;
wire n_40398;
wire n_37736;
wire n_42390;
wire n_32875;
wire n_11352;
wire n_7080;
wire n_30418;
wire n_26873;
wire n_2534;
wire newNet_2455;
wire n_7703;
wire n_23071;
wire n_12368;
wire n_21669;
wire n_11597;
wire n_25184;
wire n_4474;
wire n_12982;
wire n_13013;
wire n_42941;
wire n_34261;
wire n_984;
wire n_834;
wire n_19486;
wire FE_OCP_RBN3595_n_14785;
wire n_35214;
wire n_25778;
wire n_15447;
wire n_20649;
wire n_1020;
wire FE_OCP_RBN1728_FE_RN_1583_0;
wire n_30159;
wire newNet_1794;
wire n_34351;
wire n_30574;
wire n_46967;
wire n_29166;
wire n_12782;
wire n_21207;
wire FE_OCP_RBN2429_n_14018;
wire FE_OCP_RBN2676_n_4061;
wire n_35096;
wire FE_OCP_RBN1207_n_16814;
wire n_40626;
wire n_29475;
wire n_12289;
wire n_19753;
wire n_30155;
wire n_35746;
wire newNet_103;
wire n_31194;
wire n_25963;
wire delay_xor_ln21_unr6_stage3_stallmux_q_21_;
wire n_15284;
wire n_16709;
wire n_16778;
wire n_30221;
wire n_30233;
wire n_27332;
wire FE_RN_826_0;
wire n_16926;
wire FE_RN_848_0;
wire n_21160;
wire n_21707;
wire n_24875;
wire n_13575;
wire n_43153;
wire n_39275;
wire FE_OCP_RBN2500_n_13896;
wire n_21131;
wire n_7720;
wire n_44158;
wire newNet_1445;
wire n_6648;
wire n_11862;
wire n_7232;
wire n_32600;
wire n_38951;
wire n_1685;
wire FE_OCP_RBN3604_n_8981;
wire n_28033;
wire n_23245;
wire n_40598;
wire n_5577;
wire n_2004;
wire n_8751;
wire n_24411;
wire n_26537;
wire FE_OCPN1231_n_42201;
wire n_213;
wire n_42503;
wire n_38282;
wire n_8886;
wire n_40348;
wire n_7186;
wire newNet_1913;
wire n_30800;
wire n_22697;
wire newNet_3510;
wire n_9933;
wire n_42760;
wire n_3159;
wire FE_RN_366_0;
wire n_19980;
wire n_34828;
wire n_36072;
wire n_47009;
wire n_20293;
wire n_30672;
wire newNet_127;
wire n_14194;
wire n_20370;
wire n_7042;
wire n_5333;
wire n_6004;
wire n_19942;
wire n_28877;
wire FE_OCP_RBN2875_n_5082;
wire n_41689;
wire n_22716;
wire n_15395;
wire n_39735;
wire n_44021;
wire n_33795;
wire n_18470;
wire newNet_682;
wire n_2497;
wire n_40226;
wire newNet_1678;
wire n_24904;
wire n_5212;
wire n_19024;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_7_;
wire n_25153;
wire n_39472;
wire delay_xor_ln21_unr15_stage6_stallmux_q_3_;
wire n_36696;
wire n_24752;
wire n_15923;
wire newNet_3500;
wire n_24934;
wire n_17418;
wire FE_RN_443_0;
wire n_35345;
wire n_30139;
wire n_37538;
wire sin_out_22;
wire n_23514;
wire n_14486;
wire n_20912;
wire n_42298;
wire FE_OCP_RBN1980_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire FE_OCP_RBN2961_n_26231;
wire n_23223;
wire FE_RN_401_0;
wire n_23373;
wire n_32161;
wire n_1381;
wire n_314;
wire n_35669;
wire n_6918;
wire n_35467;
wire n_23461;
wire n_40850;
wire n_33363;
wire n_40291;
wire n_18077;
wire n_4107;
wire n_41516;
wire n_41479;
wire n_17823;
wire n_18457;
wire n_7868;
wire n_1148;
wire FE_OCPUNCON1807_n_31435;
wire n_35012;
wire newNet_2358;
wire n_1593;
wire n_22573;
wire n_44692;
wire n_25033;
wire n_10594;
wire n_10015;
wire n_27303;
wire n_16109;
wire newNet_1616;
wire newNet_1291;
wire n_31917;
wire n_3927;
wire FE_OCPN947_n_41382;
wire n_26668;
wire n_36774;
wire FE_OCP_RBN3335_n_44962;
wire n_34102;
wire n_746;
wire n_380;
wire n_31275;
wire n_30480;
wire newNet_2306;
wire n_20673;
wire n_19513;
wire n_11844;
wire n_30383;
wire FE_OCP_RBN3105_n_6358;
wire n_3631;
wire n_19792;
wire n_15610;
wire FE_RN_1220_0;
wire n_20226;
wire n_6145;
wire n_21506;
wire n_7068;
wire n_35722;
wire n_13036;
wire n_34916;
wire n_19896;
wire n_20097;
wire n_17640;
wire n_35484;
wire n_39287;
wire n_10039;
wire n_297;
wire delay_add_ln22_unr20_stage8_stallmux_q_1_;
wire n_33377;
wire n_26262;
wire n_14880;
wire FE_RN_836_0;
wire FE_OCP_RBN1685_n_18986;
wire n_31474;
wire n_42075;
wire n_21827;
wire FE_RN_142_0;
wire n_1234;
wire FE_OCP_RBN2449_n_14114;
wire n_32262;
wire n_5659;
wire n_35426;
wire n_43906;
wire n_7118;
wire n_9494;
wire n_45864;
wire n_29893;
wire n_6621;
wire n_25048;
wire n_13901;
wire FE_OFN764_n_15670;
wire newNet_3243;
wire n_30906;
wire n_9667;
wire n_26548;
wire n_20500;
wire n_41508;
wire n_1449;
wire n_27459;
wire n_5689;
wire n_11420;
wire n_41432;
wire n_33745;
wire n_24569;
wire n_41312;
wire n_26804;
wire newNet_2939;
wire n_883;
wire n_15596;
wire n_40614;
wire n_17176;
wire newNet_1284;
wire n_14557;
wire n_26164;
wire n_25464;
wire n_20160;
wire newNet_2140;
wire n_30625;
wire n_18499;
wire newNet_1896;
wire n_20307;
wire n_16739;
wire n_20950;
wire n_12209;
wire n_15463;
wire n_43300;
wire n_17381;
wire n_28966;
wire n_38635;
wire n_4385;
wire n_8519;
wire n_18663;
wire n_47268;
wire n_17395;
wire n_15397;
wire n_10997;
wire n_3274;
wire newNet_3143;
wire newNet_881;
wire n_39692;
wire n_26362;
wire n_4506;
wire n_42535;
wire n_31259;
wire newNet_868;
wire FE_RN_670_0;
wire n_24726;
wire n_11621;
wire n_12567;
wire n_23208;
wire n_31727;
wire n_17708;
wire n_41768;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_16_;
wire n_24442;
wire FE_RN_1535_0;
wire n_9952;
wire n_33822;
wire n_8848;
wire n_97;
wire n_3262;
wire n_6769;
wire n_12437;
wire n_44775;
wire n_36865;
wire n_10993;
wire n_24633;
wire n_6718;
wire n_33039;
wire n_37715;
wire n_27063;
wire n_26529;
wire n_9843;
wire n_32807;
wire n_1048;
wire n_16523;
wire FE_RN_903_0;
wire newNet_2545;
wire n_2956;
wire n_29821;
wire n_36590;
wire newNet_777;
wire newNet_357;
wire n_27778;
wire n_17862;
wire n_24148;
wire n_9739;
wire n_43531;
wire n_38483;
wire n_36650;
wire n_40246;
wire FE_RN_1687_0;
wire FE_RN_162_0;
wire n_1930;
wire n_28167;
wire n_4634;
wire n_14093;
wire n_41013;
wire n_12712;
wire n_43316;
wire n_39654;
wire n_29243;
wire n_1841;
wire n_13183;
wire n_1267;
wire n_12554;
wire n_42433;
wire n_19773;
wire FE_OCP_RBN2413_n_13960;
wire n_26911;
wire n_3466;
wire n_15534;
wire n_5924;
wire n_2587;
wire n_26604;
wire n_8032;
wire newNet_2272;
wire n_11213;
wire n_26322;
wire n_13412;
wire FE_RN_1228_0;
wire n_35693;
wire newNet_112;
wire n_9750;
wire FE_RN_1453_0;
wire n_36818;
wire n_10214;
wire n_46107;
wire n_36680;
wire n_8799;
wire n_19414;
wire n_24804;
wire n_7439;
wire n_2233;
wire n_25606;
wire n_14404;
wire n_36018;
wire n_43625;
wire n_2159;
wire n_11881;
wire n_23403;
wire n_15675;
wire n_6176;
wire n_4619;
wire n_35390;
wire n_12802;
wire n_9548;
wire n_3687;
wire FE_OCP_RBN2652_n_14684;
wire n_35003;
wire n_2948;
wire newNet_450;
wire n_6069;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_11_;
wire n_41119;
wire n_18970;
wire n_38360;
wire n_42969;
wire n_825;
wire n_22685;
wire n_37781;
wire n_12603;
wire n_15035;
wire n_30474;
wire n_4573;
wire n_37845;
wire n_28906;
wire n_32179;
wire n_38729;
wire n_3666;
wire n_4562;
wire n_21977;
wire newNet_36;
wire FE_RN_1576_0;
wire FE_RN_1722_0;
wire delay_add_ln22_unr2_stage2_stallmux_q_4_;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_5_;
wire n_42064;
wire n_29412;
wire FE_OCPN1421_n_35611;
wire newNet_3704;
wire n_41784;
wire n_13737;
wire newNet_1324;
wire n_28272;
wire n_7257;
wire n_37916;
wire n_25007;
wire n_27741;
wire n_43048;
wire newNet_3240;
wire n_12479;
wire n_9408;
wire n_3087;
wire n_4230;
wire n_14451;
wire n_6332;
wire n_32115;
wire FE_RN_1257_0;
wire n_40520;
wire n_10436;
wire newNet_258;
wire n_15356;
wire n_19588;
wire n_18657;
wire n_1964;
wire n_29787;
wire newNet_1114;
wire n_9550;
wire n_4481;
wire newNet_563;
wire FE_RN_1235_0;
wire n_13508;
wire newNet_303;
wire n_13742;
wire n_25725;
wire n_15510;
wire newNet_2808;
wire n_39989;
wire newNet_82;
wire n_28183;
wire n_7752;
wire n_11571;
wire n_18615;
wire n_45520;
wire newNet_308;
wire n_12143;
wire n_41865;
wire n_13197;
wire n_12681;
wire n_41420;
wire n_34806;
wire n_34044;
wire n_26044;
wire n_6563;
wire n_32537;
wire delay_add_ln22_unr20_stage8_stallmux_q_29_;
wire n_24319;
wire n_16474;
wire n_23519;
wire n_13471;
wire n_3295;
wire n_4886;
wire n_34980;
wire n_28574;
wire n_27961;
wire n_35595;
wire newNet_3131;
wire n_7139;
wire newNet_2957;
wire n_13207;
wire n_24232;
wire newNet_2209;
wire FE_OCP_RBN3826_n_18951;
wire n_23425;
wire n_34527;
wire n_24588;
wire newNet_1201;
wire n_10349;
wire FE_RN_93_0;
wire FE_RN_465_0;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_7_;
wire n_37191;
wire n_27376;
wire n_3061;
wire FE_OFN832_n_18287;
wire FE_OCP_RBN1910_n_20545;
wire n_29335;
wire n_6506;
wire FE_OCP_RBN2192_n_28597;
wire n_19399;
wire n_40467;
wire n_13803;
wire FE_OCP_RBN1297_n_30451;
wire newNet_1129;
wire n_34383;
wire n_3652;
wire newNet_1652;
wire n_39033;
wire n_20511;
wire n_13225;
wire n_7898;
wire n_43774;
wire n_35327;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_24_;
wire n_39908;
wire n_39969;
wire newNet_2186;
wire newNet_2154;
wire n_28952;
wire n_37099;
wire n_23184;
wire newNet_1665;
wire n_22459;
wire n_3875;
wire newNet_998;
wire FE_OCPN1258_n_25353;
wire n_39502;
wire n_14894;
wire n_7923;
wire FE_OCP_RBN3498_n_8187;
wire FE_OCPN1052_n_31674;
wire n_41536;
wire n_32242;
wire n_23587;
wire n_8722;
wire n_41147;
wire n_23619;
wire n_38724;
wire newNet_2460;
wire FE_OCP_RBN2333_n_38446;
wire n_33738;
wire n_28732;
wire n_19535;
wire n_25648;
wire n_43155;
wire n_5099;
wire n_40039;
wire n_7696;
wire n_5806;
wire cos_out_18;
wire n_3369;
wire n_39151;
wire n_2249;
wire n_28143;
wire n_12318;
wire n_34418;
wire FE_OCP_RBN3106_n_22590;
wire n_20926;
wire n_40657;
wire FE_OCP_RBN3721_n_39913;
wire n_9044;
wire n_5893;
wire n_44143;
wire n_30347;
wire FE_OCPN3786_n_22156;
wire n_45329;
wire newNet_957;
wire FE_OCP_RBN3606_n_8981;
wire n_25593;
wire n_21760;
wire n_36634;
wire FE_RN_943_0;
wire n_7870;
wire n_6051;
wire n_39578;
wire n_10574;
wire n_31147;
wire n_23634;
wire n_43335;
wire newNet_3168;
wire n_30297;
wire n_4783;
wire n_336;
wire n_26222;
wire n_15127;
wire n_36937;
wire n_8049;
wire n_6023;
wire n_9230;
wire n_38537;
wire n_19106;
wire n_10405;
wire n_39195;
wire n_16567;
wire newNet_1836;
wire n_6741;
wire newNet_1484;
wire n_32583;
wire n_40306;
wire n_19466;
wire n_11661;
wire FE_RN_1272_0;
wire n_1435;
wire n_35256;
wire n_25069;
wire n_40386;
wire n_36847;
wire n_15267;
wire FE_OCP_RBN3706_n_11146;
wire n_29171;
wire n_28072;
wire n_18986;
wire n_4743;
wire n_9292;
wire n_20776;
wire n_19325;
wire n_25573;
wire n_8316;
wire newNet_1570;
wire n_3312;
wire n_10102;
wire n_39049;
wire n_8126;
wire n_23508;
wire n_1990;
wire n_26366;
wire n_26123;
wire newNet_2125;
wire n_26968;
wire n_17726;
wire n_11125;
wire n_13703;
wire newNet_1879;
wire n_26673;
wire n_27512;
wire n_23412;
wire n_14517;
wire FE_RN_144_0;
wire delay_sub_ln22_unr24_stage9_stallmux_q_7_;
wire n_23496;
wire FE_OCP_RBN3649_n_35169;
wire n_14772;
wire FE_OCP_RBN2796_n_10106;
wire FE_OCP_RBN2503_n_13896;
wire n_17416;
wire n_25991;
wire n_7476;
wire n_30598;
wire n_11654;
wire FE_OCP_RBN2175_n_37559;
wire n_38317;
wire n_7500;
wire FE_OCP_RBN2248_n_13017;
wire n_30104;
wire n_24762;
wire n_12753;
wire n_33853;
wire n_23905;
wire newNet_2880;
wire newNet_2452;
wire newNet_609;
wire n_443;
wire n_31972;
wire n_38713;
wire n_15710;
wire n_23165;
wire n_20169;
wire n_17575;
wire n_21229;
wire n_41037;
wire n_31879;
wire n_13633;
wire n_32152;
wire n_39438;
wire n_29945;
wire n_13724;
wire n_1146;
wire n_27536;
wire n_36786;
wire n_16995;
wire FE_OCP_RBN2675_n_14991;
wire n_5639;
wire n_22998;
wire delay_xor_ln22_unr15_stage6_stallmux_q_7_;
wire n_43827;
wire n_37438;
wire n_16232;
wire n_34742;
wire FE_OCP_RBN2182_n_1916;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_23_;
wire n_10833;
wire n_870;
wire newNet_767;
wire n_9854;
wire n_24429;
wire FE_RN_1858_0;
wire n_5676;
wire n_42262;
wire n_28582;
wire n_9410;
wire n_33574;
wire newNet_1721;
wire n_37326;
wire n_14197;
wire n_34164;
wire n_9261;
wire n_21683;
wire n_39204;
wire n_22725;
wire n_6831;
wire FE_OCP_RBN3011_n_31117;
wire n_42480;
wire n_27657;
wire n_29026;
wire n_7055;
wire n_37249;
wire n_1073;
wire n_11700;
wire FE_OCP_RBN3139_n_40568;
wire n_27864;
wire newNet_2134;
wire n_42998;
wire n_14099;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_10_;
wire n_2352;
wire n_34287;
wire n_23135;
wire n_523;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_24_;
wire FE_RN_383_0;
wire newNet_620;
wire n_2204;
wire FE_OFN751_n_45003;
wire newNet_2201;
wire n_21865;
wire n_9745;
wire n_38764;
wire n_29598;
wire n_11178;
wire n_33927;
wire n_5734;
wire n_32377;
wire sin_out_27;
wire n_36431;
wire n_33970;
wire n_20761;
wire n_10749;
wire n_13650;
wire n_37059;
wire n_33693;
wire n_18848;
wire FE_RN_219_0;
wire newNet_747;
wire n_29232;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_18_;
wire n_39849;
wire n_8810;
wire n_46237;
wire n_22489;
wire newNet_1950;
wire beta_16;
wire n_22784;
wire n_36254;
wire FE_RN_1334_0;
wire FE_OCP_RBN3852_n_20848;
wire n_20660;
wire n_45858;
wire n_6425;
wire n_47186;
wire n_21922;
wire n_22592;
wire FE_OCP_RBN2915_n_42947;
wire n_4759;
wire n_6355;
wire n_22744;
wire n_4138;
wire n_10021;
wire n_16027;
wire n_8303;
wire FE_OCPN1735_n_37877;
wire n_38391;
wire n_15765;
wire n_36407;
wire FE_RN_1422_0;
wire n_32572;
wire n_32497;
wire n_43272;
wire n_41562;
wire newNet_3239;
wire FE_OCP_RBN3357_delay_xor_ln22_unr28_stage10_stallmux_q_0_;
wire n_2918;
wire n_17777;
wire n_19992;
wire n_15970;
wire FE_RN_1573_0;
wire n_41704;
wire n_32070;
wire n_18086;
wire delay_sub_ln23_0_unr22_stage8_stallmux_q;
wire n_36845;
wire n_28070;
wire n_17490;
wire n_11778;
wire n_32022;
wire n_1865;
wire n_31977;
wire n_26447;
wire n_47;
wire n_30375;
wire n_19687;
wire newNet_794;
wire n_47210;
wire n_35577;
wire newNet_2391;
wire n_43264;
wire FE_OCP_RBN3491_n_29553;
wire n_30466;
wire n_36958;
wire n_3434;
wire n_41203;
wire n_45213;
wire n_38895;
wire newNet_3578;
wire n_1916;
wire n_13424;
wire n_14292;
wire FE_RN_818_0;
wire n_37286;
wire FE_OCP_RBN2937_n_16113;
wire n_22507;
wire FE_RN_1373_0;
wire FE_OCPN3185_FE_OCP_RBN1140_n_25816;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_12_;
wire n_39190;
wire n_9881;
wire n_20984;
wire n_23688;
wire n_23749;
wire n_36965;
wire n_738;
wire n_41794;
wire n_39784;
wire n_23863;
wire n_17895;
wire newNet_3461;
wire newNet_1705;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_18_;
wire n_5404;
wire delay_xor_ln22_unr3_stage2_stallmux_q_14_;
wire n_13403;
wire n_26147;
wire n_22851;
wire n_25976;
wire n_39778;
wire n_32482;
wire FE_OCP_RBN3709_n_46337;
wire n_39442;
wire n_25050;
wire n_14606;
wire n_14317;
wire n_4378;
wire n_31744;
wire n_23836;
wire n_22253;
wire newNet_1131;
wire n_15153;
wire n_8289;
wire n_5691;
wire n_37112;
wire n_17660;
wire n_36496;
wire n_25172;
wire FE_RN_945_0;
wire n_23742;
wire n_3185;
wire n_1806;
wire n_3381;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_23_;
wire n_45821;
wire n_7352;
wire n_33397;
wire n_10393;
wire n_1126;
wire newNet_2577;
wire n_44921;
wire n_29803;
wire n_18124;
wire n_13357;
wire n_32500;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_12_;
wire n_40624;
wire n_31074;
wire n_32277;
wire n_28054;
wire n_8587;
wire n_12262;
wire n_43437;
wire newNet_568;
wire n_26627;
wire n_5066;
wire n_41040;
wire n_11801;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_10_;
wire n_13494;
wire n_42732;
wire n_18934;
wire n_1215;
wire n_40080;
wire n_25997;
wire n_15554;
wire n_26522;
wire delay_xor_ln22_unr3_stage2_stallmux_q_9_;
wire n_25142;
wire n_38056;
wire n_36450;
wire n_5579;
wire n_8085;
wire n_1169;
wire n_7515;
wire n_18551;
wire FE_RN_1052_0;
wire FE_RN_609_0;
wire newNet_1039;
wire n_1534;
wire n_33980;
wire n_12924;
wire n_40501;
wire n_25691;
wire n_34576;
wire FE_OCP_RBN3210_n_44365;
wire n_32339;
wire n_26707;
wire n_37165;
wire n_22167;
wire n_33390;
wire n_15052;
wire newNet_804;
wire n_4020;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_28_;
wire n_3514;
wire n_7346;
wire n_22079;
wire n_39896;
wire newNet_1496;
wire n_32401;
wire newNet_3102;
wire FE_OCPN1778_n_37744;
wire n_28233;
wire FE_RN_1034_0;
wire newNet_3142;
wire n_43344;
wire FE_RN_139_0;
wire n_41088;
wire newNet_26;
wire n_43177;
wire n_19160;
wire n_12877;
wire n_16007;
wire n_38166;
wire n_46373;
wire n_12183;
wire n_27953;
wire n_35591;
wire newNet_3195;
wire n_2849;
wire n_41124;
wire FE_RN_1522_0;
wire n_37582;
wire n_39928;
wire n_31063;
wire n_18717;
wire n_32776;
wire newNet_2185;
wire FE_OCP_RBN3013_n_31117;
wire n_36540;
wire n_17454;
wire n_26390;
wire n_39245;
wire n_4641;
wire n_11418;
wire n_37011;
wire newNet_1480;
wire n_9858;
wire n_38085;
wire n_5550;
wire n_35588;
wire n_159;
wire n_29440;
wire n_46427;
wire n_27918;
wire n_36692;
wire n_29777;
wire n_38663;
wire n_42058;
wire n_3785;
wire n_18658;
wire n_38605;
wire n_4589;
wire n_10965;
wire n_37308;
wire FE_OFN750_n_45003;
wire n_13397;
wire n_11384;
wire n_3769;
wire n_22293;
wire n_32627;
wire n_10740;
wire FE_OCP_RBN2708_n_15135;
wire n_6101;
wire newNet_3558;
wire n_2021;
wire n_23194;
wire n_25277;
wire n_31574;
wire n_3615;
wire n_6125;
wire n_1628;
wire n_35941;
wire n_41193;
wire n_38774;
wire n_26419;
wire n_17835;
wire n_7078;
wire n_6932;
wire n_1548;
wire n_37322;
wire n_35132;
wire n_36223;
wire n_31713;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_17_;
wire n_26008;
wire n_33447;
wire n_1181;
wire n_2245;
wire n_15113;
wire n_33232;
wire n_424;
wire n_19463;
wire n_20113;
wire newNet_3517;
wire n_5184;
wire n_21676;
wire n_14092;
wire n_9653;
wire n_32915;
wire newNet_2751;
wire n_41749;
wire n_33058;
wire n_6904;
wire n_30521;
wire n_23997;
wire n_36475;
wire n_22513;
wire n_5234;
wire n_36565;
wire n_23735;
wire FE_OCP_RBN1196_n_30926;
wire n_9699;
wire n_31778;
wire n_21353;
wire n_7326;
wire n_2617;
wire n_7680;
wire n_40191;
wire n_5267;
wire FE_RN_1289_0;
wire n_17684;
wire n_19769;
wire n_23867;
wire n_9624;
wire newNet_446;
wire newNet_762;
wire newNet_1189;
wire n_30256;
wire n_15294;
wire n_21967;
wire n_10891;
wire n_6528;
wire n_4957;
wire n_45134;
wire n_161;
wire n_24981;
wire n_34551;
wire n_29513;
wire n_15180;
wire n_18746;
wire n_37127;
wire n_14791;
wire n_36733;
wire n_5241;
wire n_41007;
wire n_4866;
wire n_12066;
wire n_23232;
wire n_28256;
wire FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire n_23122;
wire n_32815;
wire FE_OCP_RBN3554_n_44575;
wire n_3111;
wire n_31169;
wire n_6111;
wire n_1516;
wire n_10805;
wire n_8120;
wire n_21741;
wire n_16286;
wire newNet_1788;
wire n_3483;
wire newNet_3260;
wire n_29276;
wire delay_add_ln22_unr23_stage9_stallmux_q_24_;
wire n_26169;
wire n_31231;
wire n_4099;
wire n_518;
wire n_36689;
wire n_27496;
wire n_35271;
wire n_5425;
wire n_23322;
wire n_17722;
wire n_24117;
wire n_40378;
wire n_13130;
wire n_4113;
wire n_22010;
wire n_25760;
wire n_32629;
wire n_38830;
wire FE_OCP_RBN3654_n_10100;
wire n_24425;
wire n_45301;
wire n_10954;
wire n_28386;
wire n_36351;
wire n_13306;
wire n_7145;
wire n_17489;
wire n_23723;
wire n_28986;
wire n_5786;
wire n_40662;
wire n_11055;
wire n_9795;
wire n_16001;
wire n_14617;
wire n_220;
wire n_19331;
wire n_34747;
wire n_250;
wire n_36347;
wire n_9345;
wire n_11465;
wire n_26236;
wire n_8367;
wire n_17478;
wire newNet_1890;
wire n_6138;
wire n_17348;
wire n_24691;
wire delay_sub_ln22_unr24_stage9_stallmux_q_0_;
wire n_32487;
wire n_30477;
wire n_15331;
wire newNet_410;
wire n_19129;
wire n_23989;
wire n_32651;
wire n_13354;
wire FE_OCP_RBN3421_n_12879;
wire beta_5;
wire n_30422;
wire n_19347;
wire newNet_3048;
wire n_17782;
wire delay_add_ln22_unr14_stage6_stallmux_q_17_;
wire n_32895;
wire n_34020;
wire n_19071;
wire n_32454;
wire n_9003;
wire n_40484;
wire n_9352;
wire n_11246;
wire n_42336;
wire newNet_2660;
wire FE_RN_1452_0;
wire n_14783;
wire n_27089;
wire FE_RN_1101_0;
wire n_12230;
wire n_1357;
wire n_45531;
wire n_17385;
wire n_4599;
wire n_19097;
wire n_41730;
wire n_38547;
wire cos_out_6;
wire FE_OCP_RBN1190_n_14911;
wire n_39571;
wire n_5528;
wire n_17887;
wire n_30806;
wire n_2518;
wire n_28933;
wire n_4152;
wire n_15872;
wire FE_OCPN846_n_4046;
wire FE_OCP_RBN2318_n_2367;
wire n_25113;
wire n_12811;
wire n_21835;
wire n_15786;
wire FE_RN_1768_0;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_4_;
wire n_6960;
wire n_43278;
wire newNet_585;
wire n_33607;
wire n_13134;
wire FE_OCPN1390_n_9220;
wire n_6877;
wire n_35828;
wire n_33660;
wire n_31754;
wire n_14663;
wire n_19532;
wire n_5874;
wire n_18244;
wire n_16941;
wire n_40693;
wire n_24342;
wire n_1086;
wire n_43585;
wire FE_OCP_RBN2872_n_39542;
wire n_40495;
wire n_34143;
wire FE_RN_502_0;
wire newNet_1220;
wire newNet_924;
wire n_27909;
wire n_10827;
wire n_25064;
wire n_27002;
wire n_43363;
wire n_41211;
wire n_35670;
wire n_36623;
wire n_20252;
wire n_24560;
wire n_20079;
wire n_20440;
wire n_5364;
wire delay_xor_ln21_unr21_stage8_stallmux_q_6_;
wire n_29498;
wire n_18452;
wire n_43287;
wire n_19434;
wire n_42203;
wire n_23603;
wire FE_OCP_RBN2691_FE_OCPN843_n_3912;
wire n_5650;
wire n_4269;
wire n_41903;
wire n_12341;
wire n_93;
wire FE_OCPN1234_n_2414;
wire n_30492;
wire newNet_554;
wire n_20598;
wire n_20396;
wire n_42272;
wire n_40117;
wire n_27893;
wire FE_OCP_RBN2866_n_39640;
wire n_3218;
wire n_28822;
wire n_40652;
wire n_43863;
wire n_24272;
wire n_34033;
wire n_10413;
wire n_37090;
wire n_17476;
wire n_9985;
wire n_36954;
wire n_34363;
wire n_14060;
wire n_34306;
wire n_24163;
wire newNet_3147;
wire n_28451;
wire n_33202;
wire n_16591;
wire newNet_3256;
wire n_37253;
wire n_13597;
wire newNet_3423;
wire newNet_1082;
wire n_7292;
wire n_42079;
wire n_40393;
wire n_22405;
wire n_16723;
wire n_31055;
wire n_14956;
wire n_1639;
wire n_10493;
wire newNet_615;
wire n_18401;
wire n_26340;
wire n_43424;
wire n_19625;
wire newNet_2518;
wire n_41400;
wire n_37558;
wire n_15807;
wire n_1503;
wire n_39404;
wire n_34475;
wire n_20080;
wire n_16642;
wire n_22438;
wire n_42657;
wire newNet_349;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_27_;
wire n_36382;
wire n_37337;
wire n_46155;
wire n_42234;
wire FE_OCP_RBN3563_n_29857;
wire n_26115;
wire n_37463;
wire n_13112;
wire n_25940;
wire n_30861;
wire n_21063;
wire n_40460;
wire n_25635;
wire n_30428;
wire n_19528;
wire n_10718;
wire n_20328;
wire n_30328;
wire n_39845;
wire n_15975;
wire newNet_1307;
wire n_17627;
wire n_20930;
wire n_7416;
wire n_43641;
wire newNet_567;
wire newNet_1860;
wire n_37448;
wire n_13272;
wire newNet_3651;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_24_;
wire n_12940;
wire n_28174;
wire n_40732;
wire n_19823;
wire n_26946;
wire n_35749;
wire n_7486;
wire n_22133;
wire n_20271;
wire n_45739;
wire n_31305;
wire n_17497;
wire n_7097;
wire n_38090;
wire FE_OCP_RBN3636_n_47260;
wire n_22951;
wire delay_add_ln22_unr17_stage7_stallmux_q_20_;
wire n_7610;
wire n_10041;
wire n_20128;
wire n_17217;
wire n_14658;
wire FE_RN_1322_0;
wire n_39588;
wire n_35245;
wire FE_OCP_RBN2385_n_8342;
wire n_42098;
wire n_17226;
wire n_38883;
wire n_10661;
wire FE_OCP_RBN3370_n_32436;
wire newNet_1588;
wire n_10938;
wire n_16414;
wire n_32405;
wire n_7499;
wire FE_OCP_RBN2908_n_26173;
wire newNet_2628;
wire n_16837;
wire n_38865;
wire n_21405;
wire n_20662;
wire n_3904;
wire n_38720;
wire n_90;
wire n_33255;
wire n_30991;
wire n_41385;
wire n_18601;
wire newNet_2614;
wire FE_RN_1506_0;
wire n_8535;
wire newNet_9;
wire n_24088;
wire n_781;
wire n_3351;
wire n_43824;
wire n_17156;
wire n_12948;
wire newNet_2608;
wire n_32218;
wire FE_RN_1091_0;
wire n_21106;
wire n_35275;
wire n_42178;
wire newNet_3403;
wire n_27941;
wire n_1559;
wire n_29839;
wire n_8961;
wire FE_RN_410_0;
wire n_30889;
wire n_13203;
wire n_39478;
wire FE_OCP_RBN1913_n_20965;
wire n_34001;
wire n_34882;
wire n_33708;
wire n_33179;
wire n_30010;
wire n_46420;
wire n_16810;
wire n_508;
wire n_35157;
wire n_8150;
wire FE_OCP_RBN2947_n_10722;
wire n_14707;
wire n_36727;
wire n_40802;
wire newNet_1960;
wire FE_OCP_RBN2659_n_4101;
wire n_32175;
wire n_23482;
wire n_43659;
wire n_42167;
wire n_15619;
wire n_8181;
wire n_19605;
wire newNet_2983;
wire n_19798;
wire n_25281;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_26_;
wire n_15040;
wire n_16848;
wire n_12003;
wire n_43062;
wire n_16318;
wire n_46388;
wire n_6967;
wire n_10246;
wire n_4502;
wire n_25543;
wire n_19490;
wire FE_RN_926_0;
wire n_27070;
wire n_18899;
wire n_18398;
wire n_27700;
wire FE_OCP_RBN2279_n_24199;
wire n_10693;
wire n_35874;
wire n_36463;
wire n_29938;
wire n_9254;
wire FE_RN_1660_0;
wire n_39332;
wire n_25120;
wire n_18439;
wire n_25160;
wire n_28694;
wire n_42666;
wire n_9404;
wire n_6776;
wire newNet_430;
wire n_20553;
wire n_23468;
wire newNet_965;
wire n_31025;
wire n_34961;
wire n_14075;
wire n_18563;
wire n_12491;
wire FE_RN_811_0;
wire newNet_3502;
wire n_40902;
wire n_34616;
wire n_44354;
wire n_23792;
wire n_18947;
wire n_1767;
wire n_3133;
wire n_32713;
wire n_13018;
wire n_37745;
wire n_30060;
wire n_37638;
wire n_10612;
wire n_18645;
wire n_41241;
wire newNet_3284;
wire n_37317;
wire n_44710;
wire delay_add_ln22_unr8_stage4_stallmux_q_24_;
wire FE_RN_1524_0;
wire n_30957;
wire n_22085;
wire n_6192;
wire n_33322;
wire n_22655;
wire n_36707;
wire n_1466;
wire n_30286;
wire n_17547;
wire n_42494;
wire n_27365;
wire n_31296;
wire n_14924;
wire n_30987;
wire n_29831;
wire n_23201;
wire n_35218;
wire n_15440;
wire n_19078;
wire n_26900;
wire n_40646;
wire n_27481;
wire n_10573;
wire n_14045;
wire n_13860;
wire n_14609;
wire n_13046;
wire n_22263;
wire n_12095;
wire n_33303;
wire n_5236;
wire n_16499;
wire n_13481;
wire newNet_3365;
wire newNet_703;
wire newNet_1693;
wire n_39298;
wire n_20381;
wire n_36281;
wire n_8858;
wire n_31396;
wire FE_OCP_RBN2890_n_10568;
wire n_24451;
wire n_27637;
wire n_2143;
wire n_12838;
wire FE_OCPN975_n_46956;
wire n_24913;
wire n_27884;
wire FE_OCPN1790_n_18119;
wire n_42029;
wire newNet_2;
wire n_12607;
wire FE_OCP_RBN3566_n_29857;
wire n_37200;
wire n_4776;
wire n_22284;
wire n_39956;
wire n_3049;
wire FE_RN_1657_0;
wire n_24705;
wire newNet_1579;
wire n_25813;
wire n_32545;
wire n_19767;
wire n_9964;
wire FE_RN_1144_0;
wire n_16178;
wire n_26834;
wire n_5416;
wire n_25537;
wire n_24013;
wire n_27545;
wire FE_OFN759_n_45813;
wire n_10681;
wire n_1106;
wire n_12334;
wire n_22849;
wire n_39482;
wire n_34518;
wire n_30921;
wire n_13284;
wire n_4003;
wire n_16458;
wire n_8254;
wire n_40526;
wire n_6485;
wire n_36414;
wire n_41109;
wire n_11157;
wire n_15640;
wire n_22640;
wire n_21639;
wire FE_RN_464_0;
wire n_5862;
wire n_22581;
wire n_31374;
wire n_14363;
wire n_36286;
wire n_24767;
wire FE_OFN821_n_4632;
wire n_19208;
wire n_41234;
wire n_29508;
wire n_4374;
wire n_6496;
wire newNet_3091;
wire n_31682;
wire newNet_492;
wire newNet_2333;
wire FE_RN_1133_0;
wire n_2075;
wire n_43899;
wire n_46943;
wire n_13274;
wire n_11925;
wire FE_OCP_RBN2313_n_41420;
wire n_23085;
wire n_20861;
wire n_24005;
wire n_40996;
wire newNet_1295;
wire n_29762;
wire n_5725;
wire FE_RN_438_0;
wire n_36753;
wire n_35940;
wire n_4590;
wire n_22945;
wire FE_OCP_RBN1718_n_20090;
wire n_2673;
wire n_28802;
wire FE_OCP_RBN3026_n_39942;
wire n_32763;
wire FE_OCP_RBN2778_n_15595;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_23_;
wire n_20567;
wire n_42604;
wire n_19186;
wire n_8514;
wire n_30141;
wire n_22236;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_3_;
wire n_1797;
wire n_12815;
wire n_40837;
wire FE_OCPN896_n_44776;
wire n_15937;
wire n_8433;
wire n_20655;
wire n_28599;
wire n_31782;
wire n_27358;
wire n_2627;
wire n_38179;
wire FE_OCP_RBN1843_n_20910;
wire n_37953;
wire newNet_2339;
wire n_1451;
wire n_3144;
wire n_41525;
wire FE_OCP_RBN2366_n_24372;
wire n_9143;
wire n_16970;
wire n_42009;
wire n_17560;
wire n_32133;
wire FE_OCP_RBN2609_n_3807;
wire delay_add_ln22_unr2_stage2_stallmux_q_5_;
wire delay_add_ln22_unr5_stage3_stallmux_q_23_;
wire newNet_1169;
wire n_7007;
wire n_5663;
wire n_29459;
wire n_17785;
wire n_20423;
wire FE_RN_1550_0;
wire n_3967;
wire FE_OCPN984_n_25210;
wire n_20099;
wire n_11991;
wire n_29082;
wire n_17754;
wire n_32826;
wire FE_OCP_RBN2430_n_14018;
wire n_24189;
wire n_11380;
wire FE_OCP_RBN3536_n_13765;
wire n_5889;
wire n_37119;
wire FE_RN_1620_0;
wire n_28029;
wire n_17633;
wire n_19958;
wire n_9010;
wire n_17262;
wire FE_OCP_RBN2497_n_8835;
wire n_36292;
wire n_43307;
wire n_29096;
wire n_36454;
wire FE_OCP_RBN2744_n_15319;
wire n_19599;
wire n_29612;
wire n_21750;
wire n_42845;
wire n_30676;
wire newNet_2942;
wire n_35859;
wire n_19799;
wire n_26106;
wire n_33370;
wire n_25157;
wire FE_OCP_DRV_N1603_n_19961;
wire n_43591;
wire n_3039;
wire n_12035;
wire n_10385;
wire n_23329;
wire n_12542;
wire FE_OCP_RBN1838_n_19528;
wire n_5824;
wire n_5698;
wire n_41272;
wire n_30895;
wire n_26297;
wire n_17953;
wire n_9367;
wire n_21136;
wire n_7372;
wire n_8689;
wire n_20298;
wire n_16389;
wire FE_OFN776_n_17093;
wire n_8790;
wire n_16446;
wire newNet_2002;
wire n_6934;
wire n_7603;
wire n_28228;
wire n_25457;
wire n_30698;
wire n_20642;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_17_;
wire n_37903;
wire newNet_299;
wire n_33773;
wire n_20013;
wire newNet_164;
wire n_2119;
wire n_7805;
wire FE_RN_483_0;
wire n_33316;
wire n_42772;
wire n_41060;
wire n_6654;
wire n_12435;
wire n_26218;
wire n_19738;
wire n_41145;
wire n_42210;
wire n_16093;
wire n_8652;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_15_;
wire n_21870;
wire n_14348;
wire newNet_3158;
wire n_76;
wire FE_OCP_RBN2805_n_30534;
wire FE_OCPN1009_n_28439;
wire n_17647;
wire n_40330;
wire FE_RN_420_0;
wire n_27336;
wire n_40788;
wire n_21769;
wire n_37228;
wire newNet_2550;
wire n_9895;
wire FE_RN_1043_0;
wire n_23159;
wire n_9753;
wire n_19004;
wire n_38955;
wire n_19285;
wire n_19635;
wire n_36778;
wire delay_add_ln22_unr17_stage7_stallmux_q_9_;
wire n_27955;
wire n_5685;
wire n_46348;
wire newNet_1212;
wire n_1754;
wire n_26721;
wire n_19974;
wire n_14026;
wire FE_OCP_RBN3272_n_45224;
wire FE_RN_279_0;
wire n_4451;
wire n_33481;
wire newNet_519;
wire newNet_537;
wire n_25270;
wire n_24986;
wire n_43684;
wire n_31379;
wire n_31639;
wire newNet_2895;
wire n_34601;
wire n_11228;
wire n_9559;
wire n_17440;
wire n_15870;
wire n_8591;
wire n_31509;
wire n_9867;
wire n_38470;
wire n_22802;
wire n_16065;
wire n_1825;
wire FE_OCP_RBN2498_n_8835;
wire n_18893;
wire n_33367;
wire n_10982;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_2_;
wire n_36050;
wire n_12016;
wire n_26755;
wire cordic_combinational_sub_ln23_0_unr12_z_0_;
wire n_18953;
wire n_24312;
wire n_33809;
wire n_3876;
wire n_3624;
wire n_9563;
wire n_12299;
wire n_21153;
wire n_42754;
wire n_3803;
wire n_946;
wire n_7050;
wire n_38614;
wire FE_RN_931_0;
wire n_15502;
wire n_27878;
wire FE_OCP_RBN3003_n_10805;
wire n_25715;
wire n_37396;
wire n_21305;
wire n_17962;
wire n_21813;
wire n_31128;
wire n_2250;
wire n_8620;
wire n_38540;
wire n_12352;
wire n_42108;
wire n_17211;
wire FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_22173;
wire n_33210;
wire n_35259;
wire n_19906;
wire n_20604;
wire n_31017;
wire n_10237;
wire n_6661;
wire n_32208;
wire n_3009;
wire n_43145;
wire n_1947;
wire n_41157;
wire n_37865;
wire n_2090;
wire n_1205;
wire n_12591;
wire n_31103;
wire n_14950;
wire n_9441;
wire n_9908;
wire newNet_3056;
wire n_27470;
wire n_10109;
wire n_30379;
wire n_15491;
wire n_2237;
wire n_11315;
wire n_35080;
wire newNet_2468;
wire n_35649;
wire newNet_3234;
wire n_10028;
wire n_39433;
wire n_38494;
wire n_35735;
wire n_17160;
wire FE_RN_319_0;
wire n_13568;
wire n_42128;
wire n_29228;
wire n_3863;
wire n_27068;
wire n_11262;
wire n_20876;
wire n_3942;
wire n_12059;
wire n_26745;
wire n_10541;
wire n_17759;
wire FE_OCP_RBN1848_n_22068;
wire n_42582;
wire n_34906;
wire newNet_3007;
wire n_11729;
wire newNet_3120;
wire newNet_1931;
wire n_6219;
wire n_19680;
wire FE_OCP_RBN1181_n_19726;
wire n_43431;
wire newNet_2930;
wire n_12269;
wire n_45717;
wire n_16606;
wire n_39417;
wire n_34089;
wire n_39560;
wire n_33525;
wire n_24736;
wire n_7425;
wire n_47213;
wire n_31332;
wire n_42925;
wire FE_OCP_RBN2168_n_32892;
wire n_9074;
wire FE_OCP_RBN1691_n_19052;
wire n_11456;
wire n_31226;
wire n_12612;
wire n_27287;
wire n_38412;
wire n_18755;
wire n_12463;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_6_;
wire n_39519;
wire n_11718;
wire n_28341;
wire newNet_2076;
wire n_7584;
wire n_22037;
wire n_4812;
wire FE_RN_993_0;
wire n_43852;
wire n_20178;
wire n_14219;
wire n_47249;
wire n_5112;
wire newNet_3438;
wire FE_RN_1745_0;
wire n_21261;
wire n_1226;
wire n_36190;
wire n_1113;
wire n_10512;
wire n_30689;
wire n_31648;
wire n_39633;
wire n_29562;
wire n_2641;
wire n_41642;
wire n_36118;
wire n_40426;
wire n_33887;
wire n_3597;
wire delay_xor_ln21_unr6_stage3_stallmux_q_10_;
wire n_35364;
wire n_24354;
wire n_29875;
wire n_1480;
wire FE_RN_893_0;
wire n_926;
wire n_18037;
wire n_41729;
wire n_31132;
wire n_29620;
wire newNet_2313;
wire n_6394;
wire n_32156;
wire n_9827;
wire n_36913;
wire n_46165;
wire n_29632;
wire n_3270;
wire n_10522;
wire n_14720;
wire newNet_665;
wire n_13122;
wire n_8755;
wire n_4895;
wire n_3835;
wire n_41670;
wire n_7225;
wire n_24217;
wire newNet_525;
wire n_4059;
wire n_35476;
wire n_9630;
wire FE_RN_1592_0;
wire n_31821;
wire n_32443;
wire FE_OCP_RBN2395_n_8288;
wire n_26877;
wire n_29478;
wire n_8971;
wire n_35807;
wire n_34154;
wire n_35852;
wire n_16351;
wire n_43547;
wire n_41280;
wire n_12965;
wire n_34338;
wire n_2604;
wire n_43035;
wire n_44054;
wire n_37174;
wire n_31857;
wire n_15851;
wire n_38519;
wire n_11301;
wire newNet_2142;
wire n_14510;
wire n_10880;
wire FE_OCP_RBN3522_n_8242;
wire n_44875;
wire n_32939;
wire n_1957;
wire n_36943;
wire n_28138;
wire n_26683;
wire FE_OCP_RBN2655_n_9198;
wire n_30213;
wire n_33468;
wire n_19613;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_25_;
wire n_41612;
wire n_14388;
wire newNet_98;
wire n_36398;
wire n_29694;
wire newNet_206;
wire n_12441;
wire FE_RN_1686_0;
wire n_28293;
wire n_40271;
wire newNet_3316;
wire n_23658;
wire n_26583;
wire n_12123;
wire n_19778;
wire n_20074;
wire n_39216;
wire n_27788;
wire n_23606;
wire n_23641;
wire n_29824;
wire n_41053;
wire FE_OCP_RBN3729_n_43230;
wire FE_RN_1148_0;
wire newNet_2041;
wire n_3728;
wire n_26610;
wire n_30127;
wire n_17337;
wire n_37074;
wire n_3916;
wire n_27315;
wire n_31268;
wire n_2544;
wire n_29449;
wire n_26302;
wire n_34650;
wire n_7880;
wire newNet_405;
wire n_23954;
wire n_5949;
wire n_33622;
wire n_10648;
wire n_37407;
wire n_37547;
wire n_29752;
wire n_21118;
wire n_23992;
wire n_22892;
wire n_28699;
wire n_16423;
wire FE_OCP_RBN2105_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_22393;
wire FE_OCP_RBN2524_n_8951;
wire n_26084;
wire n_20635;
wire newNet_3720;
wire n_19378;
wire newNet_576;
wire n_43560;
wire n_39449;
wire n_16400;
wire n_13982;
wire n_34637;
wire newNet_3616;
wire n_32087;
wire n_4940;
wire n_12797;
wire n_40064;
wire n_12763;
wire newNet_3497;
wire newNet_3026;
wire n_1888;
wire n_36580;
wire n_12131;
wire n_3429;
wire n_37628;
wire FE_RN_915_0;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_13_;
wire n_26712;
wire n_9941;
wire n_16628;
wire n_24555;
wire n_40744;
wire n_37805;
wire FE_OCPN1387_n_11041;
wire newNet_1011;
wire n_39042;
wire n_4952;
wire n_8771;
wire n_6826;
wire n_2718;
wire FE_OCP_DRV_N1607_n_31473;
wire FE_OCP_RBN1357_n_30298;
wire n_30275;
wire n_24009;
wire n_2186;
wire n_27580;
wire n_26134;
wire newNet_2573;
wire n_36895;
wire n_30930;
wire n_16285;
wire n_21890;
wire newNet_284;
wire n_26413;
wire n_47179;
wire newNet_1072;
wire n_39312;
wire n_11709;
wire n_34668;
wire n_1068;
wire n_31435;
wire n_23803;
wire n_11647;
wire n_12234;
wire n_23814;
wire n_9522;
wire n_39343;
wire n_11878;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_19_;
wire n_625;
wire n_22358;
wire n_10486;
wire n_30408;
wire n_1751;
wire n_33501;
wire n_39163;
wire n_35617;
wire n_26326;
wire newNet_1902;
wire n_41208;
wire newNet_827;
wire n_1864;
wire n_18625;
wire n_21219;
wire n_16541;
wire n_32601;
wire n_41150;
wire n_43617;
wire n_34040;
wire n_44490;
wire n_14240;
wire n_7101;
wire FE_OCP_RBN2721_n_9494;
wire n_2761;
wire n_1159;
wire n_16668;
wire delay_xor_ln21_unr9_stage4_stallmux_q_15_;
wire n_36658;
wire n_14052;
wire n_31619;
wire newNet_918;
wire newNet_1505;
wire n_1716;
wire delay_xor_ln22_unr6_stage3_stallmux_q_13_;
wire n_13693;
wire n_18831;
wire n_24861;
wire n_23116;
wire n_13626;
wire FE_OFN734_n_22641;
wire newNet_2631;
wire n_14999;
wire n_33079;
wire n_28191;
wire n_47000;
wire n_28154;
wire n_35043;
wire n_31846;
wire n_37618;
wire n_36009;
wire n_45072;
wire n_8603;
wire newNet_1994;
wire n_17994;
wire n_36317;
wire n_9913;
wire n_10169;
wire n_28008;
wire n_19965;
wire n_35996;
wire n_31466;
wire n_36556;
wire n_14461;
wire n_26895;
wire n_30750;
wire n_3755;
wire n_28845;
wire newNet_2716;
wire FE_RN_1024_0;
wire n_31036;
wire n_3518;
wire n_38570;
wire delay_add_ln22_unr23_stage9_stallmux_q_27_;
wire n_11366;
wire n_30833;
wire newNet_783;
wire FE_OCP_RBN2140_FE_OCPN861_n_45450;
wire n_13781;
wire FE_OCPN1733_n_16143;
wire n_784;
wire delay_xor_ln21_unr6_stage3_stallmux_q_18_;
wire n_3321;
wire n_7766;
wire n_9918;
wire n_26210;
wire n_43228;
wire FE_RN_246_0;
wire n_1471;
wire n_41519;
wire n_15486;
wire n_35111;
wire n_41754;
wire n_14871;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_22_;
wire n_19700;
wire newNet_3177;
wire n_6281;
wire n_10478;
wire n_19890;
wire FE_OCP_RBN2334_n_24359;
wire FE_OCPN894_n_6521;
wire n_6643;
wire n_42945;
wire n_47267;
wire n_18133;
wire n_5096;
wire FE_RN_853_0;
wire n_16110;
wire n_35109;
wire n_20670;
wire FE_OCP_RBN2902_n_44174;
wire n_2254;
wire n_27750;
wire n_29847;
wire n_37246;
wire n_29398;
wire n_12144;
wire newNet_1831;
wire n_4646;
wire newNet_83;
wire n_20182;
wire n_7674;
wire n_22022;
wire n_22920;
wire newNet_623;
wire n_30248;
wire n_20646;
wire n_19549;
wire n_40205;
wire n_35468;
wire n_6342;
wire n_326;
wire FE_OCP_RBN2905_n_16197;
wire n_4902;
wire FE_OCP_RBN2434_n_14072;
wire FE_OCP_RBN2505_n_13896;
wire newNet_774;
wire FE_RN_439_0;
wire n_8385;
wire n_32704;
wire FE_RN_1273_0;
wire n_38515;
wire n_22761;
wire n_34403;
wire n_6388;
wire n_20481;
wire n_25764;
wire n_45318;
wire n_21288;
wire n_45760;
wire n_5638;
wire n_6310;
wire n_41016;
wire n_10282;
wire delay_sub_ln23_0_unr30_stage10_stallmux_q;
wire n_8929;
wire n_2492;
wire n_42267;
wire n_31997;
wire n_3280;
wire n_42468;
wire n_18679;
wire n_40354;
wire n_19000;
wire newNet_237;
wire newNet_1910;
wire FE_OCPN1261_n_20242;
wire n_1130;
wire n_43606;
wire n_35954;
wire newNet_369;
wire n_28363;
wire newNet_894;
wire n_5256;
wire delay_add_ln22_unr27_stage10_stallmux_q_8_;
wire newNet_817;
wire n_5157;
wire n_9137;
wire n_32483;
wire n_11114;
wire n_23761;
wire n_42043;
wire newNet_761;
wire n_31136;
wire newNet_244;
wire n_6320;
wire FE_RN_487_0;
wire n_32388;
wire n_25383;
wire n_19542;
wire n_32887;
wire n_38703;
wire newNet_660;
wire n_20594;
wire n_9681;
wire n_19945;
wire newNet_757;
wire n_40071;
wire newNet_873;
wire n_34116;
wire FE_OFN817_n_2285;
wire n_40983;
wire n_18796;
wire newNet_1878;
wire n_36033;
wire newNet_821;
wire n_8686;
wire n_39701;
wire n_25957;
wire n_12622;
wire newNet_2775;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_8_;
wire n_8453;
wire n_42136;
wire n_29497;
wire n_30220;
wire n_31956;
wire n_42692;
wire n_15948;
wire n_9198;
wire n_26373;
wire n_17409;
wire FE_OCPN942_n_44925;
wire n_9151;
wire n_29073;
wire n_6263;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_5_;
wire FE_OFN836_n_4575;
wire n_22267;
wire n_36747;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_13_;
wire n_25618;
wire FE_RN_301_0;
wire n_39529;
wire n_46213;
wire n_17618;
wire n_14281;
wire n_18335;
wire n_6670;
wire n_25336;
wire n_5773;
wire newNet_1737;
wire n_24080;
wire n_41342;
wire n_26963;
wire n_19516;
wire n_8240;
wire FE_OCP_RBN2455_n_14157;
wire n_41084;
wire newNet_3440;
wire n_25854;
wire FE_OCP_RBN1183_n_14638;
wire FE_OCP_RBN2701_n_4041;
wire n_1939;
wire n_4139;
wire n_14072;
wire n_19633;
wire n_7355;
wire n_40134;
wire n_29472;
wire n_5998;
wire n_15752;
wire n_18501;
wire n_15230;
wire n_1214;
wire n_21073;
wire n_11324;
wire n_39581;
wire n_4746;
wire n_5495;
wire n_42454;
wire n_11634;
wire n_28532;
wire n_39859;
wire n_18290;
wire n_11398;
wire n_104;
wire n_19382;
wire n_33236;
wire n_18876;
wire newNet_2172;
wire n_42506;
wire n_6554;
wire n_24957;
wire n_23119;
wire FE_RN_1256_0;
wire n_33304;
wire n_22954;
wire n_7810;
wire n_39228;
wire n_43367;
wire newNet_3658;
wire n_9936;
wire delay_xor_ln22_unr18_stage7_stallmux_q_13_;
wire n_42763;
wire n_14764;
wire n_4936;
wire n_11749;
wire n_16747;
wire n_25312;
wire n_29925;
wire delay_xor_ln22_unr3_stage2_stallmux_q_26_;
wire n_32415;
wire n_23464;
wire n_28044;
wire n_4576;
wire n_7671;
wire n_32438;
wire n_7046;
wire n_32352;
wire n_34544;
wire newNet_376;
wire FE_RN_91_0;
wire n_11972;
wire n_14185;
wire delay_xor_ln22_unr21_stage8_stallmux_q_4_;
wire n_6235;
wire FE_OCP_RBN2421_n_24505;
wire n_24412;
wire n_21114;
wire n_32967;
wire n_22941;
wire n_914;
wire FE_RN_1261_0;
wire n_38508;
wire n_1660;
wire n_7990;
wire n_38745;
wire n_33956;
wire FE_OCP_RBN3068_n_43230;
wire n_15452;
wire n_10565;
wire n_10590;
wire n_57;
wire n_43454;
wire n_34975;
wire n_13558;
wire n_21280;
wire n_39061;
wire n_28062;
wire n_11787;
wire n_639;
wire FE_OCP_RBN2369_n_38545;
wire n_34810;
wire n_4177;
wire FE_OFN627_n_34445;
wire n_37573;
wire n_10634;
wire n_13166;
wire newNet_2682;
wire n_2328;
wire newNet_1603;
wire n_47332;
wire FE_RN_365_0;
wire FE_RN_341_0;
wire n_1688;
wire n_28605;
wire n_37104;
wire n_40814;
wire n_11583;
wire FE_OCP_RBN2716_n_14982;
wire n_40196;
wire n_14547;
wire n_41985;
wire n_24867;
wire n_11022;
wire FE_OCP_DRV_N1584_n_30917;
wire n_765;
wire newNet_2742;
wire n_31884;
wire n_5701;
wire n_10267;
wire n_39453;
wire newNet_1346;
wire n_5145;
wire n_43917;
wire n_11509;
wire n_28424;
wire n_27141;
wire n_7660;
wire n_348;
wire n_2709;
wire n_3558;
wire n_2892;
wire n_8174;
wire n_39006;
wire n_12192;
wire n_31568;
wire FE_OCP_RBN2398_n_38586;
wire newNet_1216;
wire n_37441;
wire n_39086;
wire n_1246;
wire newNet_1367;
wire n_11210;
wire newNet_2388;
wire n_32562;
wire n_28480;
wire n_20721;
wire newNet_2420;
wire FE_OCPN848_n_3597;
wire n_19025;
wire n_17705;
wire n_36699;
wire newNet_1549;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_28_;
wire n_39270;
wire n_4198;
wire newNet_1089;
wire n_17924;
wire n_1902;
wire n_41602;
wire n_14732;
wire n_18049;
wire n_29263;
wire n_19609;
wire n_7599;
wire n_8099;
wire n_8769;
wire n_3542;
wire n_33964;
wire n_10776;
wire FE_RN_1005_0;
wire n_5813;
wire newNet_1979;
wire n_31431;
wire n_36056;
wire n_34097;
wire n_3659;
wire n_12538;
wire n_42725;
wire n_21950;
wire n_41248;
wire n_36510;
wire n_25304;
wire n_24617;
wire n_14835;
wire newNet_1126;
wire FE_OCPN1744_n_24962;
wire n_10711;
wire n_24770;
wire n_31806;
wire n_45209;
wire newNet_2738;
wire n_38285;
wire n_37181;
wire FE_OCP_RBN2145_FE_OCPN861_n_45450;
wire n_1019;
wire n_22244;
wire n_20570;
wire newNet_3750;
wire n_36135;
wire n_7275;
wire n_38394;
wire n_17415;
wire n_32393;
wire FE_OCP_RBN3443_n_37945;
wire n_3819;
wire n_898;
wire n_2230;
wire n_29916;
wire n_30154;
wire n_120;
wire n_1367;
wire n_30296;
wire n_24842;
wire n_17433;
wire n_9186;
wire n_20031;
wire newNet_1120;
wire n_5774;
wire n_27535;
wire n_13584;
wire n_10910;
wire n_4458;
wire n_32733;
wire n_25378;
wire n_17554;
wire n_9350;
wire n_25136;
wire n_28051;
wire n_16172;
wire n_40511;
wire n_25912;
wire n_33289;
wire n_17399;
wire FE_RN_916_0;
wire n_31344;
wire n_5011;
wire n_16338;
wire n_38186;
wire n_25477;
wire n_13456;
wire n_40847;
wire n_35119;
wire n_34327;
wire n_33217;
wire n_26189;
wire n_15891;
wire n_24055;
wire n_25735;
wire newNet_1769;
wire FE_OCP_RBN2830_n_10198;
wire newNet_3219;
wire FE_RN_855_0;
wire n_17772;
wire n_8736;
wire n_23304;
wire n_13855;
wire n_2088;
wire n_42330;
wire n_8875;
wire n_20304;
wire delay_add_ln22_unr2_stage2_stallmux_q_2_;
wire n_32238;
wire n_16369;
wire n_5482;
wire n_39132;
wire n_9102;
wire n_30944;
wire n_23874;
wire n_18016;
wire delay_add_ln22_unr20_stage8_stallmux_q_24_;
wire n_24347;
wire n_16637;
wire n_23527;
wire n_10010;
wire n_3184;
wire newNet_428;
wire n_12562;
wire newNet_2661;
wire newNet_886;
wire n_16053;
wire n_42818;
wire n_28683;
wire n_793;
wire n_33673;
wire newNet_1045;
wire n_29613;
wire n_17093;
wire newNet_2557;
wire n_28529;
wire n_9255;
wire n_43158;
wire n_15290;
wire FE_OCP_RBN1134_n_16041;
wire n_19803;
wire n_20020;
wire FE_OCP_RBN2325_n_13616;
wire n_6037;
wire n_42896;
wire n_28449;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_26_;
wire n_42005;
wire n_13783;
wire n_6161;
wire n_5921;
wire n_39790;
wire n_6913;
wire n_13411;
wire n_6329;
wire n_35207;
wire n_1852;
wire n_38863;
wire n_26020;
wire FE_RN_197_0;
wire n_2151;
wire n_25040;
wire n_7287;
wire n_25228;
wire FE_OFN0_n_43918;
wire n_41845;
wire n_5958;
wire FE_OCPN1768_n_29715;
wire newNet_2353;
wire n_5196;
wire newNet_2599;
wire newNet_709;
wire FE_OCP_RBN2456_n_13765;
wire n_33725;
wire n_13770;
wire FE_RN_450_0;
wire delay_xor_ln22_unr15_stage6_stallmux_q_4_;
wire n_23900;
wire n_20865;
wire FE_RN_1493_0;
wire n_45903;
wire FE_RN_616_0;
wire n_37835;
wire FE_RN_1500_0;
wire newNet_1404;
wire n_5719;
wire FE_OCP_RBN3001_n_42959;
wire delay_add_ln22_unr14_stage6_stallmux_q_28_;
wire n_13828;
wire n_8561;
wire n_11544;
wire n_18416;
wire n_6223;
wire n_16954;
wire n_19786;
wire n_16302;
wire n_15305;
wire n_1703;
wire n_39359;
wire n_9730;
wire newNet_1428;
wire n_2575;
wire n_23428;
wire n_22668;
wire n_27527;
wire n_7977;
wire n_18696;
wire newNet_2974;
wire n_26453;
wire n_17466;
wire n_8065;
wire n_25568;
wire FE_RN_913_0;
wire n_40051;
wire n_43473;
wire n_16102;
wire FE_OCP_RBN2128_n_6745;
wire n_3563;
wire n_36091;
wire newNet_2032;
wire n_19107;
wire FE_RN_1706_0;
wire n_37562;
wire n_23169;
wire n_7029;
wire n_11766;
wire newNet_2291;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_19_;
wire n_26770;
wire FE_OCP_RBN2135_n_11780;
wire FE_OCP_RBN2329_n_9003;
wire FE_RN_1118_0;
wire n_18456;
wire n_6398;
wire n_8831;
wire n_17136;
wire n_7221;
wire n_28474;
wire n_47253;
wire n_41099;
wire n_21446;
wire n_7853;
wire n_27962;
wire n_13240;
wire n_4368;
wire FE_RN_172_0;
wire n_30579;
wire FE_RN_1428_0;
wire n_32934;
wire n_8273;
wire n_23980;
wire n_21714;
wire n_40164;
wire FE_OCP_RBN2982_n_26767;
wire newNet_3326;
wire n_10790;
wire n_12177;
wire n_29195;
wire n_9118;
wire FE_OCP_RBN3846_FE_RN_1242_0;
wire n_24403;
wire n_21868;
wire n_33591;
wire n_45820;
wire n_26795;
wire FE_OCP_RBN3845_FE_RN_1242_0;
wire n_38686;
wire n_2353;
wire n_21238;
wire n_13892;
wire n_32241;
wire n_1763;
wire n_32694;
wire n_41616;
wire n_7267;
wire n_17679;
wire newNet_2721;
wire n_2017;
wire n_33004;
wire n_45489;
wire n_20600;
wire n_33583;
wire newNet_3551;
wire n_1332;
wire n_32182;
wire n_32451;
wire n_14456;
wire newNet_1180;
wire n_5735;
wire n_31249;
wire FE_RN_1327_0;
wire n_12137;
wire n_29882;
wire n_35659;
wire n_30593;
wire n_42054;
wire n_16572;
wire n_15580;
wire n_41360;
wire n_21095;
wire FE_RN_636_0;
wire n_35635;
wire n_42012;
wire newNet_3587;
wire n_25365;
wire n_28329;
wire n_16508;
wire n_46159;
wire n_25268;
wire FE_OFN802_n_46285;
wire FE_OCP_RBN2742_n_15206;
wire FE_OCP_RBN2763_n_25732;
wire n_4676;
wire FE_OCP_RBN3375_n_6822;
wire n_23701;
wire n_10085;
wire n_23908;
wire n_30548;
wire n_10137;
wire FE_OCP_RBN3117_n_22710;
wire n_2845;
wire n_42159;
wire n_35710;
wire n_32404;
wire FE_OCP_RBN2529_n_9044;
wire n_18386;
wire n_5440;
wire n_41266;
wire n_35173;
wire n_10696;
wire n_22617;
wire n_26466;
wire FE_OCP_RBN2801_n_15706;
wire n_2198;
wire n_28638;
wire n_11651;
wire FE_OCP_RBN2206_n_12907;
wire n_29296;
wire n_26181;
wire n_6352;
wire n_20713;
wire n_8416;
wire n_600;
wire FE_RN_1777_0;
wire n_10059;
wire n_33421;
wire n_31262;
wire n_20786;
wire FE_OCPN941_n_44925;
wire n_26607;
wire n_12649;
wire n_40659;
wire n_6687;
wire n_23516;
wire n_37468;
wire n_2983;
wire n_12892;
wire n_2446;
wire n_7202;
wire n_137;
wire n_37792;
wire n_31209;
wire n_37000;
wire n_16495;
wire newNet_2766;
wire delay_add_ln22_unr27_stage10_stallmux_q_5_;
wire n_10670;
wire newNet_2797;
wire n_29628;
wire n_20685;
wire n_13290;
wire n_32458;
wire FE_OCP_RBN2564_FE_RN_1125_0;
wire n_19863;
wire n_8195;
wire n_32446;
wire n_20336;
wire n_8696;
wire n_13360;
wire FE_RN_1375_0;
wire n_5677;
wire n_22882;
wire n_26196;
wire n_33350;
wire n_12793;
wire n_331;
wire n_2938;
wire n_32508;
wire n_23822;
wire newNet_2139;
wire n_9649;
wire delay_add_ln22_unr11_stage5_stallmux_q_1_;
wire n_25867;
wire n_20369;
wire n_36655;
wire n_1839;
wire n_40219;
wire n_32172;
wire n_46222;
wire n_15377;
wire n_23700;
wire newNet_2371;
wire n_23492;
wire newNet_2497;
wire n_40367;
wire n_34076;
wire n_2820;
wire n_31830;
wire n_1833;
wire n_40565;
wire newNet_1662;
wire FE_RN_379_0;
wire n_46186;
wire n_29572;
wire FE_OCP_RBN1336_n_20941;
wire n_40186;
wire newNet_604;
wire n_2535;
wire n_44809;
wire n_35421;
wire FE_OCP_RBN1695_n_19206;
wire n_29819;
wire n_1915;
wire newNet_214;
wire n_18022;
wire n_17913;
wire n_21012;
wire n_4997;
wire n_9775;
wire FE_RN_373_0;
wire n_22544;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_5_;
wire n_9148;
wire n_43375;
wire n_41641;
wire n_4802;
wire n_17015;
wire n_37225;
wire n_31143;
wire n_14973;
wire n_30417;
wire n_4355;
wire n_36561;
wire n_11867;
wire n_39934;
wire n_25641;
wire n_38990;
wire n_6638;
wire n_17658;
wire n_21900;
wire n_10554;
wire n_8525;
wire n_29636;
wire n_3992;
wire n_39118;
wire n_22971;
wire n_9480;
wire FE_RN_851_0;
wire n_15245;
wire n_29560;
wire newNet_3536;
wire newNet_572;
wire FE_OCP_RBN2628_n_14590;
wire n_31124;
wire n_26787;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_25_;
wire n_28758;
wire n_28358;
wire n_22411;
wire newNet_234;
wire newNet_3664;
wire n_42238;
wire n_190;
wire n_32954;
wire n_6294;
wire n_12254;
wire n_26731;
wire n_25094;
wire n_15607;
wire n_25645;
wire n_40736;
wire n_7572;
wire n_12707;
wire n_37423;
wire FE_RN_1042_0;
wire newNet_2191;
wire delay_add_ln22_unr23_stage9_stallmux_q_14_;
wire n_28624;
wire n_20834;
wire n_19144;
wire FE_OCPN1476_n_23708;
wire newNet_522;
wire n_36532;
wire n_29593;
wire n_41501;
wire n_6276;
wire n_21579;
wire n_2027;
wire FE_OCPN946_n_1780;
wire n_20760;
wire newNet_2534;
wire n_10842;
wire n_21082;
wire n_22119;
wire newNet_2067;
wire n_33879;
wire n_19408;
wire n_36681;
wire n_25323;
wire n_22787;
wire newNet_1256;
wire n_41322;
wire n_10182;
wire n_33922;
wire n_8237;
wire n_34817;
wire n_4106;
wire newNet_742;
wire n_4868;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_14_;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_22_;
wire n_36379;
wire n_30712;
wire delay_xor_ln22_unr18_stage7_stallmux_q_7_;
wire n_40862;
wire n_25994;
wire n_20826;
wire newNet_2204;
wire n_14067;
wire n_38269;
wire n_19924;
wire n_37377;
wire n_43189;
wire n_3576;
wire FE_RN_1631_0;
wire n_41359;
wire FE_OCPN3166_n_44267;
wire FE_OCP_RBN2949_n_10852;
wire n_20526;
wire newNet_545;
wire FE_RN_398_0;
wire newNet_330;
wire n_7381;
wire FE_OCP_RBN2632_n_30170;
wire n_9824;
wire n_24965;
wire n_30114;
wire n_21371;
wire newNet_3321;
wire n_47181;
wire FE_OCP_RBN2626_n_3848;
wire n_40541;
wire n_9295;
wire n_31875;
wire n_16530;
wire n_5576;
wire n_28798;
wire n_2061;
wire n_33529;
wire n_23282;
wire FE_OCP_RBN2636_n_38806;
wire FE_RN_1294_0;
wire FE_OFN765_n_15670;
wire n_16123;
wire n_19428;
wire n_4939;
wire n_32464;
wire n_35984;
wire newNet_2826;
wire n_8967;
wire n_40302;
wire n_1614;
wire n_5935;
wire n_38736;
wire n_15599;
wire n_41170;
wire n_28737;
wire n_20119;
wire n_23505;
wire n_27602;
wire newNet_3259;
wire n_1002;
wire newNet_1281;
wire n_39445;
wire n_4558;
wire n_22826;
wire n_40476;
wire n_40266;
wire n_40885;
wire n_28289;
wire n_22357;
wire newNet_2867;
wire n_6592;
wire n_4063;
wire n_18981;
wire n_26972;
wire newNet_643;
wire n_39537;
wire FE_OFN780_n_17093;
wire n_15551;
wire n_17847;
wire newNet_1105;
wire n_41666;
wire n_6697;
wire n_32106;
wire n_22939;
wire n_31643;
wire n_21438;
wire n_19912;
wire newNet_3084;
wire n_4149;
wire n_7305;
wire n_10022;
wire n_27922;
wire n_40619;
wire n_25054;
wire n_21318;
wire n_17509;
wire n_17579;
wire n_13177;
wire FE_RN_1219_0;
wire n_43353;
wire n_38796;
wire n_33027;
wire n_46356;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_18_;
wire n_2267;
wire n_34955;
wire n_38003;
wire n_1802;
wire FE_RN_1044_0;
wire FE_OCP_RBN2270_n_13489;
wire n_41018;
wire n_15768;
wire n_21797;
wire n_12827;
wire n_1520;
wire n_39496;
wire n_27340;
wire newNet_3697;
wire n_1078;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_10_;
wire n_36802;
wire n_5594;
wire n_10688;
wire n_33558;
wire FE_OCP_RBN2809_n_35285;
wire n_31420;
wire FE_OCP_DRV_N1595_n_21458;
wire n_39952;
wire newNet_3208;
wire n_27569;
wire n_36881;
wire n_16321;
wire n_4594;
wire n_12516;
wire n_31959;
wire n_17054;
wire n_34528;
wire n_28164;
wire n_34384;
wire n_29868;
wire n_12596;
wire n_2698;
wire n_26914;
wire n_25885;
wire n_38818;
wire FE_RN_380_0;
wire n_18091;
wire newNet_3356;
wire n_333;
wire n_27693;
wire n_39320;
wire n_35191;
wire n_23332;
wire n_36410;
wire newNet_22;
wire n_1737;
wire n_39301;
wire n_33618;
wire newNet_1204;
wire FE_RN_358_0;
wire n_24296;
wire n_28928;
wire n_37046;
wire FE_OCP_RBN3839_n_19513;
wire n_15840;
wire n_37455;
wire n_37543;
wire n_45898;
wire n_31429;
wire n_16071;
wire n_8281;
wire n_40962;
wire n_4898;
wire n_39467;
wire n_34244;
wire n_20073;
wire n_18853;
wire n_36191;
wire n_36140;
wire n_12638;
wire newNet_3548;
wire newNet_976;
wire n_14460;
wire n_43909;
wire n_22673;
wire n_43240;
wire n_36765;
wire newNet_455;
wire n_31151;
wire n_46988;
wire n_41445;
wire n_3837;
wire newNet_1989;
wire n_23808;
wire n_16745;
wire n_21622;
wire n_32728;
wire n_28347;
wire n_20538;
wire FE_OCP_RBN2256_n_37844;
wire n_38890;
wire n_24909;
wire n_40711;
wire FE_RN_1585_0;
wire n_23923;
wire n_21166;
wire n_36402;
wire n_27349;
wire n_2860;
wire n_28651;
wire n_18616;
wire n_12333;
wire n_27490;
wire n_41435;
wire n_14041;
wire n_41876;
wire n_8068;
wire n_35570;
wire newNet_2289;
wire newNet_1589;
wire n_13683;
wire n_5473;
wire n_22065;
wire n_28109;
wire n_17255;
wire n_35889;
wire n_14868;
wire n_1343;
wire n_17820;
wire n_20321;
wire n_9573;
wire n_21721;
wire FE_RN_1618_0;
wire n_39986;
wire n_33454;
wire FE_RN_1783_0;
wire n_37230;
wire n_24603;
wire n_36144;
wire n_36046;
wire n_33126;
wire n_4297;
wire n_22914;
wire FE_OCP_RBN3539_n_3335;
wire n_30637;
wire n_14642;
wire n_44818;
wire n_47019;
wire n_8742;
wire n_34771;
wire n_13765;
wire n_5895;
wire n_10998;
wire n_1873;
wire n_41271;
wire n_27164;
wire newNet_1007;
wire n_358;
wire n_16712;
wire n_1984;
wire n_17533;
wire n_3024;
wire n_31440;
wire n_21909;
wire n_28901;
wire n_7913;
wire n_36303;
wire n_3765;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_17_;
wire n_43297;
wire n_12678;
wire n_20280;
wire n_14895;
wire n_8723;
wire n_43325;
wire n_21853;
wire n_22595;
wire n_13888;
wire n_16391;
wire delay_xor_ln21_unr6_stage3_stallmux_q_7_;
wire newNet_327;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_10_;
wire n_32803;
wire n_2896;
wire n_12550;
wire FE_RN_1246_0;
wire n_6578;
wire n_15250;
wire delay_add_ln22_unr8_stage4_stallmux_q_31_;
wire n_1960;
wire n_43028;
wire n_20262;
wire n_43330;
wire n_43638;
wire n_27033;
wire FE_OCP_RBN2853_n_26169;
wire n_14883;
wire n_9129;
wire newNet_677;
wire n_30758;
wire n_1969;
wire n_4683;
wire n_26628;
wire n_32554;
wire n_7129;
wire n_13367;
wire n_3137;
wire n_40588;
wire n_17186;
wire n_36615;
wire n_23098;
wire n_11737;
wire n_31403;
wire n_11263;
wire n_37752;
wire n_21121;
wire n_35945;
wire newNet_2359;
wire FE_OCPN3753_n_1448;
wire n_22818;
wire n_42900;
wire n_25711;
wire n_11335;
wire n_22620;
wire n_42595;
wire newNet_2153;
wire n_11388;
wire n_35189;
wire n_38190;
wire n_23034;
wire n_4009;
wire n_14250;
wire n_21726;
wire n_3928;
wire n_4736;
wire n_38482;
wire n_38055;
wire newNet_3241;
wire n_10165;
wire FE_RN_824_0;
wire n_5059;
wire n_2589;
wire newNet_1196;
wire n_15926;
wire n_4128;
wire newNet_3214;
wire n_24910;
wire n_30941;
wire n_40798;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_26_;
wire n_40453;
wire n_6723;
wire newNet_1390;
wire FE_RN_1354_0;
wire n_15514;
wire n_19035;
wire n_42191;
wire n_28782;
wire n_689;
wire n_33072;
wire n_23212;
wire n_41169;
wire newNet_1410;
wire n_27224;
wire n_46951;
wire n_16146;
wire n_32838;
wire n_43534;
wire n_43508;
wire n_25156;
wire n_44811;
wire n_42386;
wire n_569;
wire n_35099;
wire n_44221;
wire n_29125;
wire n_39179;
wire newNet_863;
wire FE_OCP_RBN3283_n_44365;
wire FE_OCP_DRV_N1560_n_34288;
wire n_3629;
wire n_9970;
wire newNet_3511;
wire n_1171;
wire n_26809;
wire n_38140;
wire n_11791;
wire newNet_792;
wire n_2103;
wire n_15200;
wire n_24305;
wire newNet_2778;
wire newNet_990;
wire n_24447;
wire n_10877;
wire FE_OCPN1497_n_26360;
wire FE_RN_456_0;
wire n_15408;
wire n_12805;
wire n_7237;
wire n_30092;
wire n_3849;
wire FE_OCP_RBN2536_n_3645;
wire n_12483;
wire newNet_3248;
wire newNet_595;
wire n_21464;
wire n_24626;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_17_;
wire n_21930;
wire n_28316;
wire n_19585;
wire newNet_69;
wire n_41250;
wire n_13386;
wire n_6949;
wire n_24257;
wire newNet_1262;
wire n_35404;
wire newNet_2464;
wire n_3062;
wire n_26860;
wire n_35319;
wire n_4080;
wire n_36645;
wire n_33184;
wire n_15001;
wire FE_OCP_DRV_N1590_n_21343;
wire n_35225;
wire delay_xor_ln21_unr9_stage4_stallmux_q_5_;
wire n_34893;
wire n_12998;
wire FE_RN_1238_0;
wire n_20068;
wire n_15375;
wire FE_RN_1059_0;
wire n_7179;
wire n_38354;
wire n_24664;
wire n_38039;
wire n_19848;
wire n_24472;
wire n_19979;
wire n_45190;
wire n_254;
wire n_4752;
wire n_9020;
wire n_27500;
wire FE_RN_1217_0;
wire FE_OCP_RBN2348_n_13702;
wire newNet_1354;
wire n_12686;
wire n_998;
wire FE_OCP_RBN3372_n_6745;
wire n_43654;
wire n_39489;
wire n_11510;
wire n_21503;
wire n_36660;
wire n_240;
wire n_4281;
wire n_17312;
wire n_38365;
wire n_42677;
wire n_35723;
wire n_14487;
wire n_5310;
wire n_16346;
wire n_24316;
wire newNet_3529;
wire n_37784;
wire n_9061;
wire n_17179;
wire n_15468;
wire n_6600;
wire n_40769;
wire n_36868;
wire n_26317;
wire n_4103;
wire n_12512;
wire n_30339;
wire n_617;
wire n_16968;
wire n_14112;
wire n_3851;
wire newNet_2956;
wire n_10105;
wire n_38952;
wire n_28075;
wire n_20180;
wire n_1590;
wire FE_RN_706_0;
wire n_26050;
wire n_33334;
wire n_17980;
wire n_29411;
wire n_5555;
wire n_32751;
wire n_28216;
wire n_33102;
wire FE_RN_1156_0;
wire n_12085;
wire n_29457;
wire n_39260;
wire n_31670;
wire n_10971;
wire n_18000;
wire n_33359;
wire n_26813;
wire n_28001;
wire n_36073;
wire n_36789;
wire newNet_945;
wire n_23056;
wire n_10054;
wire n_39109;
wire n_24453;
wire n_4990;
wire n_24063;
wire FE_OCP_DRV_N3739_n_29439;
wire n_25883;
wire newNet_3701;
wire n_11027;
wire n_27204;
wire n_26601;
wire n_4842;
wire newNet_1171;
wire n_43006;
wire newNet_3160;
wire n_4621;
wire n_26640;
wire n_23566;
wire n_42980;
wire n_24276;
wire n_493;
wire n_21880;
wire newNet_1512;
wire FE_RN_1847_0;
wire n_19291;
wire n_23747;
wire n_20341;
wire n_12572;
wire n_20805;
wire n_31588;
wire n_15287;
wire n_43118;
wire n_19652;
wire n_7710;
wire n_18202;
wire n_16195;
wire n_37649;
wire n_14330;
wire n_30905;
wire delay_xor_ln21_unr12_stage5_stallmux_q_5_;
wire n_39881;
wire FE_OCP_RBN1162_n_24701;
wire n_43866;
wire n_8938;
wire newNet_2099;
wire n_13592;
wire newNet_3600;
wire n_12786;
wire n_34532;
wire n_20933;
wire n_13445;
wire newNet_1540;
wire n_42270;
wire n_10639;
wire n_39772;
wire n_42694;
wire n_42202;
wire n_11391;
wire n_44211;
wire newNet_1758;
wire n_45622;
wire newNet_318;
wire n_32656;
wire n_28993;
wire newNet_2089;
wire n_8575;
wire n_41932;
wire n_24105;
wire n_39875;
wire newNet_101;
wire n_18438;
wire n_46957;
wire n_32798;
wire FE_RN_1437_0;
wire n_27240;
wire n_45032;
wire n_21701;
wire n_17824;
wire n_2261;
wire n_26120;
wire n_17544;
wire delay_add_ln22_unr17_stage7_stallmux_q_8_;
wire n_15439;
wire n_22814;
wire n_9790;
wire n_30994;
wire n_7782;
wire n_29328;
wire n_1554;
wire n_20958;
wire FE_OCPN845_n_4046;
wire n_7568;
wire FE_OCP_RBN3622_n_15135;
wire n_32686;
wire newNet_1085;
wire n_37445;
wire n_28649;
wire FE_OCP_RBN1341_n_19077;
wire n_23421;
wire n_15209;
wire n_16191;
wire n_32670;
wire n_13714;
wire n_13239;
wire n_37298;
wire newNet_2515;
wire n_24582;
wire n_23927;
wire n_40048;
wire n_41371;
wire n_34259;
wire n_40641;
wire n_21429;
wire n_34303;
wire n_22524;
wire newNet_1223;
wire newNet_618;
wire n_26992;
wire FE_OFN360_n_9391;
wire n_13221;
wire FE_OCP_RBN2963_n_26231;
wire n_19387;
wire newNet_3081;
wire n_16166;
wire newNet_2892;
wire n_12417;
wire n_44696;
wire n_7385;
wire n_36214;
wire n_34564;
wire FE_RN_402_0;
wire n_47337;
wire n_17473;
wire n_6523;
wire FE_OCP_RBN3091_n_11475;
wire n_42846;
wire n_33266;
wire n_4920;
wire n_24362;
wire n_13139;
wire n_29931;
wire n_25375;
wire FE_OCP_RBN3556_n_44575;
wire n_22134;
wire n_15922;
wire n_6156;
wire n_30708;
wire n_39761;
wire FE_RN_453_0;
wire n_42783;
wire n_19696;
wire n_4838;
wire FE_OCPN915_n_7832;
wire n_28496;
wire n_17517;
wire n_33080;
wire n_31913;
wire newNet_116;
wire n_32782;
wire n_26207;
wire n_23793;
wire n_24114;
wire FE_OCP_RBN3579_n_44944;
wire n_4808;
wire n_30278;
wire n_19830;
wire n_31868;
wire n_12475;
wire n_5613;
wire n_20028;
wire n_22196;
wire n_2373;
wire n_38835;
wire n_21115;
wire n_17806;
wire newNet_2706;
wire n_28619;
wire newNet_41;
wire n_23171;
wire n_7819;
wire n_21434;
wire n_21893;
wire n_1454;
wire n_14123;
wire n_38497;
wire n_22585;
wire n_30096;
wire n_42716;
wire n_218;
wire n_46385;
wire n_28868;
wire n_27098;
wire newNet_1053;
wire n_44866;
wire n_25804;
wire newNet_3303;
wire n_24825;
wire n_12466;
wire n_3407;
wire n_3760;
wire n_22368;
wire n_42599;
wire n_20222;
wire n_40516;
wire n_35352;
wire n_5572;
wire n_10511;
wire n_630;
wire n_43162;
wire n_36885;
wire n_21200;
wire FE_OCP_RBN2950_n_21363;
wire n_18870;
wire n_43816;
wire newNet_431;
wire n_4815;
wire newNet_1394;
wire n_27683;
wire newNet_2363;
wire n_25638;
wire n_9974;
wire n_5763;
wire n_6509;
wire n_30261;
wire FE_OCP_RBN3041_n_46337;
wire newNet_1019;
wire n_4779;
wire n_9355;
wire n_25515;
wire n_19493;
wire newNet_3281;
wire n_40725;
wire FE_RN_285_0;
wire n_42701;
wire n_17026;
wire n_26383;
wire n_27219;
wire newNet_2479;
wire newNet_2681;
wire n_6773;
wire newNet_3179;
wire n_17942;
wire n_17195;
wire n_37464;
wire n_2797;
wire n_37397;
wire n_22548;
wire n_20981;
wire n_14929;
wire n_2319;
wire n_13266;
wire n_29406;
wire n_14700;
wire n_1238;
wire newNet_363;
wire FE_RN_1063_0;
wire FE_OCP_RBN2603_n_39126;
wire n_2710;
wire newNet_2239;
wire n_19020;
wire n_13075;
wire newNet_1033;
wire n_10469;
wire n_5752;
wire n_39662;
wire n_20856;
wire n_19356;
wire n_19459;
wire n_32948;
wire n_674;
wire n_30079;
wire n_19183;
wire n_5619;
wire n_40692;
wire n_28842;
wire FE_OCPN3790_n_36069;
wire n_43114;
wire n_33401;
wire newNet_2255;
wire n_28015;
wire n_10496;
wire n_29879;
wire n_27312;
wire n_16540;
wire n_44358;
wire n_18825;
wire newNet_2759;
wire n_1723;
wire n_40317;
wire newNet_3482;
wire n_15239;
wire n_18240;
wire n_29236;
wire n_2520;
wire n_25522;
wire n_31304;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_17_;
wire n_42495;
wire newNet_3235;
wire newNet_2590;
wire newNet_596;
wire n_24788;
wire newNet_1471;
wire n_33385;
wire n_38424;
wire n_35916;
wire n_28644;
wire n_40407;
wire n_769;
wire n_24539;
wire n_16903;
wire n_5627;
wire FE_OCP_RBN2727_n_4219;
wire n_19714;
wire n_5018;
wire n_43582;
wire n_38752;
wire n_20579;
wire n_15144;
wire n_12870;
wire n_7615;
wire n_10242;
wire n_42472;
wire n_37585;
wire newNet_2181;
wire n_39508;
wire n_37886;
wire n_16264;
wire n_37084;
wire n_16551;
wire n_17581;
wire n_23559;
wire n_32578;
wire n_20345;
wire n_35752;
wire n_35557;
wire n_14162;
wire FE_RN_1160_0;
wire n_32257;
wire n_40110;
wire n_13574;
wire n_40875;
wire n_28157;
wire n_36282;
wire n_13898;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_26_;
wire n_39183;
wire n_37053;
wire n_9239;
wire n_19871;
wire n_13418;
wire n_40896;
wire n_40792;
wire n_9157;
wire delay_add_ln22_unr27_stage10_stallmux_q_24_;
wire n_40116;
wire n_42512;
wire newNet_2762;
wire n_4308;
wire n_15578;
wire newNet_1026;
wire n_7624;
wire n_42300;
wire n_25504;
wire n_19502;
wire FE_OCPN1400_n_8670;
wire n_11278;
wire n_42047;
wire n_10888;
wire FE_RN_899_0;
wire n_39832;
wire n_25257;
wire FE_OCP_RBN3801_delay_xor_ln22_unr12_stage5_stallmux_q_1_;
wire n_13757;
wire n_25499;
wire n_15565;
wire n_7489;
wire n_33496;
wire n_11691;
wire n_472;
wire n_5328;
wire n_15933;
wire n_1156;
wire n_1634;
wire n_18010;
wire n_30589;
wire n_7498;
wire n_13825;
wire n_31903;
wire n_39337;
wire n_5723;
wire n_2679;
wire n_34847;
wire n_16201;
wire n_3447;
wire n_12519;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_0_;
wire n_23300;
wire n_5189;
wire n_36659;
wire FE_RN_328_0;
wire n_31432;
wire n_16136;
wire n_40391;
wire newNet_1271;
wire n_26664;
wire n_36267;
wire n_23190;
wire n_36251;
wire newNet_507;
wire n_3114;
wire n_39756;
wire n_14821;
wire n_26779;
wire n_14879;
wire FE_OCP_RBN2363_n_13785;
wire n_38868;
wire n_34643;
wire n_6059;
wire n_29161;
wire n_10068;
wire n_9325;
wire n_35804;
wire n_7409;
wire newNet_3449;
wire n_25010;
wire n_408;
wire n_15297;
wire n_42031;
wire n_16615;
wire n_38876;
wire n_6077;
wire n_25751;
wire n_25127;
wire n_9626;
wire n_22375;
wire n_29273;
wire n_11012;
wire n_5899;
wire newNet_491;
wire n_24112;
wire n_15093;
wire FE_OCP_RBN2218_FE_OCPN950_n_28595;
wire n_15412;
wire n_14861;
wire n_6806;
wire n_38584;
wire n_9892;
wire n_27995;
wire newNet_719;
wire n_44025;
wire n_33547;
wire n_35853;
wire n_34183;
wire n_31049;
wire n_23893;
wire newNet_2017;
wire n_27831;
wire n_10062;
wire n_4142;
wire n_26849;
wire n_39745;
wire n_16216;
wire n_1497;
wire FE_OCPN1475_n_23708;
wire FE_RN_1004_0;
wire n_10600;
wire FE_RN_1159_0;
wire n_32525;
wire n_19292;
wire n_26387;
wire n_18196;
wire n_5248;
wire newNet_3492;
wire n_22435;
wire n_3356;
wire n_6391;
wire n_9702;
wire n_46143;
wire n_16352;
wire n_25355;
wire n_42371;
wire n_37007;
wire n_7512;
wire n_25284;
wire FE_OCP_RBN2548_n_44944;
wire n_39939;
wire n_25683;
wire n_33125;
wire n_26829;
wire FE_OCP_RBN2351_n_38534;
wire n_22924;
wire n_15320;
wire n_3743;
wire n_12673;
wire n_22650;
wire newNet_1305;
wire FE_OCP_RBN2226_n_7531;
wire newNet_2365;
wire n_29423;
wire n_36833;
wire n_6042;
wire n_26704;
wire n_33416;
wire FE_OCP_RBN2724_n_4219;
wire n_24258;
wire n_8134;
wire n_37166;
wire n_1597;
wire FE_OCPN868_n_16086;
wire n_9761;
wire newNet_2197;
wire n_12862;
wire FE_OCP_RBN1203_n_26121;
wire n_13392;
wire n_38578;
wire delay_add_ln22_unr11_stage5_stallmux_q_23_;
wire n_38640;
wire newNet_3637;
wire n_21944;
wire n_38415;
wire n_18301;
wire n_15962;
wire n_12521;
wire n_12583;
wire n_38074;
wire n_45625;
wire n_20141;
wire n_9899;
wire FE_RN_820_0;
wire n_35200;
wire newNet_1353;
wire n_15671;
wire n_31768;
wire n_1817;
wire n_5346;
wire n_40446;
wire n_36576;
wire n_35542;
wire n_8419;
wire n_26349;
wire newNet_1165;
wire newNet_988;
wire n_16640;
wire n_1568;
wire n_2452;
wire n_21055;
wire n_34365;
wire n_17971;
wire n_38161;
wire n_16918;
wire n_14273;
wire n_28082;
wire n_15416;
wire n_15117;
wire n_16700;
wire n_17758;
wire n_36471;
wire n_33472;
wire n_38215;
wire n_46231;
wire n_33685;
wire n_9121;
wire n_19140;
wire n_40423;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_28_;
wire n_12250;
wire n_22883;
wire n_21020;
wire n_38970;
wire n_38395;
wire n_33997;
wire n_37161;
wire n_36669;
wire n_3792;
wire n_46991;
wire n_31503;
wire n_13674;
wire n_40609;
wire n_25369;
wire n_34402;
wire FE_RN_1404_0;
wire n_13331;
wire newNet_1389;
wire n_14032;
wire n_40429;
wire n_41192;
wire n_37314;
wire n_29515;
wire n_10578;
wire n_22214;
wire delay_add_ln22_unr5_stage3_stallmux_q_19_;
wire n_36711;
wire FE_OFN749_n_45003;
wire FE_OCPN871_n_2737;
wire n_24128;
wire newNet_510;
wire n_30809;
wire n_15860;
wire newNet_1192;
wire n_26752;
wire FE_OCP_RBN1988_delay_xor_ln23_unr6_stage3_stallmux_q;
wire n_1092;
wire n_31550;
wire n_3945;
wire n_9786;
wire n_20234;
wire n_7280;
wire n_22036;
wire n_40504;
wire n_35135;
wire n_4093;
wire n_62;
wire n_8364;
wire newNet_3546;
wire n_37334;
wire n_3879;
wire FE_RN_1536_0;
wire n_38324;
wire FE_RN_1077_0;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_3_;
wire n_3207;
wire n_42311;
wire n_24974;
wire n_22045;
wire n_28978;
wire n_27133;
wire n_15207;
wire n_22168;
wire FE_OCPN1517_n_26752;
wire n_36760;
wire newNet_3757;
wire n_34390;
wire FE_OCP_RBN3217_n_19781;
wire n_19764;
wire n_28243;
wire n_6753;
wire n_13637;
wire FE_OCP_RBN1725_FE_RN_422_0;
wire n_40106;
wire n_35270;
wire n_15177;
wire n_31465;
wire n_20790;
wire FE_OCP_RBN3083_n_31819;
wire n_24833;
wire n_12823;
wire n_12943;
wire n_5272;
wire n_22019;
wire FE_RN_471_0;
wire n_32841;
wire n_7777;
wire n_40021;
wire n_37390;
wire n_41965;
wire n_22774;
wire n_8058;
wire n_2801;
wire n_12275;
wire n_8455;
wire FE_RN_948_0;
wire n_2325;
wire n_26173;
wire newNet_340;
wire n_41121;
wire newNet_3045;
wire n_26039;
wire n_38069;
wire n_22272;
wire n_956;
wire n_22396;
wire n_41872;
wire cos_out_7;
wire n_34717;
wire n_37906;
wire FE_OCPN927_n_26231;
wire n_42220;
wire n_37627;
wire newNet_737;
wire FE_RN_1598_0;
wire n_13550;
wire n_42323;
wire n_29701;
wire FE_RN_1068_0;
wire n_41945;
wire n_6338;
wire n_33006;
wire n_6133;
wire n_14156;
wire n_60;
wire n_1656;
wire n_2129;
wire n_41275;
wire n_31948;
wire n_37180;
wire n_8635;
wire delay_xor_ln21_unr12_stage5_stallmux_q_7_;
wire newNet_1094;
wire n_7341;
wire n_34727;
wire newNet_3378;
wire newNet_2566;
wire n_2474;
wire n_40909;
wire n_31383;
wire n_43835;
wire n_45875;
wire n_38293;
wire n_893;
wire n_12231;
wire n_40911;
wire n_41572;
wire n_42723;
wire FE_OCP_RBN2580_n_3734;
wire n_33113;
wire n_9719;
wire cos_out_10;
wire n_1587;
wire n_31234;
wire n_24552;
wire FE_RN_316_0;
wire n_18596;
wire n_46370;
wire n_37943;
wire n_19365;
wire n_26398;
wire n_18547;
wire FE_RN_1860_0;
wire n_13513;
wire n_10154;
wire n_31809;
wire n_41063;
wire FE_RN_716_0;
wire n_26889;
wire n_42102;
wire n_35236;
wire n_3599;
wire n_9695;
wire n_9756;
wire n_35523;
wire n_9275;
wire n_18461;
wire n_4361;
wire n_23263;
wire n_429;
wire n_9362;
wire n_23804;
wire delay_xor_ln22_unr6_stage3_stallmux_q_15_;
wire n_12180;
wire n_12617;
wire n_14799;
wire n_39378;
wire n_29984;
wire n_34990;
wire n_29721;
wire n_4949;
wire cos_out_27;
wire n_36701;
wire n_18521;
wire n_1810;
wire n_9348;
wire n_33444;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_11_;
wire n_41078;
wire n_14029;
wire n_28751;
wire newNet_2611;
wire FE_RN_863_0;
wire n_40607;
wire n_33520;
wire n_30688;
wire newNet_2829;
wire n_33277;
wire n_3075;
wire n_34606;
wire n_19372;
wire n_362;
wire n_47014;
wire n_40061;
wire n_20300;
wire n_341;
wire n_15090;
wire FE_RN_331_0;
wire FE_RN_1784_0;
wire n_17991;
wire n_23950;
wire n_4327;
wire n_43217;
wire n_21604;
wire n_9623;
wire n_22613;
wire n_21148;
wire FE_OFN626_n_34445;
wire newNet_149;
wire n_42154;
wire n_9764;
wire n_31337;
wire n_17411;
wire n_22556;
wire n_41262;
wire n_35287;
wire FE_RN_335_0;
wire n_29205;
wire n_43524;
wire newNet_1038;
wire n_3179;
wire n_25316;
wire n_24263;
wire n_7111;
wire newNet_1817;
wire n_3307;
wire n_9776;
wire newNet_670;
wire n_233;
wire n_6814;
wire n_1154;
wire n_30063;
wire n_6525;
wire n_30355;
wire n_9726;
wire n_38372;
wire newNet_3611;
wire newNet_174;
wire n_31335;
wire newNet_1576;
wire n_2394;
wire n_26369;
wire n_30495;
wire n_43893;
wire n_29976;
wire newNet_917;
wire n_34667;
wire n_22388;
wire n_17572;
wire n_37450;
wire n_42291;
wire n_34663;
wire n_3481;
wire n_34273;
wire n_3199;
wire n_32880;
wire n_15787;
wire n_27396;
wire n_14464;
wire n_22564;
wire newNet_1790;
wire n_15737;
wire n_29360;
wire n_17423;
wire n_14425;
wire n_2869;
wire n_10544;
wire n_38999;
wire n_36423;
wire FE_OCP_RBN2978_n_5555;
wire n_23380;
wire newNet_313;
wire n_29210;
wire FE_RN_1581_0;
wire n_31557;
wire n_3316;
wire delay_add_ln22_unr14_stage6_stallmux_q_16_;
wire n_32419;
wire n_42609;
wire n_9240;
wire n_42445;
wire n_6092;
wire n_7460;
wire n_46171;
wire n_1210;
wire n_31525;
wire n_27715;
wire n_26932;
wire n_208;
wire n_39971;
wire newNet_3644;
wire n_39168;
wire newNet_3355;
wire newNet_3308;
wire n_25721;
wire n_10398;
wire n_13259;
wire n_29807;
wire newNet_654;
wire newNet_2790;
wire n_10428;
wire n_25207;
wire n_14475;
wire newNet_2810;
wire n_3584;
wire n_43019;
wire n_21665;
wire n_8861;
wire n_15072;
wire newNet_2150;
wire n_27464;
wire n_19244;
wire newNet_2342;
wire n_10489;
wire FE_RN_756_0;
wire n_39823;
wire n_9826;
wire newNet_3072;
wire FE_OCP_RBN3574_n_44563;
wire n_18974;
wire n_41029;
wire n_12930;
wire n_22496;
wire FE_RN_94_0;
wire FE_RN_1665_0;
wire n_6959;
wire n_12936;
wire n_881;
wire FE_RN_218_0;
wire n_43857;
wire n_36951;
wire n_42566;
wire n_30840;
wire n_936;
wire n_10452;
wire n_26685;
wire n_5024;
wire n_31629;
wire n_10940;
wire newNet_2130;
wire n_12326;
wire n_5466;
wire n_42521;
wire newNet_2295;
wire n_35602;
wire newNet_3265;
wire n_8608;
wire n_7843;
wire n_31730;
wire n_4351;
wire n_18670;
wire FE_RN_199_0;
wire n_14513;
wire n_5548;
wire n_14526;
wire newNet_398;
wire n_33757;
wire n_2817;
wire FE_OCP_RBN1206_n_16814;
wire n_5006;
wire n_39846;
wire n_13535;
wire n_3971;
wire n_3271;
wire n_8654;
wire newNet_294;
wire n_140;
wire n_40122;
wire n_21693;
wire n_10380;
wire n_10677;
wire FE_OCP_RBN3038_n_47269;
wire n_2442;
wire n_1942;
wire n_5227;
wire n_37237;
wire n_27016;
wire FE_RN_1161_0;
wire newNet_1743;
wire FE_OCP_RBN3672_n_30820;
wire n_31736;
wire FE_RN_1342_0;
wire FE_RN_673_0;
wire FE_OCPN3764_FE_OCP_RBN2222_n_13010;
wire FE_OCP_RBN3043_n_46337;
wire n_26353;
wire FE_RN_299_0;
wire n_8813;
wire n_7206;
wire newNet_1888;
wire FE_OCPN1471_n_13434;
wire n_2277;
wire n_20968;
wire n_28065;
wire n_26239;
wire n_36246;
wire n_25403;
wire n_21679;
wire n_41799;
wire FE_RN_1000_0;
wire FE_RN_1700_0;
wire newNet_3414;
wire n_32455;
wire n_11171;
wire n_21790;
wire n_8430;
wire FE_OCP_RBN2277_n_24173;
wire n_42036;
wire n_13647;
wire n_35433;
wire FE_OCP_RBN3418_n_12739;
wire n_22893;
wire n_18818;
wire n_35930;
wire n_28396;
wire n_17999;
wire FE_OCPN3751_n_44222;
wire n_44717;
wire n_21985;
wire n_17445;
wire n_37523;
wire n_29292;
wire n_5518;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_9_;
wire n_22347;
wire n_26586;
wire n_30292;
wire n_33870;
wire n_38147;
wire n_28738;
wire FE_RN_226_0;
wire n_28607;
wire FE_RN_1838_0;
wire n_34912;
wire FE_RN_1092_0;
wire n_23969;
wire n_39516;
wire n_32718;
wire n_14995;
wire n_8481;
wire n_42263;
wire n_7762;
wire n_34038;
wire n_15198;
wire n_35282;
wire n_18112;
wire n_12509;
wire n_32850;
wire FE_OCP_RBN3593_n_8902;
wire delay_add_ln22_unr11_stage5_stallmux_q_4_;
wire n_34314;
wire n_27667;
wire n_33864;
wire n_244;
wire newNet_2434;
wire n_30146;
wire FE_OCP_RBN2762_n_15200;
wire n_2140;
wire n_19711;
wire n_8141;
wire n_14413;
wire n_5152;
wire n_3750;
wire n_29947;
wire n_29997;
wire n_30644;
wire n_34695;
wire n_4270;
wire n_12645;
wire n_24175;
wire n_33198;
wire n_12247;
wire n_14496;
wire n_24657;
wire n_8606;
wire n_149;
wire n_32442;
wire n_43071;
wire n_32768;
wire n_4523;
wire n_30484;
wire n_1711;
wire n_19856;
wire newNet_1611;
wire n_38390;
wire n_22422;
wire FE_OCP_RBN1704_n_22740;
wire newNet_3073;
wire newNet_1991;
wire n_27889;
wire n_11205;
wire n_3625;
wire n_7552;
wire n_30249;
wire delay_add_ln22_unr27_stage10_stallmux_q_2_;
wire n_41285;
wire n_3300;
wire newNet_3383;
wire n_18130;
wire n_25763;
wire FE_RN_19_0;
wire newNet_697;
wire newNet_59;
wire n_18931;
wire FE_OCP_RBN2782_n_25997;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_11_;
wire n_29372;
wire n_31399;
wire n_17265;
wire n_14385;
wire n_30838;
wire n_19578;
wire FE_OCP_RBN2487_n_3338;
wire n_1890;
wire n_12394;
wire n_43613;
wire n_813;
wire n_25088;
wire n_33259;
wire n_38369;
wire n_34894;
wire n_21382;
wire n_44661;
wire n_26674;
wire n_8038;
wire n_39806;
wire n_19209;
wire n_19084;
wire newNet_191;
wire n_27172;
wire n_8334;
wire n_30319;
wire FE_RN_1002_0;
wire n_25708;
wire n_24609;
wire n_30935;
wire FE_OCP_RBN1152_n_29053;
wire n_13776;
wire n_8202;
wire n_30455;
wire newNet_2964;
wire n_7089;
wire n_27675;
wire n_38501;
wire n_47259;
wire n_23770;
wire n_2976;
wire n_15728;
wire n_14084;
wire FE_OFN818_n_4575;
wire FE_RN_1158_0;
wire FE_RN_733_0;
wire n_6385;
wire n_13257;
wire n_23646;
wire n_42988;
wire n_4503;
wire n_43877;
wire n_39710;
wire n_1645;
wire n_4798;
wire n_1163;
wire n_9845;
wire n_42634;
wire n_24395;
wire n_7747;
wire newNet_3514;
wire n_8671;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_26_;
wire FE_OCP_RBN2852_n_26169;
wire n_29586;
wire n_17046;
wire FE_RN_435_0;
wire n_43670;
wire FE_RN_344_0;
wire newNet_550;
wire n_4037;
wire n_38707;
wire n_15896;
wire n_5413;
wire n_15660;
wire n_37763;
wire n_9178;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_23_;
wire FE_RN_488_0;
wire n_18352;
wire n_41708;
wire FE_OCP_RBN3430_n_13245;
wire n_23868;
wire n_11500;
wire newNet_1801;
wire n_13271;
wire n_25149;
wire n_11594;
wire FE_OCP_RBN2343_FE_OCPN870_n_2737;
wire n_22866;
wire n_30976;
wire n_8429;
wire n_5873;
wire n_39423;
wire n_8782;
wire n_43502;
wire n_43281;
wire n_8255;
wire n_15257;
wire FE_OCPN1018_n_23078;
wire n_42160;
wire n_31952;
wire n_32195;
wire FE_RN_707_0;
wire n_15589;
wire n_27232;
wire n_45508;
wire n_28883;
wire n_23026;
wire newNet_1399;
wire n_25441;
wire n_25782;
wire n_3090;
wire newNet_810;
wire n_33647;
wire n_33841;
wire n_39540;
wire n_37175;
wire newNet_553;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_4_;
wire n_23369;
wire FE_OCPN1224_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire FE_OCP_RBN3507_n_13860;
wire n_12430;
wire n_7072;
wire newNet_2520;
wire n_448;
wire n_31685;
wire n_31155;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_28_;
wire n_37229;
wire n_38400;
wire newNet_242;
wire n_31022;
wire n_30175;
wire n_21647;
wire n_35791;
wire n_6623;
wire n_16374;
wire n_21488;
wire n_8637;
wire n_44429;
wire FE_OCP_RBN1714_n_20734;
wire n_15275;
wire n_4225;
wire n_9440;
wire n_36321;
wire n_8169;
wire n_2055;
wire n_41412;
wire n_36444;
wire n_9581;
wire n_46345;
wire n_5130;
wire FE_RN_256_0;
wire n_23737;
wire n_19280;
wire n_19909;
wire n_8242;
wire n_43729;
wire n_39915;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_22_;
wire n_43780;
wire newNet_3723;
wire n_5651;
wire FE_OCPN954_n_44460;
wire newNet_2899;
wire n_21632;
wire n_16036;
wire n_31114;
wire n_13731;
wire n_23922;
wire n_14360;
wire n_35809;
wire n_20083;
wire FE_RN_1335_0;
wire n_12444;
wire n_7533;
wire n_23305;
wire n_4133;
wire newNet_463;
wire n_24095;
wire n_31162;
wire n_17105;
wire n_8104;
wire n_32130;
wire n_28102;
wire n_43894;
wire n_29345;
wire n_21937;
wire n_17832;
wire n_24677;
wire FE_RN_789_0;
wire FE_OCP_RBN2735_n_14985;
wire FE_OCPN1526_n_26587;
wire newNet_3268;
wire n_4964;
wire n_32660;
wire n_4932;
wire n_21475;
wire n_571;
wire FE_RN_364_0;
wire n_30167;
wire n_35622;
wire newNet_3503;
wire FE_RN_784_0;
wire n_3287;
wire n_28385;
wire n_36309;
wire n_47027;
wire n_33484;
wire n_22245;
wire n_29249;
wire n_2206;
wire sin_out_6;
wire FE_OCP_RBN3819_n_44061;
wire n_33721;
wire n_36063;
wire n_128;
wire newNet_2771;
wire n_3842;
wire n_41512;
wire n_39895;
wire n_26551;
wire n_2224;
wire FE_OCP_RBN3560_n_8809;
wire n_4544;
wire n_6346;
wire n_11952;
wire FE_RN_584_0;
wire n_45050;
wire n_18276;
wire FE_RN_1688_0;
wire n_33012;
wire n_43306;
wire n_41775;
wire delay_add_ln22_unr11_stage5_stallmux_q_30_;
wire n_2944;
wire newNet_334;
wire n_7393;
wire FE_OCP_RBN2494_n_8641;
wire FE_OCP_RBN2680_n_14768;
wire n_21620;
wire n_910;
wire n_5830;
wire n_7008;
wire n_3882;
wire n_3220;
wire n_30021;
wire newNet_3654;
wire n_17713;
wire n_15828;
wire n_20458;
wire n_5634;
wire n_33602;
wire n_6703;
wire FE_OCP_RBN3251_delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire n_466;
wire n_6607;
wire n_14220;
wire n_43120;
wire n_14345;
wire n_35312;
wire n_38308;
wire n_31505;
wire n_31140;
wire n_25062;
wire n_281;
wire n_28560;
wire n_9946;
wire n_8400;
wire n_8793;
wire n_2840;
wire n_38250;
wire n_24739;
wire FE_OCPN1765_n_33447;
wire n_25193;
wire FE_RN_825_0;
wire n_37434;
wire FE_OCP_RBN1723_n_21004;
wire n_2212;
wire n_28298;
wire n_42175;
wire n_43879;
wire delay_add_ln22_unr8_stage4_stallmux_q_27_;
wire n_6865;
wire newNet_2074;
wire n_29018;
wire n_26822;
wire delay_add_ln22_unr2_stage2_stallmux_q_3_;
wire n_35046;
wire FE_OCPN1443_n_45050;
wire n_44721;
wire n_14543;
wire n_30526;
wire FE_RN_302_0;
wire newNet_3524;
wire n_15856;
wire n_20041;
wire n_8710;
wire n_28913;
wire n_14962;
wire n_20198;
wire n_29546;
wire n_18505;
wire n_38256;
wire n_39236;
wire n_1728;
wire n_33101;
wire n_18743;
wire n_16445;
wire n_9013;
wire n_24570;
wire n_13096;
wire n_3047;
wire newNet_91;
wire n_42618;
wire n_41999;
wire n_27933;
wire FE_RN_1563_0;
wire n_39267;
wire n_28428;
wire newNet_2804;
wire n_11451;
wire n_7609;
wire n_20005;
wire n_11745;
wire n_15845;
wire n_18294;
wire n_22231;
wire n_36905;
wire n_1798;
wire n_30770;
wire newNet_194;
wire newNet_2116;
wire n_9526;
wire n_43097;
wire n_1003;
wire n_14351;
wire FE_OCP_RBN2522_n_8951;
wire n_1304;
wire n_23570;
wire n_7125;
wire n_23068;
wire FE_OCP_RBN3066_n_36547;
wire n_42627;
wire FE_RN_1380_0;
wire n_1044;
wire n_4654;
wire n_15342;
wire n_11220;
wire FE_OCP_RBN2433_n_14018;
wire n_2920;
wire delay_xor_ln21_unr3_stage2_stallmux_q_3_;
wire n_42398;
wire n_15235;
wire newNet_1460;
wire n_707;
wire FE_RN_1496_0;
wire n_14403;
wire newNet_2156;
wire FE_RN_1145_0;
wire n_9947;
wire n_21125;
wire n_27875;
wire newNet_73;
wire FE_OCP_RBN3725_n_16975;
wire n_19558;
wire n_23574;
wire n_6717;
wire n_17605;
wire FE_OCP_RBN3048_n_6013;
wire delay_add_ln22_unr11_stage5_stallmux_q_22_;
wire n_31692;
wire n_22705;
wire n_8849;
wire n_26553;
wire n_1452;
wire n_5700;
wire n_31816;
wire n_5853;
wire n_35069;
wire n_20654;
wire n_10149;
wire n_7959;
wire newNet_2853;
wire n_7563;
wire n_6417;
wire n_29013;
wire n_31100;
wire n_13035;
wire n_38603;
wire newNet_1213;
wire n_44083;
wire n_2226;
wire FE_OCP_DRV_N1552_n_19010;
wire n_41118;
wire FE_RN_870_0;
wire n_20002;
wire n_8091;
wire FE_OCP_RBN2630_n_14912;
wire n_36318;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_8_;
wire n_31716;
wire n_2979;
wire n_18288;
wire n_21530;
wire newNet_674;
wire n_4262;
wire n_20399;
wire n_8084;
wire newNet_3526;
wire newNet_2281;
wire n_9566;
wire n_18379;
wire n_22738;
wire FE_OFN841_n_15791;
wire n_36240;
wire n_27314;
wire n_31352;
wire newNet_2730;
wire n_15474;
wire n_7588;
wire n_38234;
wire delay_add_ln22_unr23_stage9_stallmux_q_12_;
wire n_1948;
wire n_17243;
wire n_16524;
wire newNet_346;
wire n_21810;
wire n_36982;
wire delay_sub_ln23_0_unr28_stage10_stallmux_q;
wire n_45894;
wire n_20542;
wire n_23697;
wire n_36356;
wire n_7240;
wire n_20096;
wire n_12434;
wire n_12530;
wire n_2999;
wire FE_OCP_RBN3040_n_46337;
wire n_31138;
wire FE_RN_704_0;
wire n_3398;
wire n_37307;
wire n_28066;
wire newNet_927;
wire n_13913;
wire newNet_1615;
wire delay_add_ln22_unr23_stage9_stallmux_q_30_;
wire n_36586;
wire n_5419;
wire n_24507;
wire n_42670;
wire n_37509;
wire n_7438;
wire n_35190;
wire n_2925;
wire n_38665;
wire n_39286;
wire FE_OCP_RBN1324_n_29056;
wire n_21341;
wire n_796;
wire n_10079;
wire n_39714;
wire n_20299;
wire n_41083;
wire newNet_1651;
wire n_35315;
wire n_28787;
wire n_26669;
wire n_2601;
wire n_34669;
wire n_29100;
wire n_10666;
wire n_32324;
wire n_12346;
wire n_31755;
wire n_21818;
wire n_11935;
wire n_11158;
wire n_8992;
wire n_41971;
wire FE_RN_1143_0;
wire n_22751;
wire newNet_2802;
wire FE_OCP_RBN3508_n_13860;
wire n_16379;
wire n_42534;
wire n_17389;
wire n_33746;
wire n_20559;
wire n_22803;
wire n_6655;
wire n_11715;
wire n_7001;
wire n_12566;
wire n_26165;
wire n_9650;
wire n_6261;
wire n_13277;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_12_;
wire n_21940;
wire FE_OCP_RBN3625_n_38870;
wire n_39348;
wire n_30179;
wire FE_OCP_RBN2264_n_29033;
wire n_43092;
wire n_298;
wire n_43504;
wire n_27375;
wire newNet_177;
wire n_2293;
wire n_40700;
wire n_42072;
wire n_27230;
wire n_39111;
wire FE_OCP_RBN1337_n_20941;
wire n_32343;
wire n_28508;
wire n_27559;
wire n_29354;
wire n_40907;
wire n_25029;
wire newNet_2531;
wire newNet_811;
wire n_29460;
wire n_31086;
wire n_6975;
wire n_35582;
wire n_5755;
wire n_12754;
wire n_41473;
wire n_24207;
wire n_26045;
wire n_3790;
wire n_31018;
wire n_4033;
wire n_40521;
wire n_24154;
wire n_26840;
wire n_5262;
wire FE_OCP_RBN2464_n_4336;
wire n_28700;
wire n_23712;
wire n_16257;
wire n_817;
wire n_12174;
wire n_28598;
wire newNet_2187;
wire n_28573;
wire n_30882;
wire FE_OCPN1776_n_18263;
wire n_28303;
wire n_33208;
wire n_32666;
wire n_8296;
wire newNet_2404;
wire n_1069;
wire n_32149;
wire n_22145;
wire n_4885;
wire n_39186;
wire n_26582;
wire n_4051;
wire n_692;
wire n_12040;
wire n_1643;
wire n_28734;
wire n_20549;
wire newNet_3071;
wire n_43003;
wire n_9484;
wire newNet_1458;
wire n_35152;
wire n_36890;
wire n_14857;
wire n_2912;
wire beta_15;
wire n_37222;
wire n_124;
wire n_11024;
wire n_35683;
wire n_28119;
wire n_20956;
wire n_10396;
wire n_14788;
wire n_5091;
wire n_14429;
wire n_22869;
wire n_26153;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_2_;
wire n_1923;
wire n_24184;
wire n_36625;
wire n_12011;
wire n_27661;
wire n_3788;
wire n_31395;
wire n_36049;
wire newNet_3074;
wire n_19669;
wire n_15380;
wire n_18676;
wire n_29132;
wire n_45505;
wire newNet_2323;
wire n_25724;
wire n_35906;
wire n_43310;
wire newNet_836;
wire n_522;
wire n_16388;
wire n_3212;
wire n_8699;
wire n_35383;
wire n_3359;
wire FE_OCP_DRV_N1576_n_28829;
wire FE_OCP_RBN3490_n_3390;
wire n_1422;
wire n_1794;
wire n_37077;
wire n_11097;
wire n_43053;
wire n_11194;
wire n_4843;
wire n_41717;
wire n_17104;
wire n_4927;
wire n_12081;
wire n_20053;
wire newNet_1842;
wire n_44877;
wire n_40452;
wire n_36916;
wire n_9505;
wire n_12914;
wire n_20581;
wire n_21682;
wire n_43830;
wire n_7702;
wire n_11272;
wire newNet_1528;
wire n_4221;
wire n_17201;
wire n_37631;
wire n_38355;
wire n_35339;
wire n_22458;
wire n_33758;
wire n_29772;
wire FE_OCPN1253_n_8348;
wire n_20441;
wire n_4276;
wire n_43225;
wire n_43542;
wire n_29526;
wire newNet_1387;
wire n_24273;
wire n_14368;
wire n_43892;
wire newNet_2695;
wire n_22233;
wire n_8489;
wire n_30849;
wire n_25049;
wire n_21495;
wire n_17837;
wire n_12235;
wire n_13769;
wire FE_RN_436_0;
wire n_18614;
wire newNet_356;
wire n_19772;
wire n_15895;
wire n_24845;
wire FE_OCP_RBN1182_n_19726;
wire n_25524;
wire n_41769;
wire n_42918;
wire FE_RN_1715_0;
wire n_29986;
wire n_40884;
wire n_17808;
wire n_3296;
wire n_12008;
wire n_30354;
wire FE_RN_989_0;
wire n_32689;
wire n_13140;
wire newNet_2058;
wire n_7964;
wire n_17180;
wire n_30614;
wire n_17121;
wire n_9720;
wire n_5072;
wire n_18935;
wire n_814;
wire n_14241;
wire n_11202;
wire n_33854;
wire n_15172;
wire n_5373;
wire n_40350;
wire newNet_571;
wire n_3378;
wire n_7820;
wire n_43759;
wire n_28767;
wire n_8522;
wire n_35026;
wire n_10073;
wire n_12370;
wire FE_OCP_RBN3212_n_44365;
wire n_35358;
wire n_14471;
wire n_39463;
wire n_32908;
wire newNet_443;
wire n_13634;
wire n_20036;
wire n_36429;
wire n_6032;
wire n_25102;
wire n_17576;
wire n_10832;
wire n_1158;
wire n_24070;
wire n_17993;
wire n_33199;
wire n_22294;
wire n_11779;
wire newNet_2980;
wire n_17266;
wire n_5382;
wire n_33070;
wire n_37159;
wire n_32363;
wire n_41902;
wire n_33714;
wire n_31686;
wire n_3324;
wire newNet_784;
wire newNet_1559;
wire n_23047;
wire n_19703;
wire n_37456;
wire n_21698;
wire n_5673;
wire n_44288;
wire n_24571;
wire n_35165;
wire newNet_1251;
wire n_17552;
wire FE_OCPN1751_n_29420;
wire n_37439;
wire n_4317;
wire n_5796;
wire n_29044;
wire n_24501;
wire n_16461;
wire n_28166;
wire n_38277;
wire n_43469;
wire n_28761;
wire newNet_195;
wire newNet_1744;
wire n_21933;
wire FE_RN_338_0;
wire n_2649;
wire n_30818;
wire n_26325;
wire n_42950;
wire n_11492;
wire newNet_171;
wire n_37325;
wire n_22053;
wire n_14556;
wire n_40559;
wire n_29929;
wire n_26960;
wire n_33258;
wire n_2669;
wire n_2624;
wire n_36360;
wire n_6830;
wire n_26736;
wire n_24396;
wire n_27578;
wire n_5461;
wire newNet_2288;
wire n_2014;
wire n_40815;
wire n_23045;
wire n_28144;
wire n_40432;
wire n_43895;
wire n_11068;
wire n_44344;
wire n_18215;
wire n_34693;
wire newNet_3640;
wire n_10721;
wire n_34454;
wire n_20710;
wire newNet_2475;
wire n_35228;
wire n_38571;
wire n_1774;
wire n_19391;
wire n_36772;
wire n_1943;
wire n_9744;
wire n_35451;
wire n_6635;
wire n_25187;
wire n_4554;
wire n_26081;
wire n_17714;
wire n_40741;
wire n_12026;
wire newNet_530;
wire n_21332;
wire n_6020;
wire n_23440;
wire n_35178;
wire n_6347;
wire n_10101;
wire n_39311;
wire n_34246;
wire n_24547;
wire n_15843;
wire n_10484;
wire n_5510;
wire n_25345;
wire n_33011;
wire n_13889;
wire n_10647;
wire n_33894;
wire n_39970;
wire newNet_3167;
wire n_1436;
wire n_2746;
wire newNet_590;
wire n_41288;
wire n_615;
wire n_14812;
wire n_48;
wire n_41522;
wire n_42423;
wire n_20578;
wire n_29751;
wire FE_RN_1132_0;
wire n_18884;
wire n_8427;
wire n_18148;
wire n_18855;
wire FE_RN_1169_0;
wire n_29407;
wire n_42180;
wire n_17448;
wire delay_xor_ln21_unr21_stage8_stallmux_q_5_;
wire n_39648;
wire n_6399;
wire n_40688;
wire n_726;
wire n_42750;
wire n_15192;
wire n_6304;
wire FE_OCP_RBN2186_n_37686;
wire n_25412;
wire n_25204;
wire n_11354;
wire n_12468;
wire n_12643;
wire FE_RN_1353_0;
wire n_39140;
wire n_14387;
wire n_22491;
wire n_37101;
wire n_41028;
wire n_34337;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_6_;
wire n_34101;
wire n_36550;
wire n_19435;
wire n_12140;
wire n_42314;
wire n_30537;
wire n_35808;
wire newNet_1130;
wire n_3273;
wire n_39866;
wire n_14723;
wire n_20877;
wire n_11701;
wire n_39441;
wire n_29802;
wire n_24970;
wire n_14474;
wire FE_RN_774_0;
wire n_33467;
wire n_20636;
wire n_38646;
wire n_21141;
wire newNet_387;
wire n_30459;
wire n_22875;
wire n_673;
wire n_36573;
wire n_31434;
wire n_2966;
wire n_30498;
wire n_22636;
wire FE_OCP_RBN2653_n_14684;
wire n_28469;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_13_;
wire n_12440;
wire n_31847;
wire n_43436;
wire newNet_3231;
wire n_41581;
wire FE_OCP_DRV_N1602_n_21639;
wire n_22428;
wire n_288;
wire n_41703;
wire n_42997;
wire newNet_203;
wire n_1206;
wire n_40123;
wire n_19897;
wire n_26862;
wire n_344;
wire n_40300;
wire n_11929;
wire newNet_2576;
wire n_36420;
wire n_12263;
wire n_18739;
wire n_39219;
wire FE_OCP_DRV_N1606_n_31445;
wire n_17366;
wire n_10568;
wire newNet_2879;
wire n_39779;
wire n_10060;
wire FE_OCP_RBN3140_n_6477;
wire n_11287;
wire n_30441;
wire n_7056;
wire n_18707;
wire n_6253;
wire n_2049;
wire n_19037;
wire n_18087;
wire n_239;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_2_;
wire n_7465;
wire n_1118;
wire n_31192;
wire n_38879;
wire n_13716;
wire n_3000;
wire delay_xor_ln22_unr12_stage5_stallmux_q_3_;
wire n_47211;
wire n_41238;
wire n_43754;
wire n_30721;
wire n_4609;
wire n_3981;
wire n_40472;
wire n_31824;
wire n_29077;
wire n_32573;
wire n_21174;
wire n_23993;
wire n_36938;
wire n_25916;
wire FE_OCP_RBN2480_n_8595;
wire FE_OCP_RBN3422_n_12879;
wire n_9439;
wire newNet_3349;
wire n_5216;
wire n_22407;
wire n_37864;
wire n_31331;
wire n_4204;
wire n_20210;
wire n_31560;
wire n_42147;
wire n_10020;
wire n_32682;
wire n_11189;
wire n_8302;
wire n_35086;
wire n_14438;
wire n_36432;
wire n_31064;
wire n_41731;
wire n_4243;
wire n_9305;
wire delay_add_ln22_unr8_stage4_stallmux_q_29_;
wire n_29547;
wire n_15499;
wire n_13788;
wire n_7625;
wire n_30919;
wire n_14023;
wire n_5937;
wire n_10006;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_13_;
wire FE_RN_188_0;
wire n_31759;
wire n_12803;
wire n_14442;
wire n_31258;
wire n_28905;
wire n_39211;
wire n_43271;
wire n_43752;
wire n_14144;
wire n_37806;
wire newNet_1163;
wire n_10230;
wire n_14108;
wire n_13658;
wire n_900;
wire n_34711;
wire FE_RN_1320_0;
wire n_29202;
wire FE_RN_1197_0;
wire delay_add_ln22_unr20_stage8_stallmux_q_2_;
wire n_43263;
wire FE_OCP_RBN3115_n_6379;
wire n_42189;
wire n_24405;
wire FE_OCP_RBN2765_n_25895;
wire n_12771;
wire n_27006;
wire FE_OCP_RBN2831_n_10198;
wire n_15577;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_10_;
wire n_24050;
wire n_3158;
wire n_46169;
wire n_1372;
wire n_22221;
wire n_7211;
wire FE_RN_1232_0;
wire n_19775;
wire n_30659;
wire n_32206;
wire n_30961;
wire n_26710;
wire n_4930;
wire n_10252;
wire n_29719;
wire n_24708;
wire n_45747;
wire n_11617;
wire FE_RN_591_0;
wire newNet_940;
wire n_3204;
wire n_41834;
wire n_854;
wire n_41991;
wire n_12271;
wire newNet_1783;
wire n_16575;
wire newNet_494;
wire n_4580;
wire n_23266;
wire FE_OCP_RBN1176_n_18981;
wire n_31223;
wire n_17233;
wire n_5436;
wire n_39074;
wire n_44636;
wire n_1354;
wire n_31160;
wire n_13576;
wire n_21134;
wire n_14954;
wire n_43267;
wire n_25563;
wire n_21421;
wire n_29940;
wire FE_RN_359_0;
wire n_36160;
wire n_20983;
wire n_1619;
wire newNet_1413;
wire n_1046;
wire n_18600;
wire FE_OCP_RBN3647_n_44490;
wire n_39741;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_1_;
wire n_35230;
wire n_227;
wire n_5609;
wire n_39797;
wire n_42748;
wire n_21476;
wire FE_OCP_RBN2305_n_7817;
wire n_33109;
wire n_31655;
wire n_1855;
wire n_35491;
wire n_17740;
wire FE_OCPN1417_n_31504;
wire n_4892;
wire n_13670;
wire newNet_139;
wire newNet_1591;
wire n_5909;
wire n_5428;
wire FE_RN_1704_0;
wire newNet_2632;
wire n_7405;
wire n_22034;
wire n_12553;
wire n_4391;
wire n_2488;
wire n_42359;
wire n_29144;
wire FE_OCP_RBN2644_n_34980;
wire n_8937;
wire newNet_2553;
wire newNet_2480;
wire n_20997;
wire n_41279;
wire n_21794;
wire n_20624;
wire n_7850;
wire n_11538;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_22_;
wire delay_xor_ln21_unr3_stage2_stallmux_q_24_;
wire FE_RN_1668_0;
wire newNet_2220;
wire n_16987;
wire n_36675;
wire n_17610;
wire n_1513;
wire n_2091;
wire newNet_1810;
wire n_6114;
wire n_5385;
wire n_26753;
wire n_23953;
wire n_20202;
wire n_11146;
wire n_38061;
wire n_25639;
wire n_31801;
wire n_18566;
wire n_42415;
wire n_33682;
wire n_115;
wire n_13588;
wire n_9694;
wire n_36397;
wire n_33391;
wire n_26708;
wire n_18559;
wire n_31243;
wire n_1312;
wire n_31494;
wire n_19873;
wire n_36539;
wire n_14798;
wire newNet_2270;
wire n_21181;
wire n_17302;
wire n_36358;
wire n_10856;
wire n_43010;
wire n_11675;
wire n_36437;
wire n_9839;
wire n_34861;
wire n_34122;
wire n_26290;
wire n_8825;
wire newNet_2224;
wire n_43032;
wire n_42838;
wire n_77;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_7_;
wire n_43721;
wire n_32315;
wire n_27274;
wire FE_OCPN1006_n_13962;
wire n_22843;
wire n_35840;
wire n_4146;
wire n_37808;
wire n_33911;
wire n_40097;
wire FE_OCPN1423_delay_sub_ln23_0_unr21_stage8_stallmux_q;
wire FE_RN_1525_0;
wire n_12375;
wire n_25195;
wire n_12664;
wire n_42478;
wire n_43115;
wire n_21045;
wire n_41245;
wire n_42859;
wire n_4158;
wire n_6177;
wire n_9782;
wire n_29279;
wire n_16415;
wire n_13425;
wire n_37369;
wire n_20889;
wire n_22777;
wire n_35525;
wire n_20385;
wire n_565;
wire n_42283;
wire n_8000;
wire n_34889;
wire n_41568;
wire n_41392;
wire n_42729;
wire n_2462;
wire newNet_619;
wire n_69;
wire n_22298;
wire FE_OCP_RBN2235_n_29055;
wire n_4186;
wire n_7491;
wire n_16337;
wire n_26213;
wire n_39848;
wire FE_OCP_RBN1137_n_11779;
wire n_40915;
wire n_11804;
wire n_41607;
wire n_19761;
wire newNet_274;
wire n_21915;
wire FE_RN_722_0;
wire FE_RN_157_0;
wire n_25030;
wire n_38930;
wire n_23911;
wire n_39725;
wire FE_RN_1677_0;
wire n_36228;
wire cos_out_14;
wire n_24254;
wire newNet_2312;
wire delay_sub_ln23_unr29_stage9_stallmux_q_2_;
wire n_24592;
wire n_543;
wire n_1502;
wire n_34994;
wire n_2790;
wire n_12242;
wire n_3855;
wire n_22089;
wire n_32529;
wire newNet_1866;
wire newNet_3554;
wire n_25362;
wire n_39732;
wire n_37762;
wire n_6130;
wire n_13675;
wire n_7284;
wire n_38779;
wire n_25404;
wire n_36445;
wire n_29007;
wire n_9659;
wire n_10575;
wire n_2322;
wire n_13398;
wire n_34510;
wire FE_OCP_RBN2991_n_35539;
wire newNet_408;
wire n_26176;
wire n_31763;
wire n_14970;
wire n_15696;
wire n_30423;
wire n_45194;
wire n_16532;
wire newNet_3498;
wire n_1560;
wire n_34896;
wire FE_OCPN3174_n_38799;
wire n_1182;
wire n_27767;
wire n_37687;
wire n_16049;
wire n_39891;
wire n_15963;
wire n_40889;
wire FE_OCP_RBN3640_n_44490;
wire n_22130;
wire n_21352;
wire n_25702;
wire newNet_1395;
wire n_45300;
wire n_25709;
wire n_21783;
wire n_13560;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_3_;
wire n_10153;
wire n_4039;
wire delay_add_ln22_unr27_stage10_stallmux_q_7_;
wire n_16977;
wire newNet_1184;
wire n_690;
wire n_7686;
wire n_9203;
wire newNet_3313;
wire n_33573;
wire n_25243;
wire delay_xor_ln21_unr9_stage4_stallmux_q_13_;
wire n_26544;
wire n_18104;
wire FE_RN_500_0;
wire n_6493;
wire n_7745;
wire n_5137;
wire n_38378;
wire n_34017;
wire n_39422;
wire n_13119;
wire n_41006;
wire n_21490;
wire n_43383;
wire n_26299;
wire n_39361;
wire n_4526;
wire n_26420;
wire n_6921;
wire n_42864;
wire n_36155;
wire n_4642;
wire n_8630;
wire n_4698;
wire newNet_1809;
wire newNet_3108;
wire n_26230;
wire n_18776;
wire n_6197;
wire FE_RN_1876_0;
wire n_41613;
wire FE_OCP_DRV_N1588_n_31012;
wire n_25019;
wire n_16866;
wire FE_RN_648_0;
wire n_42363;
wire n_19930;
wire n_6044;
wire FE_RN_200_0;
wire n_35920;
wire FE_RN_427_0;
wire n_20719;
wire n_23984;
wire FE_OCP_RBN2816_n_4459;
wire newNet_1455;
wire n_41226;
wire n_25396;
wire n_21569;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_28_;
wire n_7034;
wire n_22185;
wire n_30101;
wire FE_RN_1575_0;
wire n_38221;
wire n_8136;
wire n_42718;
wire FE_RN_1513_0;
wire n_37880;
wire n_18801;
wire n_14398;
wire n_16293;
wire n_7264;
wire n_38198;
wire FE_OCP_RBN2246_n_13017;
wire n_37010;
wire n_32198;
wire n_23976;
wire newNet_690;
wire n_24025;
wire n_41515;
wire n_11329;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_19_;
wire newNet_1580;
wire n_4624;
wire FE_OCP_RBN2367_n_24408;
wire n_4475;
wire n_27931;
wire n_8484;
wire n_22656;
wire n_30071;
wire n_21968;
wire n_12492;
wire n_34903;
wire newNet_3400;
wire n_38833;
wire newNet_2344;
wire n_14925;
wire n_14875;
wire n_14168;
wire n_14419;
wire n_40269;
wire n_33413;
wire n_650;
wire n_18358;
wire n_1425;
wire n_38421;
wire n_2043;
wire n_24196;
wire n_6867;
wire n_7349;
wire n_18948;
wire n_7902;
wire n_30429;
wire n_21500;
wire n_4703;
wire n_38260;
wire n_20846;
wire n_18714;
wire FE_OCP_RBN2884_n_26292;
wire n_24083;
wire n_11958;
wire n_33321;
wire n_18940;
wire n_27025;
wire n_21051;
wire FE_RN_1678_0;
wire FE_RN_987_0;
wire n_32501;
wire n_24797;
wire cos_out_26;
wire newNet_418;
wire FE_OCP_RBN3594_n_44561;
wire n_29935;
wire n_28710;
wire n_23937;
wire n_3744;
wire n_32078;
wire n_18420;
wire n_9794;
wire n_11051;
wire n_46137;
wire n_18971;
wire FE_OCP_RBN3025_n_39942;
wire n_34929;
wire n_35213;
wire n_15521;
wire n_2526;
wire newNet_2096;
wire newNet_688;
wire newNet_252;
wire n_387;
wire n_2231;
wire n_25514;
wire sin_out_19;
wire n_2712;
wire n_20243;
wire n_28858;
wire newNet_852;
wire n_43810;
wire FE_OCP_RBN2173_n_1813;
wire n_23766;
wire FE_OCP_RBN3079_n_16977;
wire n_22057;
wire n_43563;
wire n_10490;
wire n_21069;
wire n_40950;
wire n_2185;
wire n_2413;
wire n_16589;
wire n_24803;
wire n_4563;
wire n_40633;
wire n_16218;
wire newNet_1822;
wire n_44268;
wire n_32090;
wire n_18261;
wire n_33262;
wire n_41297;
wire n_42623;
wire newNet_1963;
wire n_35744;
wire n_45512;
wire n_8964;
wire n_45002;
wire n_32916;
wire n_34676;
wire n_27987;
wire n_36716;
wire n_23629;
wire n_19533;
wire delay_xor_ln22_unr18_stage7_stallmux_q_0_;
wire n_40518;
wire newNet_2719;
wire n_27696;
wire n_37747;
wire n_37726;
wire n_18592;
wire n_13552;
wire n_4363;
wire FE_RN_615_0;
wire newNet_1525;
wire n_17340;
wire newNet_3718;
wire n_842;
wire n_30266;
wire FE_RN_727_0;
wire newNet_126;
wire n_10868;
wire n_22528;
wire n_17297;
wire newNet_2079;
wire n_8538;
wire n_38327;
wire n_23467;
wire n_24101;
wire FE_RN_414_0;
wire n_34330;
wire n_38398;
wire n_33821;
wire n_15332;
wire n_5230;
wire n_5825;
wire FE_OCP_RBN2649_n_3840;
wire n_31371;
wire n_34725;
wire n_21087;
wire n_12949;
wire n_2383;
wire n_15836;
wire n_6096;
wire n_43140;
wire n_22354;
wire n_14668;
wire n_12696;
wire n_20793;
wire newNet_557;
wire n_4710;
wire n_43730;
wire n_34718;
wire n_11697;
wire FE_OCP_RBN2938_n_26456;
wire n_26882;
wire n_28657;
wire n_9447;
wire n_40361;
wire FE_OCP_RBN2956_n_26231;
wire n_37537;
wire n_21662;
wire n_21100;
wire n_28458;
wire n_44423;
wire n_33362;
wire n_29729;
wire n_28691;
wire n_32990;
wire n_14450;
wire n_20225;
wire n_1007;
wire n_40890;
wire n_2872;
wire n_40290;
wire n_42603;
wire newNet_3565;
wire n_34960;
wire n_10922;
wire n_22962;
wire newNet_3481;
wire n_38068;
wire n_31938;
wire n_11588;
wire n_27062;
wire n_32044;
wire n_41967;
wire FE_RN_1007_0;
wire n_38291;
wire n_28891;
wire n_1638;
wire n_40227;
wire n_21070;
wire n_11402;
wire n_42144;
wire n_20617;
wire n_13133;
wire FE_RN_884_0;
wire newNet_736;
wire n_19811;
wire n_14374;
wire n_32942;
wire n_34203;
wire delay_add_ln22_unr2_stage2_stallmux_q_20_;
wire n_5244;
wire n_26508;
wire n_20752;
wire n_23224;
wire n_26599;
wire n_15081;
wire FE_RN_873_0;
wire delay_xor_ln22_unr21_stage8_stallmux_q_1_;
wire n_9099;
wire newNet_3598;
wire FE_RN_1030_0;
wire FE_OCP_RBN2303_n_7817;
wire n_7966;
wire n_2317;
wire n_43579;
wire FE_OCPN877_n_44734;
wire n_32335;
wire n_13;
wire n_5748;
wire n_45738;
wire n_7169;
wire n_40319;
wire n_25058;
wire sin_out_23;
wire FE_OFN756_n_44461;
wire n_27482;
wire n_32624;
wire n_3177;
wire n_5946;
wire n_28634;
wire n_37737;
wire n_41637;
wire n_5211;
wire n_39143;
wire newNet_3642;
wire n_6266;
wire n_36346;
wire n_39667;
wire n_3686;
wire n_35776;
wire n_23757;
wire n_39407;
wire n_12472;
wire n_24265;
wire n_38450;
wire n_29670;
wire n_37666;
wire n_20026;
wire n_3634;
wire n_35663;
wire n_19087;
wire n_35757;
wire n_24326;
wire n_19793;
wire n_6668;
wire FE_OCPN3763_n_34222;
wire newNet_2027;
wire n_11986;
wire n_39665;
wire newNet_1200;
wire n_6146;
wire n_669;
wire n_2733;
wire n_40207;
wire FE_RN_250_0;
wire n_11295;
wire FE_OCP_RBN2874_n_10477;
wire n_23100;
wire FE_OCPN3782_n_16463;
wire n_34940;
wire n_2271;
wire newNet_3096;
wire newNet_2836;
wire n_13515;
wire n_215;
wire n_22625;
wire n_34540;
wire n_1259;
wire FE_RN_107_0;
wire n_4810;
wire n_25832;
wire n_17082;
wire n_23672;
wire n_1223;
wire n_34189;
wire n_33796;
wire newNet_2510;
wire n_40910;
wire n_27631;
wire FE_OCP_RBN3485_n_13667;
wire n_21380;
wire n_16632;
wire n_2038;
wire n_7271;
wire n_12783;
wire n_582;
wire n_34066;
wire n_39855;
wire n_5174;
wire n_32849;
wire n_33950;
wire n_34144;
wire n_35276;
wire newNet_438;
wire n_14826;
wire n_101;
wire FE_RN_847_0;
wire newNet_2594;
wire n_5521;
wire n_31098;
wire n_30990;
wire newNet_1299;
wire n_38409;
wire n_38092;
wire n_54;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_13_;
wire delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire n_12863;
wire n_4500;
wire n_38457;
wire n_24985;
wire n_20939;
wire n_38744;
wire n_27822;
wire n_13137;
wire n_41123;
wire n_29836;
wire n_29266;
wire n_31112;
wire n_20294;
wire newNet_2580;
wire newNet_1546;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_9_;
wire n_36204;
wire n_41741;
wire n_17514;
wire n_22558;
wire n_7162;
wire n_16317;
wire n_26792;
wire n_12873;
wire n_26068;
wire beta_18;
wire newNet_2463;
wire n_46953;
wire n_20371;
wire n_5116;
wire n_7636;
wire n_39473;
wire n_20161;
wire newNet_3251;
wire n_6463;
wire newNet_3306;
wire n_6756;
wire n_11964;
wire newNet_298;
wire newNet_3058;
wire n_6340;
wire n_6740;
wire n_22944;
wire n_39783;
wire n_43791;
wire n_42648;
wire n_33317;
wire n_41892;
wire n_23483;
wire n_10555;
wire n_22466;
wire n_24740;
wire n_34698;
wire newNet_973;
wire n_29956;
wire FE_RN_1613_0;
wire n_24069;
wire n_47278;
wire n_20098;
wire n_33600;
wire n_27156;
wire n_26296;
wire n_8158;
wire n_21636;
wire n_29533;
wire n_1931;
wire n_31967;
wire n_27226;
wire n_19195;
wire n_14489;
wire n_9888;
wire FE_OCP_RBN2901_n_44174;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_21_;
wire FE_OCPN1446_n_31473;
wire n_247;
wire n_41270;
wire FE_OCP_RBN3799_delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire n_40949;
wire FE_RN_821_0;
wire FE_RN_864_0;
wire cos_out_17;
wire n_11212;
wire n_47182;
wire n_27692;
wire n_38973;
wire n_5707;
wire n_27587;
wire n_24034;
wire n_2695;
wire n_29129;
wire FE_OCP_RBN2208_n_12907;
wire n_32723;
wire n_18205;
wire n_19049;
wire newNet_1858;
wire n_27357;
wire n_3238;
wire n_9574;
wire n_43592;
wire n_14339;
wire n_38964;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_29_;
wire FE_RN_963_0;
wire n_39251;
wire n_5345;
wire n_18694;
wire n_36293;
wire delay_xor_ln22_unr15_stage6_stallmux_q_2_;
wire FE_RN_1526_0;
wire n_17580;
wire n_25167;
wire n_8082;
wire FE_RN_1833_0;
wire newNet_220;
wire n_21370;
wire FE_OCP_RBN2665_n_35207;
wire n_20908;
wire n_17786;
wire n_35574;
wire n_32630;
wire n_6395;
wire n_28951;
wire n_8857;
wire newNet_3202;
wire n_3393;
wire n_38249;
wire n_6569;
wire FE_OCP_RBN3727_FE_RN_1787_0;
wire n_33817;
wire n_42569;
wire newNet_119;
wire n_826;
wire n_5294;
wire n_31547;
wire n_13877;
wire n_24311;
wire n_10206;
wire FE_OCP_RBN2355_n_13858;
wire n_24672;
wire n_27935;
wire n_9666;
wire n_32033;
wire n_24010;
wire n_22654;
wire newNet_2954;
wire FE_OCPN1488_n_23447;
wire newNet_3249;
wire n_37672;
wire newNet_257;
wire delay_add_ln22_unr27_stage10_stallmux_q_28_;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_19_;
wire n_4616;
wire FE_OCP_RBN3284_n_44365;
wire n_42842;
wire n_1301;
wire n_9142;
wire FE_OFN804_n_46196;
wire n_15858;
wire n_37526;
wire newNet_1357;
wire n_12764;
wire FE_RN_1290_0;
wire n_45841;
wire n_19237;
wire n_24448;
wire n_6055;
wire FE_RN_276_0;
wire newNet_1207;
wire n_19273;
wire n_15482;
wire n_7526;
wire n_18989;
wire n_39483;
wire n_6721;
wire n_36921;
wire newNet_2003;
wire n_18051;
wire n_25151;
wire n_11141;
wire n_27714;
wire n_29815;
wire n_44797;
wire FE_OCP_RBN1164_n_13726;
wire n_38231;
wire n_36182;
wire n_13506;
wire n_12335;
wire n_30208;
wire n_2642;
wire n_6856;
wire n_39102;
wire n_28153;
wire FE_RN_112_0;
wire n_29083;
wire n_21516;
wire n_8725;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_29_;
wire n_36277;
wire n_24479;
wire newNet_3134;
wire FE_OCP_RBN1368_n_20763;
wire n_12365;
wire FE_RN_24_0;
wire n_12684;
wire n_19321;
wire n_39041;
wire newNet_3092;
wire n_11519;
wire n_40527;
wire n_28319;
wire newNet_1578;
wire n_39968;
wire newNet_2332;
wire n_10907;
wire FE_OCP_RBN2532_n_47018;
wire n_15004;
wire n_20282;
wire n_40587;
wire n_4252;
wire n_6585;
wire n_5596;
wire n_315;
wire n_38486;
wire newNet_1687;
wire n_12424;
wire n_24587;
wire n_3887;
wire n_22150;
wire n_15888;
wire n_39940;
wire n_35878;
wire FE_OCP_RBN2244_n_13017;
wire n_12628;
wire n_16715;
wire n_40992;
wire FE_OCP_RBN2894_n_39575;
wire newNet_770;
wire n_16710;
wire n_33201;
wire n_36785;
wire n_33354;
wire newNet_3561;
wire delay_sub_ln22_unr24_stage9_stallmux_q_2_;
wire n_12353;
wire n_40987;
wire n_31364;
wire n_22574;
wire n_42253;
wire FE_RN_682_0;
wire n_34981;
wire n_27879;
wire n_31421;
wire n_42442;
wire FE_RN_1788_0;
wire n_30163;
wire n_5923;
wire newNet_1919;
wire n_8720;
wire n_34232;
wire n_11606;
wire n_3957;
wire n_28534;
wire n_40459;
wire FE_OCP_RBN1141_n_25816;
wire n_42737;
wire n_21828;
wire n_13213;
wire n_26605;
wire n_22629;
wire n_4388;
wire n_6997;
wire n_9951;
wire n_36234;
wire n_41593;
wire n_9457;
wire n_42434;
wire n_42686;
wire n_14697;
wire n_32959;
wire n_16224;
wire n_34220;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_18_;
wire n_31700;
wire n_23370;
wire n_38480;
wire n_39110;
wire n_4305;
wire newNet_1442;
wire n_36651;
wire n_24149;
wire delay_xor_ln22_unr6_stage3_stallmux_q_0_;
wire n_24777;
wire newNet_869;
wire n_1218;
wire n_36497;
wire n_28212;
wire n_7265;
wire n_40365;
wire n_28220;
wire n_31688;
wire n_46191;
wire n_7120;
wire n_33453;
wire newNet_287;
wire n_116;
wire FE_OFN815_n_19807;
wire n_21452;
wire n_19271;
wire n_19698;
wire n_21987;
wire n_40714;
wire n_31412;
wire n_7233;
wire FE_RN_693_0;
wire FE_OCP_RBN3036_n_47269;
wire n_27676;
wire n_29725;
wire n_16066;
wire newNet_3370;
wire newNet_1448;
wire n_43319;
wire n_29048;
wire n_14754;
wire n_8805;
wire n_39072;
wire n_7943;
wire n_8043;
wire newNet_180;
wire n_41235;
wire n_856;
wire n_22648;
wire FE_RN_878_0;
wire n_39426;
wire n_28032;
wire n_2209;
wire n_10307;
wire n_40789;
wire FE_RN_1341_0;
wire n_19191;
wire n_43277;
wire n_18167;
wire n_30900;
wire n_19402;
wire FE_OCP_RBN3851_n_20848;
wire n_4058;
wire newNet_1893;
wire n_11624;
wire n_12561;
wire FE_RN_1743_0;
wire FE_OCP_RBN2842_n_4784;
wire n_15050;
wire FE_OCP_RBN3510_n_19599;
wire n_36637;
wire n_6447;
wire n_40211;
wire FE_OCPN1008_n_28439;
wire n_18047;
wire n_26363;
wire newNet_3255;
wire n_9806;
wire n_24818;
wire n_40914;
wire n_19894;
wire n_24049;
wire n_14424;
wire n_13941;
wire n_23097;
wire newNet_2881;
wire n_14468;
wire n_20641;
wire n_39781;
wire n_4658;
wire n_6626;
wire n_3974;
wire n_5843;
wire n_5941;
wire n_13421;
wire n_33461;
wire newNet_694;
wire FE_OCPUNCON1804_n_18111;
wire n_35819;
wire n_27780;
wire n_40182;
wire n_27200;
wire n_4018;
wire n_42033;
wire n_22635;
wire n_1732;
wire n_444;
wire n_23826;
wire newNet_1988;
wire n_29865;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_19_;
wire n_31227;
wire n_7010;
wire n_31858;
wire n_16350;
wire n_47001;
wire newNet_3207;
wire n_30857;
wire newNet_518;
wire n_10852;
wire n_12170;
wire n_25083;
wire n_26915;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_27_;
wire n_12770;
wire n_22747;
wire n_31775;
wire n_17597;
wire n_8756;
wire n_41793;
wire FE_OCPN1477_n_28775;
wire n_12668;
wire n_38135;
wire FE_OCP_RBN2756_FE_RN_722_0;
wire n_10176;
wire n_39914;
wire n_16749;
wire n_43187;
wire newNet_1720;
wire n_42810;
wire n_31481;
wire n_35221;
wire n_1610;
wire n_28817;
wire n_26204;
wire n_24291;
wire n_26526;
wire n_2503;
wire newNet_3639;
wire n_37623;
wire n_31341;
wire n_37440;
wire n_21744;
wire newNet_404;
wire n_17840;
wire FE_OCP_RBN2578_n_47017;
wire n_38678;
wire n_37041;
wire n_1815;
wire n_5335;
wire n_1956;
wire n_8288;
wire n_18153;
wire n_43430;
wire n_22989;
wire n_5995;
wire n_3571;
wire n_27600;
wire n_10096;
wire n_3955;
wire n_2728;
wire n_9631;
wire n_24997;
wire n_4371;
wire n_17008;
wire n_17306;
wire n_12018;
wire newNet_3317;
wire n_23339;
wire n_28780;
wire n_32855;
wire n_335;
wire n_26412;
wire FE_OCPN1255_n_8499;
wire n_29340;
wire n_13315;
wire n_3997;
wire n_36453;
wire n_14506;
wire n_4719;
wire n_12590;
wire n_4081;
wire FE_OCP_RBN3467_n_7886;
wire n_25649;
wire n_24894;
wire n_19500;
wire n_32072;
wire n_3223;
wire n_28894;
wire n_34892;
wire newNet_1706;
wire n_4192;
wire n_23490;
wire n_36955;
wire n_9366;
wire n_30965;
wire n_2329;
wire FE_RN_657_0;
wire FE_OCP_RBN3460_n_7886;
wire n_12058;
wire n_24815;
wire newNet_2103;
wire n_8889;
wire n_34879;
wire n_36255;
wire n_18754;
wire n_12397;
wire n_7926;
wire n_43622;
wire n_31606;
wire n_21866;
wire n_7799;
wire n_34350;
wire n_37453;
wire n_26648;
wire n_39229;
wire n_20715;
wire newNet_210;
wire newNet_1285;
wire n_970;
wire n_16518;
wire FE_OCP_DRV_N3740_n_29576;
wire n_1734;
wire newNet_2049;
wire n_18339;
wire n_28865;
wire newNet_3439;
wire n_25973;
wire newNet_540;
wire FE_RN_1324_0;
wire n_12613;
wire n_23138;
wire n_42289;
wire n_43242;
wire n_2792;
wire n_31898;
wire n_14933;
wire n_19380;
wire FE_OCP_RBN2777_n_15595;
wire n_36408;
wire n_33906;
wire n_8239;
wire n_913;
wire n_7411;
wire n_31071;
wire n_17441;
wire n_10211;
wire n_39518;
wire n_21111;
wire n_10116;
wire FE_OCP_RBN3441_n_37945;
wire n_3995;
wire n_38812;
wire n_37940;
wire n_43783;
wire n_22027;
wire n_20682;
wire n_7693;
wire n_19348;
wire newNet_1550;
wire n_11664;
wire newNet_524;
wire n_8028;
wire n_26359;
wire n_3343;
wire newNet_2685;
wire n_7194;
wire n_2751;
wire n_9857;
wire n_8511;
wire n_36527;
wire FE_OCP_RBN3050_n_11329;
wire n_2539;
wire FE_OCP_RBN1342_n_19077;
wire n_2685;
wire n_29631;
wire n_11997;
wire n_35044;
wire n_32203;
wire n_41526;
wire newNet_919;
wire n_45080;
wire n_12849;
wire FE_OCP_RBN1165_n_13726;
wire n_32481;
wire n_43411;
wire newNet_2436;
wire n_7503;
wire n_20688;
wire n_992;
wire n_34071;
wire newNet_1504;
wire n_8979;
wire n_3368;
wire n_37143;
wire n_13400;
wire n_14611;
wire FE_OFN507_n_25938;
wire n_44498;
wire n_30105;
wire newNet_283;
wire n_28190;
wire newNet_2425;
wire n_8037;
wire n_7628;
wire n_7477;
wire n_26935;
wire newNet_394;
wire n_14529;
wire n_31044;
wire n_13694;
wire n_34627;
wire n_17986;
wire n_34952;
wire n_3669;
wire n_45322;
wire n_11126;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_19_;
wire n_28834;
wire n_8821;
wire FE_OCP_RBN2883_n_26292;
wire n_25556;
wire n_30510;
wire n_37508;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_20_;
wire n_13808;
wire FE_RN_254_0;
wire n_1690;
wire n_11199;
wire n_42795;
wire n_41043;
wire n_35933;
wire n_16731;
wire n_28898;
wire n_4233;
wire n_24382;
wire FE_OCPN1441_n_45060;
wire FE_RN_1138_0;
wire n_25599;
wire n_22810;
wire delay_add_ln22_unr5_stage3_stallmux_q_12_;
wire n_1474;
wire n_13609;
wire n_20349;
wire newNet_2145;
wire n_10930;
wire n_39408;
wire n_31251;
wire n_42798;
wire n_13296;
wire n_41924;
wire n_36860;
wire n_34145;
wire n_11646;
wire n_33331;
wire n_42898;
wire n_3797;
wire n_4439;
wire n_25222;
wire n_12674;
wire n_46969;
wire n_17661;
wire n_28704;
wire n_23682;
wire n_4887;
wire newNet_2265;
wire n_34651;
wire newNet_1009;
wire n_28009;
wire n_4994;
wire n_40381;
wire n_5712;
wire n_42883;
wire n_13602;
wire n_8660;
wire n_36855;
wire FE_OCP_RBN3127_n_43752;
wire n_15126;
wire n_164;
wire n_28762;
wire n_7030;
wire n_37665;
wire n_1648;
wire n_4775;
wire n_17951;
wire n_5324;
wire FE_RN_1839_0;
wire n_1441;
wire n_20501;
wire n_25575;
wire n_43191;
wire n_15905;
wire n_14848;
wire FE_OCP_RBN1697_n_19206;
wire n_22593;
wire n_21226;
wire n_11415;
wire FE_RN_1330_0;
wire n_1678;
wire n_28128;
wire FE_OCP_RBN2633_n_30170;
wire n_34041;
wire n_3862;
wire n_30875;
wire n_34819;
wire n_35952;
wire FE_OCPN902_n_44581;
wire n_20469;
wire n_5554;
wire n_3768;
wire n_6002;
wire n_29894;
wire FE_OCP_RBN1922_cordic_combinational_sub_ln23_0_unr12_z_0__;
wire n_16077;
wire n_18024;
wire n_42850;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_24_;
wire n_5122;
wire newNet_1310;
wire FE_RN_761_0;
wire n_17144;
wire n_9643;
wire n_40865;
wire n_2532;
wire n_7555;
wire FE_OCP_DRV_N1553_n_19314;
wire n_35729;
wire n_27495;
wire n_11286;
wire n_38900;
wire n_41161;
wire n_39693;
wire n_8479;
wire FE_RN_18_0;
wire FE_RN_1010_0;
wire FE_OCP_RBN3118_n_22755;
wire n_32729;
wire n_30529;
wire n_26477;
wire n_23633;
wire n_10978;
wire n_40389;
wire n_19052;
wire n_34130;
wire n_1838;
wire n_41753;
wire n_38896;
wire n_14756;
wire n_6576;
wire n_21648;
wire n_3163;
wire n_16952;
wire n_36529;
wire newNet_1092;
wire n_36172;
wire n_42059;
wire n_9463;
wire n_24715;
wire n_18832;
wire n_1282;
wire n_32122;
wire n_9253;
wire n_13625;
wire n_41177;
wire n_6382;
wire n_27117;
wire n_15712;
wire FE_RN_828_0;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_14_;
wire FE_RN_1869_0;
wire n_509;
wire FE_RN_1025_0;
wire n_3123;
wire n_23189;
wire n_3616;
wire n_10737;
wire FE_RN_962_0;
wire n_34654;
wire n_4168;
wire n_9907;
wire n_3568;
wire n_13885;
wire n_18795;
wire newNet_715;
wire n_15310;
wire n_14944;
wire n_28305;
wire n_45635;
wire n_36373;
wire n_33231;
wire n_19541;
wire newNet_1043;
wire n_17377;
wire n_25171;
wire FE_RN_455_0;
wire n_33055;
wire newNet_2729;
wire n_2337;
wire n_7679;
wire newNet_2442;
wire n_5177;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_10_;
wire FE_RN_925_0;
wire delay_add_ln22_unr2_stage2_stallmux_q_21_;
wire n_35834;
wire n_38316;
wire FE_RN_61_0;
wire n_20754;
wire n_5527;
wire n_14091;
wire newNet_3576;
wire newNet_2352;
wire n_12053;
wire n_17130;
wire n_23998;
wire newNet_3634;
wire newNet_763;
wire n_23864;
wire FE_OCPUNCON3146_n_21058;
wire n_16431;
wire n_25525;
wire n_1823;
wire n_21712;
wire n_11690;
wire n_13569;
wire n_30481;
wire n_26185;
wire n_10792;
wire n_17159;
wire n_22888;
wire n_1360;
wire n_22701;
wire n_21947;
wire n_4976;
wire n_11078;
wire n_22712;
wire n_558;
wire n_6135;
wire n_19889;
wire n_38994;
wire n_17781;
wire n_1177;
wire n_12484;
wire n_20435;
wire n_26281;
wire newNet_2088;
wire n_43127;
wire FE_RN_1134_0;
wire FE_OCP_RBN3602_n_3913;
wire FE_OCPN1046_n_13570;
wire n_22436;
wire n_15586;
wire n_5964;
wire n_7363;
wire n_41332;
wire n_30546;
wire FE_RN_390_0;
wire n_24074;
wire n_39748;
wire newNet_8;
wire n_96;
wire n_8277;
wire newNet_1276;
wire FE_OCPN1254_n_8499;
wire n_26119;
wire n_18256;
wire n_42122;
wire n_20820;
wire n_32492;
wire n_31200;
wire n_21015;
wire n_1405;
wire n_42134;
wire n_11802;
wire FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire newNet_1170;
wire n_39448;
wire n_14104;
wire n_37775;
wire n_34161;
wire FE_OCP_RBN2912_n_30908;
wire n_1096;
wire n_35264;
wire n_15157;
wire n_13937;
wire n_35687;
wire n_34423;
wire FE_RN_1146_0;
wire n_32904;
wire newNet_1064;
wire n_405;
wire n_34597;
wire n_39927;
wire n_38460;
wire n_30591;
wire n_3101;
wire n_258;
wire n_27218;
wire n_29031;
wire n_37471;
wire n_34756;
wire n_22852;
wire n_32735;
wire newNet_1111;
wire n_659;
wire n_21090;
wire n_21936;
wire n_18302;
wire n_1765;
wire n_43539;
wire n_5354;
wire n_807;
wire FE_OCPN1452_n_27518;
wire n_36960;
wire n_30476;
wire n_24946;
wire n_12586;
wire n_28219;
wire n_3138;
wire n_15648;
wire n_7353;
wire n_17884;
wire n_5003;
wire n_32302;
wire n_27836;
wire n_38142;
wire n_39154;
wire n_25431;
wire n_14591;
wire n_39008;
wire FE_OCP_RBN2664_n_20333;
wire n_7516;
wire FE_OCP_RBN3608_n_14905;
wire n_317;
wire newNet_1108;
wire n_15958;
wire n_5767;
wire n_42427;
wire n_9028;
wire n_40753;
wire n_20006;
wire delay_xor_ln22_unr12_stage5_stallmux_q_5_;
wire n_23906;
wire newNet_549;
wire n_23249;
wire n_23631;
wire n_28465;
wire n_8719;
wire FE_OCP_RBN2103_n_44962;
wire n_23724;
wire n_36352;
wire n_17776;
wire n_11879;
wire n_41779;
wire FE_OCP_RBN2596_n_25181;
wire n_24379;
wire n_35477;
wire n_18019;
wire n_41838;
wire n_40416;
wire n_2981;
wire n_31553;
wire n_17347;
wire n_9547;
wire FE_RN_1178_0;
wire newNet_2605;
wire n_284;
wire n_11292;
wire newNet_2212;
wire n_19809;
wire n_5955;
wire n_22785;
wire newNet_628;
wire n_20991;
wire n_14586;
wire n_2866;
wire FE_RN_44_0;
wire newNet_3749;
wire n_11261;
wire n_39393;
wire n_19825;
wire n_10826;
wire n_30599;
wire n_38986;
wire FE_OCPN1514_FE_OFN738_n_22641;
wire n_41626;
wire newNet_1971;
wire n_5914;
wire n_16465;
wire n_12570;
wire n_13826;
wire n_45486;
wire n_13664;
wire FE_OCP_RBN1684_n_33491;
wire n_28852;
wire n_13287;
wire n_16733;
wire n_37515;
wire n_15704;
wire n_21339;
wire n_9606;
wire n_37300;
wire n_13376;
wire n_18412;
wire FE_OCP_RBN2710_n_35075;
wire FE_RN_1199_0;
wire FE_OCP_RBN1209_n_16814;
wire n_39130;
wire n_31325;
wire n_9358;
wire delay_xor_ln21_unr6_stage3_stallmux_q_9_;
wire n_38606;
wire n_23988;
wire n_9638;
wire n_10694;
wire n_18703;
wire newNet_2831;
wire n_40343;
wire n_20873;
wire newNet_1922;
wire n_6271;
wire n_31380;
wire delay_xor_ln21_unr3_stage2_stallmux_q_23_;
wire n_863;
wire n_10561;
wire n_43352;
wire n_10340;
wire newNet_884;
wire n_2000;
wire n_7570;
wire n_5426;
wire FE_OCP_RBN3611_FE_OCPN1797_n_20333;
wire n_619;
wire n_7597;
wire n_8832;
wire newNet_167;
wire n_3174;
wire n_31295;
wire n_9714;
wire n_10134;
wire n_13441;
wire n_40554;
wire n_8131;
wire FE_RN_239_0;
wire n_33160;
wire n_35055;
wire n_4116;
wire n_38388;
wire newNet_1249;
wire n_2469;
wire n_14975;
wire n_17608;
wire n_6017;
wire n_10902;
wire n_41302;
wire FE_OCP_RBN2728_n_4219;
wire n_18537;
wire n_37348;
wire n_33425;
wire n_11656;
wire FE_OCP_RBN2191_n_28597;
wire n_35496;
wire n_13614;
wire newNet_1134;
wire n_2358;
wire n_10974;
wire FE_RN_837_0;
wire newNet_1684;
wire n_19062;
wire FE_OCPN1479_n_23872;
wire n_14434;
wire n_28030;
wire newNet_1392;
wire n_43807;
wire n_36734;
wire newNet_2168;
wire delay_xor_ln22_unr6_stage3_stallmux_q_21_;
wire n_34328;
wire n_30336;
wire newNet_3342;
wire FE_OCP_RBN3516_n_8498;
wire FE_OCPN1487_n_23447;
wire n_33960;
wire n_18660;
wire n_21007;
wire n_32422;
wire n_42712;
wire n_20742;
wire n_34129;
wire n_1123;
wire n_10167;
wire n_11941;
wire n_9517;
wire n_1379;
wire n_5481;
wire n_8925;
wire FE_RN_361_0;
wire n_30554;
wire n_46374;
wire n_31998;
wire n_8390;
wire n_42910;
wire n_40963;
wire n_13305;
wire n_26774;
wire n_38664;
wire n_16287;
wire FE_OCP_RBN2698_n_4238;
wire n_36513;
wire n_10180;
wire FE_RN_1514_0;
wire n_5451;
wire n_36824;
wire n_8864;
wire newNet_310;
wire n_37073;
wire newNet_2615;
wire n_38753;
wire cos_out_5;
wire n_4160;
wire n_11772;
wire n_13414;
wire n_3408;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_22_;
wire n_34962;
wire n_2256;
wire n_46204;
wire n_22404;
wire n_35466;
wire n_40733;
wire n_30244;
wire newNet_2170;
wire n_13113;
wire n_37857;
wire n_20913;
wire n_25075;
wire n_23528;
wire FE_RN_1231_0;
wire n_34481;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_2_;
wire n_22523;
wire n_34812;
wire n_11320;
wire n_23878;
wire n_22328;
wire n_12722;
wire n_38762;
wire n_14002;
wire n_30046;
wire n_3630;
wire n_31054;
wire n_19986;
wire n_19691;
wire n_3705;
wire n_41376;
wire n_23386;
wire n_36381;
wire n_1594;
wire n_10861;
wire n_37057;
wire n_5642;
wire n_7069;
wire n_5102;
wire n_28203;
wire n_29270;
wire n_21507;
wire n_32287;
wire n_25349;
wire n_42948;
wire n_2829;
wire FE_OCP_RBN3732_n_31819;
wire n_32433;
wire n_19080;
wire n_33083;
wire n_7855;
wire n_27611;
wire n_43708;
wire n_19431;
wire delay_xor_ln21_unr3_stage2_stallmux_q_15_;
wire n_2494;
wire n_43550;
wire n_10717;
wire n_32980;
wire n_14076;
wire n_633;
wire n_42699;
wire FE_OCP_RBN3333_n_44962;
wire n_23424;
wire n_24648;
wire FE_OCP_RBN2635_n_38806;
wire n_25233;
wire n_24876;
wire n_37560;
wire n_39802;
wire n_16826;
wire n_15479;
wire n_15806;
wire n_29968;
wire n_1134;
wire newNet_1188;
wire n_19512;
wire n_15638;
wire FE_RN_369_0;
wire n_12278;
wire n_29580;
wire n_26943;
wire FE_RN_995_0;
wire n_32462;
wire n_10525;
wire n_40851;
wire n_44155;
wire n_29403;
wire n_41010;
wire n_37725;
wire n_6784;
wire n_2109;
wire n_23359;
wire FE_OCP_RBN2599_n_34388;
wire n_16103;
wire n_11555;
wire n_24625;
wire n_12810;
wire n_37004;
wire n_1475;
wire n_41885;
wire n_3036;
wire n_8245;
wire n_19138;
wire newNet_3097;
wire n_44568;
wire newNet_2374;
wire n_40496;
wire n_44033;
wire FE_OCPN3797_n_26115;
wire n_26061;
wire n_9930;
wire n_1785;
wire n_42491;
wire n_38153;
wire n_7771;
wire n_6868;
wire n_13038;
wire n_7784;
wire n_3496;
wire n_6775;
wire n_8732;
wire n_42397;
wire n_38123;
wire n_28729;
wire n_37918;
wire n_13989;
wire n_27684;
wire n_42469;
wire delay_add_ln22_unr20_stage8_stallmux_q_18_;
wire n_26579;
wire n_18451;
wire FE_OCP_RBN2931_n_5307;
wire newNet_2825;
wire n_4750;
wire n_6222;
wire n_18736;
wire n_33589;
wire n_26908;
wire n_29143;
wire n_29662;
wire n_9405;
wire n_23297;
wire n_20726;
wire n_13959;
wire n_30790;
wire n_26536;
wire n_30224;
wire newNet_3035;
wire n_13241;
wire n_17693;
wire FE_RN_1603_0;
wire n_1203;
wire n_13745;
wire n_2484;
wire n_2804;
wire FE_RN_208_0;
wire n_5815;
wire n_12284;
wire n_25421;
wire n_32176;
wire delay_add_ln22_unr2_stage2_stallmux_q_7_;
wire n_29883;
wire n_4530;
wire n_37488;
wire n_33491;
wire n_31564;
wire n_19574;
wire n_41585;
wire newNet_2734;
wire n_30604;
wire n_12868;
wire FE_RN_921_0;
wire n_41425;
wire FE_RN_1122_0;
wire FE_OCPN1521_n_26054;
wire n_43844;
wire n_29194;
wire FE_RN_1249_0;
wire n_31751;
wire n_22553;
wire n_33700;
wire n_21485;
wire n_4207;
wire n_42886;
wire newNet_3586;
wire n_32382;
wire FE_RN_1641_0;
wire n_25386;
wire n_24601;
wire n_37744;
wire FE_OCP_RBN2233_n_13141;
wire n_7083;
wire n_37241;
wire n_11087;
wire n_36515;
wire n_34617;
wire n_23895;
wire FE_RN_220_0;
wire n_32129;
wire n_26158;
wire n_24029;
wire n_39479;
wire n_39586;
wire n_40404;
wire n_19143;
wire n_27476;
wire newNet_758;
wire n_40855;
wire n_24164;
wire newNet_906;
wire n_1846;
wire n_32565;
wire n_31119;
wire n_28668;
wire n_35217;
wire FE_RN_1130_0;
wire n_31002;
wire FE_OCP_RBN2488_n_3338;
wire newNet_3331;
wire FE_OCP_RBN2838_n_4692;
wire n_20574;
wire n_20599;
wire newNet_621;
wire n_18126;
wire n_21034;
wire n_7156;
wire n_22287;
wire n_35113;
wire n_23376;
wire n_16206;
wire n_17863;
wire n_2304;
wire newNet_2456;
wire n_37447;
wire n_15283;
wire n_25851;
wire newNet_3261;
wire FE_RN_1595_0;
wire n_17023;
wire n_24921;
wire FE_RN_1481_0;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_10_;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_25_;
wire n_3058;
wire n_36749;
wire n_34262;
wire n_1913;
wire n_13458;
wire delay_add_ln22_unr5_stage3_stallmux_q_29_;
wire n_40643;
wire n_37359;
wire n_24341;
wire n_30823;
wire n_22995;
wire n_14533;
wire n_13797;
wire n_42825;
wire n_3639;
wire n_3084;
wire n_15227;
wire n_3313;
wire n_35303;
wire newNet_2544;
wire n_18851;
wire n_13364;
wire n_36220;
wire n_6327;
wire newNet_3478;
wire n_24933;
wire n_34547;
wire n_4741;
wire n_42970;
wire n_38506;
wire n_3328;
wire n_40812;
wire n_19943;
wire n_35097;
wire n_547;
wire n_25494;
wire newNet_350;
wire n_31608;
wire n_14187;
wire newNet_896;
wire n_9297;
wire n_30239;
wire newNet_1087;
wire n_33144;
wire n_3547;
wire n_21658;
wire n_38040;
wire FE_RN_1807_0;
wire n_27020;
wire n_19783;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_30_;
wire n_2029;
wire newNet_1587;
wire n_19250;
wire n_7721;
wire n_37754;
wire n_18787;
wire n_7102;
wire n_8845;
wire n_27803;
wire n_25296;
wire n_23752;
wire n_7365;
wire n_26442;
wire n_17878;
wire n_35692;
wire FE_OCP_RBN2592_n_25181;
wire n_39960;
wire n_43185;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_29_;
wire n_19058;
wire n_10265;
wire n_20676;
wire n_37698;
wire n_33298;
wire n_36440;
wire n_23567;
wire n_33146;
wire n_34115;
wire newNet_1776;
wire n_10284;
wire n_26660;
wire n_32406;
wire FE_RN_571_0;
wire n_22003;
wire n_16639;
wire n_36798;
wire n_37460;
wire n_31300;
wire n_1558;
wire n_12371;
wire n_3292;
wire n_32709;
wire newNet_962;
wire FE_OFN781_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire n_30801;
wire n_32944;
wire n_45132;
wire n_33689;
wire n_16592;
wire n_40651;
wire n_36613;
wire newNet_1906;
wire newNet_2190;
wire n_5989;
wire newNet_235;
wire n_16180;
wire n_43102;
wire newNet_10;
wire n_38680;
wire n_6217;
wire n_5782;
wire n_42237;
wire n_43744;
wire n_1090;
wire n_24682;
wire FE_OCP_DRV_N3148_n_33225;
wire newNet_1318;
wire n_6864;
wire n_37190;
wire newNet_2347;
wire n_35163;
wire n_15606;
wire n_31791;
wire n_30741;
wire n_4858;
wire n_29635;
wire FE_RN_1840_0;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_9_;
wire n_29118;
wire n_47233;
wire n_20633;
wire n_35725;
wire n_30124;
wire n_14477;
wire n_38722;
wire n_29996;
wire n_35251;
wire n_20731;
wire n_35438;
wire n_1505;
wire n_34664;
wire n_43635;
wire n_11258;
wire n_19857;
wire n_25342;
wire newNet_3619;
wire n_31735;
wire n_5870;
wire newNet_92;
wire FE_OCP_RBN2740_n_20565;
wire n_13028;
wire n_27236;
wire n_15244;
wire n_41023;
wire FE_RN_0_0;
wire n_4715;
wire n_28186;
wire n_9180;
wire n_18724;
wire n_21849;
wire n_27871;
wire n_36603;
wire n_21413;
wire n_14384;
wire n_23417;
wire n_44347;
wire n_2854;
wire n_7541;
wire n_4765;
wire n_19962;
wire n_43566;
wire n_20125;
wire n_17129;
wire n_4577;
wire n_36433;
wire n_22776;
wire newNet_3381;
wire n_28756;
wire newNet_2070;
wire n_3965;
wire n_22707;
wire n_30837;
wire n_10822;
wire n_27668;
wire n_27429;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_8_;
wire n_41388;
wire n_26467;
wire newNet_268;
wire n_14340;
wire n_42317;
wire n_9149;
wire n_25584;
wire n_40062;
wire newNet_2133;
wire n_36738;
wire n_4358;
wire n_17729;
wire n_6303;
wire n_31576;
wire newNet_2765;
wire FE_OCP_RBN3434_n_2224;
wire n_28887;
wire n_10859;
wire n_12126;
wire n_41306;
wire newNet_2711;
wire FE_OCPN939_n_7712;
wire n_31144;
wire n_8439;
wire n_28093;
wire n_34947;
wire n_780;
wire newNet_2294;
wire n_4399;
wire n_8773;
wire n_40475;
wire n_24527;
wire n_17732;
wire FE_OCP_RBN2001_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_34639;
wire n_27543;
wire n_32171;
wire n_12997;
wire n_43484;
wire FE_OFN822_n_4597;
wire n_28399;
wire n_13749;
wire n_14901;
wire FE_OCP_RBN2757_FE_RN_722_0;
wire n_30678;
wire n_38690;
wire n_2825;
wire n_23443;
wire n_44872;
wire n_41523;
wire n_33475;
wire n_3512;
wire newNet_1013;
wire n_2743;
wire n_13145;
wire FE_RN_553_0;
wire FE_OCP_RBN1133_n_16041;
wire n_14841;
wire n_19739;
wire n_4127;
wire n_15931;
wire newNet_3617;
wire mux_while_ln12_psv_q_1_;
wire n_46189;
wire n_30724;
wire n_24262;
wire n_26701;
wire n_5658;
wire n_1153;
wire n_23195;
wire newNet_3299;
wire newNet_3093;
wire FE_OCPN1755_n_16923;
wire FE_OCP_RBN1212_n_32142;
wire n_29520;
wire n_27621;
wire FE_OCP_RBN3629_n_38870;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_7_;
wire n_43036;
wire delay_xor_ln22_unr9_stage4_stallmux_q_21_;
wire n_1222;
wire n_1719;
wire n_12918;
wire n_39511;
wire n_40774;
wire n_14785;
wire n_36949;
wire FE_RN_1664_0;
wire FE_OCP_DRV_N1587_n_31012;
wire n_40806;
wire n_23488;
wire n_15736;
wire n_1399;
wire n_16886;
wire n_12105;
wire newNet_2554;
wire n_43785;
wire FE_OCP_RBN3833_n_19241;
wire n_22698;
wire newNet_3227;
wire n_28163;
wire newNet_691;
wire FE_OCP_RBN1375_n_20889;
wire n_34831;
wire n_4998;
wire n_13538;
wire n_31556;
wire n_31334;
wire n_31237;
wire n_12672;
wire n_303;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_7_;
wire n_42094;
wire FE_RN_134_0;
wire n_4780;
wire n_41155;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_28_;
wire n_42758;
wire FE_RN_1515_0;
wire FE_RN_674_0;
wire n_32752;
wire n_37402;
wire n_3838;
wire n_26617;
wire FE_RN_1740_0;
wire n_36013;
wire n_34311;
wire n_33718;
wire FE_OCP_RBN2473_n_8664;
wire n_6924;
wire n_46355;
wire n_38805;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_4_;
wire n_16267;
wire n_33617;
wire n_27056;
wire n_29363;
wire n_31355;
wire n_23832;
wire n_26439;
wire n_30204;
wire n_41722;
wire n_11370;
wire n_36555;
wire n_23609;
wire n_17128;
wire n_6848;
wire newNet_205;
wire n_2937;
wire n_35824;
wire n_44329;
wire FE_OCP_RBN3267_n_45224;
wire n_18212;
wire n_9816;
wire n_36332;
wire n_18036;
wire n_19036;
wire FE_RN_457_0;
wire n_8122;
wire n_35087;
wire n_38817;
wire n_25922;
wire newNet_3485;
wire n_30951;
wire n_9208;
wire n_28929;
wire n_34514;
wire n_5593;
wire n_40038;
wire n_26306;
wire n_7683;
wire delay_add_ln22_unr23_stage9_stallmux_q_16_;
wire n_26138;
wire FE_OCP_RBN2323_n_33942;
wire n_31065;
wire n_39495;
wire n_6958;
wire n_29609;
wire newNet_3549;
wire n_10408;
wire n_39602;
wire n_11847;
wire n_30212;
wire newNet_1117;
wire n_31773;
wire n_13120;
wire n_2420;
wire n_3912;
wire n_10302;
wire beta_26;
wire n_18090;
wire n_45205;
wire n_40260;
wire n_39679;
wire n_37596;
wire n_25037;
wire n_36467;
wire n_22938;
wire n_39466;
wire n_43849;
wire n_20407;
wire n_8609;
wire n_42021;
wire n_34477;
wire FE_OCP_RBN3665_n_4604;
wire n_34660;
wire FE_OCP_RBN2452_n_38537;
wire n_24521;
wire n_4332;
wire n_28269;
wire n_20164;
wire n_12332;
wire n_32617;
wire n_4593;
wire newNet_2637;
wire n_40395;
wire FE_RN_1369_0;
wire n_25146;
wire n_28371;
wire n_779;
wire FE_RN_238_0;
wire n_27271;
wire n_26321;
wire n_31640;
wire n_24781;
wire n_34805;
wire n_27452;
wire n_37593;
wire n_6669;
wire n_43649;
wire n_30718;
wire FE_OCP_RBN2417_n_24720;
wire n_181;
wire n_11758;
wire n_23281;
wire n_24399;
wire FE_RN_312_0;
wire n_38495;
wire FE_OCP_RBN3542_n_44575;
wire FE_OCP_RBN3219_n_21358;
wire FE_RN_111_0;
wire FE_OCP_DRV_N1596_n_21458;
wire n_20879;
wire n_7457;
wire n_20460;
wire n_22639;
wire n_35141;
wire n_9788;
wire n_2268;
wire n_29187;
wire n_22171;
wire n_39414;
wire n_20409;
wire n_42747;
wire sin_out_1;
wire n_19593;
wire n_30912;
wire FE_OCPN1519_n_31403;
wire n_8226;
wire n_31357;
wire n_36114;
wire newNet_202;
wire delay_xor_ln22_unr21_stage8_stallmux_q_8_;
wire n_45819;
wire n_22979;
wire n_32883;
wire n_10025;
wire n_18313;
wire n_7304;
wire n_7912;
wire n_38795;
wire n_24765;
wire n_3149;
wire FE_RN_293_0;
wire n_36583;
wire delay_xor_ln22_unr18_stage7_stallmux_q_8_;
wire n_28425;
wire n_27198;
wire n_12844;
wire n_5950;
wire n_9197;
wire n_26892;
wire n_33743;
wire n_37557;
wire n_16225;
wire n_37545;
wire n_2062;
wire n_11736;
wire n_18954;
wire n_32952;
wire n_482;
wire newNet_558;
wire n_25789;
wire n_10726;
wire n_43029;
wire n_12358;
wire FE_RN_1795_0;
wire n_8542;
wire FE_OCP_RBN2972_n_31239;
wire n_25478;
wire n_36872;
wire n_41947;
wire n_42574;
wire FE_RN_1275_0;
wire n_26498;
wire n_12480;
wire n_41702;
wire FE_RN_1056_0;
wire n_13490;
wire FE_RN_1841_0;
wire n_948;
wire n_18595;
wire newNet_3388;
wire n_2412;
wire n_33071;
wire n_36908;
wire n_3896;
wire n_5973;
wire n_40918;
wire n_31220;
wire n_10985;
wire n_12834;
wire n_11227;
wire n_18582;
wire n_22817;
wire FE_OCP_RBN3046_n_40231;
wire n_10158;
wire FE_OCP_RBN3073_n_43230;
wire n_33914;
wire newNet_2859;
wire n_4918;
wire n_12527;
wire n_28973;
wire n_14342;
wire n_31827;
wire n_8258;
wire newNet_1533;
wire n_20342;
wire n_39371;
wire n_37399;
wire n_33215;
wire n_15272;
wire n_1275;
wire FE_RN_9_0;
wire n_38253;
wire n_19968;
wire n_568;
wire n_35551;
wire newNet_30;
wire n_40213;
wire newNet_21;
wire n_2058;
wire n_8711;
wire newNet_823;
wire n_3888;
wire n_36920;
wire n_2921;
wire FE_RN_897_0;
wire n_32107;
wire n_43724;
wire FE_OCPN1012_n_41478;
wire n_42755;
wire n_31931;
wire n_29215;
wire n_26077;
wire delay_xor_ln22_unr3_stage2_stallmux_q_11_;
wire n_9893;
wire n_42926;
wire n_38083;
wire n_23851;
wire n_24454;
wire n_2557;
wire n_34868;
wire n_14377;
wire n_35363;
wire n_386;
wire n_10547;
wire n_33643;
wire FE_OCPN994_n_15552;
wire n_35340;
wire n_37383;
wire newNet_675;
wire newNet_326;
wire n_22733;
wire n_9434;
wire FE_RN_1402_0;
wire n_22750;
wire n_18285;
wire n_39283;
wire n_29982;
wire n_23157;
wire FE_OCPN977_n_31594;
wire n_5361;
wire n_23738;
wire FE_OCP_RBN3506_n_13860;
wire n_14225;
wire n_36364;
wire n_33235;
wire n_40018;
wire n_347;
wire n_39295;
wire n_40575;
wire n_27739;
wire n_34266;
wire n_7375;
wire FE_OCP_DRV_N1580_n_35482;
wire newNet_1434;
wire n_31150;
wire FE_OCP_RBN1056_n_18267;
wire n_24185;
wire n_1254;
wire n_10538;
wire n_12390;
wire n_22335;
wire n_32368;
wire n_22230;
wire n_17258;
wire n_18001;
wire n_30140;
wire newNet_3213;
wire n_19228;
wire n_43298;
wire newNet_1166;
wire n_32135;
wire n_1066;
wire n_36910;
wire FE_OCP_RBN2674_n_14991;
wire n_43342;
wire n_33957;
wire FE_OCP_RBN3060_FE_RN_640_0;
wire n_43313;
wire n_42606;
wire n_36304;
wire n_1769;
wire n_2928;
wire n_27951;
wire FE_OCP_RBN2297_n_2438;
wire n_27032;
wire n_17665;
wire n_27880;
wire n_30940;
wire n_7002;
wire n_33036;
wire n_24983;
wire n_32661;
wire n_35008;
wire n_39444;
wire n_27554;
wire n_17281;
wire newNet_1459;
wire n_26969;
wire n_8071;
wire n_9734;
wire n_33859;
wire n_31907;
wire n_25374;
wire newNet_3464;
wire n_13945;
wire n_5297;
wire n_12021;
wire FE_RN_1547_0;
wire n_37908;
wire n_30161;
wire n_2762;
wire n_4552;
wire n_19351;
wire n_39428;
wire n_35720;
wire newNet_1847;
wire newNet_1625;
wire delay_add_ln22_unr11_stage5_stallmux_q_0_;
wire n_13955;
wire n_33417;
wire n_198;
wire delay_sub_ln21_unr24_stage9_stallmux_q_6_;
wire FE_RN_1652_0;
wire n_31506;
wire n_26144;
wire n_26876;
wire n_18109;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_2_;
wire newNet_1513;
wire n_13530;
wire n_465;
wire n_27593;
wire n_31533;
wire FE_OCP_RBN2047_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire n_2050;
wire n_21881;
wire n_43091;
wire n_12345;
wire n_6885;
wire n_2182;
wire n_36418;
wire n_17819;
wire n_4022;
wire n_12791;
wire n_23067;
wire n_12621;
wire n_42914;
wire n_19953;
wire n_2959;
wire newNet_3350;
wire n_1601;
wire n_23932;
wire n_11593;
wire FE_OCPN1458_n_18426;
wire n_6562;
wire n_9582;
wire n_21872;
wire n_13431;
wire newNet_1637;
wire n_20155;
wire newNet_3535;
wire n_4400;
wire n_13685;
wire newNet_842;
wire n_36533;
wire newNet_471;
wire n_33347;
wire n_417;
wire n_15875;
wire n_35384;
wire n_7043;
wire n_11044;
wire FE_RN_1019_0;
wire n_649;
wire n_2123;
wire n_7713;
wire n_30100;
wire n_7740;
wire n_24576;
wire n_5690;
wire FE_OCP_RBN3461_n_7886;
wire FE_RN_1113_0;
wire n_27932;
wire n_8694;
wire n_1927;
wire n_40945;
wire n_34439;
wire n_11712;
wire n_15054;
wire n_14372;
wire n_33804;
wire n_33063;
wire newNet_2969;
wire n_12179;
wire n_43074;
wire n_30218;
wire n_8783;
wire FE_OFN738_n_22641;
wire FE_OCPN1026_n_25481;
wire n_8166;
wire n_22806;
wire newNet_2014;
wire FE_OCPN1480_n_23872;
wire n_45880;
wire FE_OCPN1422_n_35611;
wire n_6976;
wire n_19297;
wire n_6409;
wire n_10334;
wire n_1168;
wire n_28830;
wire n_21895;
wire delay_add_ln22_unr11_stage5_stallmux_q_20_;
wire n_17269;
wire n_36053;
wire n_2144;
wire n_4421;
wire n_39055;
wire n_32607;
wire n_12547;
wire n_28199;
wire newNet_3161;
wire n_13476;
wire newNet_3366;
wire n_8405;
wire n_36289;
wire n_35077;
wire n_13298;
wire n_32445;
wire n_3671;
wire n_37957;
wire n_5414;
wire n_8860;
wire n_31122;
wire n_7917;
wire n_36066;
wire n_40768;
wire FE_OCP_RBN2285_n_2433;
wire n_30093;
wire n_37954;
wire newNet_1826;
wire n_25221;
wire n_42931;
wire n_11190;
wire n_13270;
wire n_38015;
wire n_327;
wire newNet_2075;
wire n_7585;
wire n_41669;
wire n_9928;
wire n_15548;
wire n_4795;
wire n_11264;
wire n_6850;
wire FE_OCP_RBN2760_n_15180;
wire n_21831;
wire n_24315;
wire n_10104;
wire n_46148;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_12_;
wire newNet_1889;
wire n_15725;
wire n_33290;
wire n_33410;
wire n_35590;
wire delay_sub_ln23_0_unr21_stage8_stallmux_q;
wire n_26550;
wire n_20473;
wire n_5838;
wire n_43200;
wire FE_RN_148_0;
wire FE_OFN793_n_45813;
wire n_16347;
wire n_3400;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_13192;
wire n_10883;
wire n_40649;
wire n_37392;
wire n_14081;
wire n_12494;
wire n_24041;
wire n_13966;
wire n_27028;
wire FE_OCP_RBN3829_n_19204;
wire FE_RN_901_0;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_13_;
wire n_43397;
wire FE_OCPN1758_n_33213;
wire n_19014;
wire n_9136;
wire n_8943;
wire n_9150;
wire n_9317;
wire n_3749;
wire n_38706;
wire newNet_413;
wire n_39760;
wire n_16412;
wire n_37611;
wire n_42042;
wire n_36585;
wire newNet_818;
wire n_30247;
wire n_20665;
wire newNet_2774;
wire n_39702;
wire n_10570;
wire n_43869;
wire FE_OCP_DRV_N1568_n_19751;
wire n_18431;
wire n_43658;
wire n_4071;
wire n_32266;
wire newNet_1966;
wire n_9596;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_0_;
wire n_30471;
wire n_11363;
wire n_36748;
wire n_6630;
wire FE_RN_1032_0;
wire n_35910;
wire n_4462;
wire n_24566;
wire n_34464;
wire n_15136;
wire n_395;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_17_;
wire n_11138;
wire n_46977;
wire n_34369;
wire n_30015;
wire n_8572;
wire n_10503;
wire FE_OCP_RBN2695_n_14814;
wire n_30036;
wire n_5231;
wire n_30885;
wire n_22021;
wire n_4790;
wire n_30608;
wire n_33003;
wire FE_OCP_RBN1175_n_18981;
wire n_23665;
wire n_46212;
wire n_33305;
wire n_42700;
wire FE_OCP_DRV_N1592_n_34327;
wire n_45066;
wire newNet_3601;
wire newNet_279;
wire n_3113;
wire n_10724;
wire n_34535;
wire n_11080;
wire n_39368;
wire n_1484;
wire FE_RN_50_0;
wire n_9910;
wire newNet_2362;
wire n_20595;
wire n_10417;
wire n_13514;
wire n_30696;
wire n_29652;
wire n_42349;
wire n_39528;
wire newNet_2756;
wire n_29123;
wire n_40696;
wire delay_add_ln22_unr11_stage5_stallmux_q_26_;
wire n_4958;
wire delay_xor_ln21_unr9_stage4_stallmux_q_7_;
wire n_24127;
wire newNet_3178;
wire n_25133;
wire newNet_3588;
wire FE_RN_1349_0;
wire n_33170;
wire n_11967;
wire n_1510;
wire n_561;
wire n_33994;
wire FE_OCPN1472_n_13434;
wire newNet_1562;
wire FE_RN_1209_0;
wire n_39402;
wire n_20107;
wire n_5904;
wire n_33169;
wire n_39974;
wire n_37850;
wire n_16842;
wire newNet_1388;
wire n_26332;
wire n_19355;
wire n_7801;
wire n_26070;
wire n_9771;
wire n_31027;
wire n_29399;
wire n_7849;
wire n_35273;
wire n_36646;
wire n_25258;
wire n_41484;
wire n_19283;
wire n_29010;
wire newNet_3675;
wire delay_add_ln22_unr8_stage4_stallmux_q_12_;
wire n_32711;
wire n_7095;
wire n_12701;
wire n_24536;
wire newNet_3390;
wire n_14242;
wire n_11830;
wire n_13260;
wire n_27703;
wire newNet_2850;
wire n_2046;
wire n_10760;
wire n_38431;
wire FE_OCPN3774_n_14730;
wire n_9169;
wire FE_OCP_RBN1193_n_22542;
wire n_40006;
wire n_33085;
wire n_31038;
wire n_5089;
wire n_34081;
wire newNet_368;
wire n_11789;
wire FE_RN_1749_0;
wire FE_OCP_RBN2951_n_21489;
wire n_17185;
wire n_27827;
wire n_36198;
wire newNet_2128;
wire n_27129;
wire n_34069;
wire n_11056;
wire FE_OCP_RBN2384_n_8342;
wire n_16263;
wire n_8375;
wire n_15708;
wire n_13238;
wire n_43695;
wire n_23471;
wire n_12502;
wire n_11364;
wire n_6688;
wire n_32281;
wire FE_OCPN1386_n_470;
wire n_7767;
wire n_9086;
wire n_30564;
wire n_34292;
wire newNet_3623;
wire n_5526;
wire n_36596;
wire n_40824;
wire n_36213;
wire newNet_236;
wire n_23843;
wire n_6466;
wire n_15781;
wire n_6102;
wire n_29932;
wire n_5616;
wire n_26596;
wire newNet_1543;
wire newNet_901;
wire n_31270;
wire n_1207;
wire n_14469;
wire newNet_245;
wire FE_OCP_RBN2214_FE_OCPN950_n_28595;
wire n_32437;
wire n_2656;
wire n_13138;
wire n_39220;
wire n_11983;
wire n_13462;
wire n_45721;
wire n_764;
wire n_36723;
wire n_22730;
wire FE_OCP_RBN1839_n_19528;
wire FE_OCP_RBN2314_n_41420;
wire newNet_2421;
wire n_6871;
wire n_12154;
wire n_14269;
wire n_20254;
wire n_36348;
wire n_29873;
wire newNet_2084;
wire n_17689;
wire n_6008;
wire n_15429;
wire n_31955;
wire n_43538;
wire n_7930;
wire n_8532;
wire n_10923;
wire FE_RN_168_0;
wire n_28604;
wire newNet_1121;
wire n_9884;
wire n_39324;
wire FE_OCP_RBN1837_FE_RN_1542_0;
wire n_24094;
wire n_13756;
wire n_40206;
wire n_44955;
wire n_18473;
wire n_15805;
wire n_31863;
wire FE_RN_1297_0;
wire n_279;
wire n_27519;
wire n_1023;
wire FE_RN_283_0;
wire n_25947;
wire n_30863;
wire n_17541;
wire n_4585;
wire n_40270;
wire FE_RN_1126_0;
wire FE_OCP_RBN3214_n_44365;
wire n_23309;
wire n_32685;
wire n_10631;
wire n_7443;
wire n_46380;
wire FE_OCP_RBN3075_FE_OFN807_n_46195;
wire n_35180;
wire n_25937;
wire n_25311;
wire n_38888;
wire n_22431;
wire n_23354;
wire FE_OCP_RBN3058_n_36515;
wire n_34442;
wire newNet_3289;
wire n_4197;
wire n_23348;
wire n_21128;
wire newNet_3304;
wire n_19649;
wire n_20659;
wire n_31567;
wire newNet_1418;
wire n_24199;
wire n_39100;
wire n_19315;
wire n_43702;
wire n_25510;
wire n_20127;
wire n_18480;
wire n_30022;
wire FE_OCP_RBN3130_n_17591;
wire n_35964;
wire n_39730;
wire n_18812;
wire n_27443;
wire delay_add_ln22_unr11_stage5_stallmux_q_5_;
wire FE_OCPN1239_n_37945;
wire n_536;
wire n_31664;
wire n_33393;
wire n_3771;
wire n_39005;
wire n_37371;
wire FE_OCP_RBN3670_n_46982;
wire n_43040;
wire n_15636;
wire n_7166;
wire FE_OCP_DRV_N1608_n_31473;
wire n_5197;
wire n_1644;
wire n_36874;
wire n_34379;
wire n_26624;
wire n_2772;
wire FE_RN_1085_0;
wire n_16972;
wire n_16895;
wire n_7783;
wire n_3490;
wire n_22980;
wire n_38062;
wire FE_OCP_RBN2119_n_45224;
wire n_11390;
wire n_30281;
wire n_32353;
wire n_27949;
wire n_23109;
wire n_40878;
wire newNet_683;
wire n_32774;
wire n_31082;
wire FE_OCP_RBN1844_n_20910;
wire n_40135;
wire n_9293;
wire n_37734;
wire n_16254;
wire n_41954;
wire n_6876;
wire n_36950;
wire n_3371;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_1_;
wire n_23320;
wire n_5876;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_10_;
wire n_23101;
wire n_37209;
wire n_12776;
wire n_11993;
wire n_38719;
wire n_33975;
wire n_33888;
wire n_34355;
wire n_33515;
wire n_10746;
wire n_14874;
wire n_22719;
wire n_10598;
wire n_37753;
wire n_24155;
wire n_44037;
wire n_216;
wire FE_RN_1845_0;
wire n_1961;
wire FE_RN_683_0;
wire n_1535;
wire n_20145;
wire n_20374;
wire n_18875;
wire n_33690;
wire n_37680;
wire n_13590;
wire n_1663;
wire FE_OCP_RBN3848_FE_RN_1548_0;
wire n_26988;
wire n_9288;
wire n_10368;
wire n_10468;
wire FE_RN_440_0;
wire n_23303;
wire n_13336;
wire FE_OCP_DRV_N3156_n_15342;
wire n_39131;
wire n_2846;
wire n_38747;
wire n_8064;
wire n_9324;
wire n_9381;
wire n_3469;
wire n_42475;
wire newNet_2569;
wire n_2113;
wire n_38685;
wire n_2364;
wire FE_RN_7_0;
wire FE_OCP_RBN3124_n_6557;
wire n_16041;
wire n_1351;
wire n_27187;
wire n_26160;
wire n_19454;
wire n_21439;
wire FE_RN_1809_0;
wire n_32595;
wire FE_OCP_RBN2903_n_44174;
wire newNet_1768;
wire n_40144;
wire n_16366;
wire n_16046;
wire cos_out_20;
wire n_554;
wire n_28226;
wire n_14781;
wire newNet_2662;
wire n_21558;
wire n_22225;
wire newNet_1095;
wire n_26346;
wire n_7536;
wire n_13489;
wire n_34307;
wire newNet_2844;
wire n_3811;
wire FE_OCP_RBN3737_n_12027;
wire n_2190;
wire n_2170;
wire n_29327;
wire newNet_2561;
wire n_29902;
wire FE_RN_122_0;
wire n_39021;
wire n_38296;
wire n_37605;
wire n_43232;
wire n_15141;
wire n_757;
wire n_38522;
wire n_34694;
wire n_30432;
wire n_11896;
wire n_831;
wire n_14659;
wire n_31813;
wire n_12202;
wire n_30138;
wire newNet_3375;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_3_;
wire FE_OCP_RBN3586_n_25295;
wire n_16566;
wire n_32927;
wire n_30635;
wire n_19476;
wire n_26021;
wire n_34245;
wire n_22860;
wire n_46233;
wire n_18548;
wire FE_RN_919_0;
wire n_41062;
wire FE_RN_155_0;
wire n_6351;
wire n_19164;
wire newNet_977;
wire n_34609;
wire n_29444;
wire n_12921;
wire n_31439;
wire n_17909;
wire n_35118;
wire n_45532;
wire n_20021;
wire newNet_1151;
wire n_8934;
wire n_26019;
wire n_10775;
wire newNet_447;
wire n_5713;
wire FE_OCPN991_n_22249;
wire FE_OCP_RBN3518_n_8498;
wire n_2835;
wire n_9654;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_23_;
wire n_43758;
wire n_32641;
wire n_1017;
wire n_16004;
wire n_30254;
wire n_844;
wire FE_OCPN1028_n_4182;
wire n_22300;
wire n_40258;
wire n_10710;
wire FE_OCPN969_n_19342;
wire n_10629;
wire n_3733;
wire n_40848;
wire n_16942;
wire n_7591;
wire n_4155;
wire n_43136;
wire n_1694;
wire n_39272;
wire n_13178;
wire newNet_1240;
wire FE_OCPN1522_n_26054;
wire n_27940;
wire n_38755;
wire n_21247;
wire n_3530;
wire n_9110;
wire n_15528;
wire n_40998;
wire n_6833;
wire n_21309;
wire FE_OCP_RBN3112_n_32254;
wire n_25713;
wire FE_RN_426_0;
wire n_47017;
wire n_29438;
wire n_2875;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_22_;
wire n_20011;
wire n_504;
wire n_8059;
wire n_45891;
wire FE_OCP_RBN2576_n_47017;
wire n_17930;
wire n_31989;
wire n_26810;
wire n_33402;
wire n_24336;
wire n_33863;
wire n_29878;
wire n_21772;
wire n_26267;
wire FE_RN_1779_0;
wire n_36579;
wire n_31048;
wire n_8217;
wire newNet_3109;
wire n_5181;
wire n_19442;
wire n_12147;
wire n_17432;
wire n_1935;
wire n_29781;
wire n_23407;
wire n_43514;
wire n_17391;
wire FE_RN_1140_0;
wire n_36480;
wire n_16469;
wire n_26694;
wire n_27815;
wire n_47252;
wire n_38843;
wire n_44718;
wire n_9359;
wire n_29380;
wire n_25095;
wire n_35515;
wire n_41196;
wire n_22280;
wire delay_xor_ln21_unr3_stage2_stallmux_q_5_;
wire n_4309;
wire n_38597;
wire n_43770;
wire n_23943;
wire FE_RN_794_0;
wire newNet_3495;
wire n_32278;
wire newNet_500;
wire n_39922;
wire n_32403;
wire n_33106;
wire n_22330;
wire n_39370;
wire n_26032;
wire n_41458;
wire n_17743;
wire FE_RN_1772_0;
wire n_3532;
wire n_38414;
wire n_1581;
wire n_39838;
wire n_29239;
wire n_21094;
wire n_41934;
wire newNet_987;
wire n_27723;
wire n_66;
wire n_27043;
wire FE_OCPN1752_n_29420;
wire n_35127;
wire n_16037;
wire n_37516;
wire n_25244;
wire n_21023;
wire newNet_2093;
wire newNet_3435;
wire n_12717;
wire n_6899;
wire newNet_1183;
wire n_27142;
wire n_14455;
wire n_35071;
wire newNet_2901;
wire n_8415;
wire n_12412;
wire n_2445;
wire FE_OCP_RBN3639_n_44490;
wire FE_RN_1761_0;
wire newNet_300;
wire FE_RN_766_0;
wire n_25669;
wire newNet_2233;
wire n_25275;
wire n_13583;
wire n_14280;
wire n_9535;
wire n_29203;
wire n_37013;
wire n_5109;
wire n_16820;
wire n_11305;
wire n_34362;
wire n_40435;
wire n_238;
wire n_791;
wire FE_RN_1430_0;
wire n_15328;
wire n_12381;
wire n_37834;
wire n_18455;
wire delay_xor_ln22_unr6_stage3_stallmux_q_10_;
wire n_42055;
wire n_18065;
wire n_42726;
wire n_16545;
wire n_33917;
wire n_9318;
wire n_37469;
wire n_44434;
wire newNet_3222;
wire n_40050;
wire n_660;
wire n_43472;
wire n_24820;
wire newNet_642;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_2_;
wire n_1287;
wire n_37867;
wire n_32876;
wire newNet_3734;
wire n_1879;
wire newNet_3448;
wire n_40668;
wire newNet_3047;
wire n_12588;
wire n_5185;
wire n_14750;
wire n_18245;
wire n_25024;
wire FE_RN_1267_0;
wire n_24722;
wire n_20088;
wire newNet_3341;
wire FE_OCP_RBN1842_n_20910;
wire newNet_1375;
wire n_38169;
wire newNet_2251;
wire n_5929;
wire newNet_1527;
wire n_3215;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_5_;
wire n_18187;
wire n_12699;
wire delay_add_ln22_unr27_stage10_stallmux_q_17_;
wire n_23914;
wire newNet_512;
wire n_45146;
wire n_19498;
wire n_9901;
wire n_19802;
wire n_10803;
wire n_21531;
wire n_19108;
wire n_37008;
wire n_32216;
wire n_27326;
wire n_25280;
wire n_19249;
wire n_5000;
wire n_15574;
wire newNet_1027;
wire n_2596;
wire n_33092;
wire n_33314;
wire n_42837;
wire delay_xor_ln22_unr3_stage2_stallmux_q_18_;
wire n_25519;
wire n_13846;
wire n_33557;
wire n_15335;
wire FE_OCP_RBN3331_n_44962;
wire newNet_3327;
wire n_15402;
wire n_45506;
wire n_6078;
wire newNet_3407;
wire n_10063;
wire n_10667;
wire n_29353;
wire n_7222;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_13_;
wire newNet_1079;
wire n_6194;
wire FE_OCPN3791_n_36069;
wire n_29969;
wire n_38555;
wire n_22970;
wire n_28095;
wire FE_OCP_RBN3817_n_44061;
wire n_8941;
wire n_9241;
wire n_26225;
wire n_36026;
wire n_31182;
wire newNet_745;
wire n_4828;
wire newNet_1952;
wire n_12165;
wire n_18508;
wire newNet_2990;
wire n_18866;
wire FE_OCPN3775_n_14730;
wire n_36768;
wire newNet_3665;
wire n_21140;
wire n_37184;
wire FE_OCP_RBN2166_n_32892;
wire n_30392;
wire n_11331;
wire newNet_2435;
wire n_35047;
wire FE_OCP_RBN3080_n_16977;
wire n_34772;
wire newNet_2781;
wire n_616;
wire FE_OCP_RBN3489_n_3390;
wire n_33026;
wire newNet_1137;
wire n_20519;
wire n_37626;
wire n_1591;
wire newNet_653;
wire n_40628;
wire n_13909;
wire delay_add_ln22_unr20_stage8_stallmux_q_6_;
wire n_29156;
wire n_22596;
wire n_22630;
wire n_35732;
wire n_19053;
wire n_29806;
wire FE_OCPN956_n_39096;
wire n_7245;
wire n_977;
wire FE_RN_1484_0;
wire n_38723;
wire n_30250;
wire n_16601;
wire n_23743;
wire FE_OCPN1461_n_23759;
wire n_22687;
wire FE_OCP_RBN2371_n_8221;
wire n_38244;
wire n_38656;
wire n_37259;
wire n_35288;
wire n_38893;
wire n_26058;
wire n_31561;
wire n_23678;
wire n_40867;
wire FE_RN_1776_0;
wire n_42221;
wire n_17164;
wire n_15557;
wire n_17221;
wire n_37121;
wire n_22395;
wire n_12744;
wire FE_RN_914_0;
wire n_14602;
wire n_44040;
wire n_11302;
wire delay_xor_ln22_unr12_stage5_stallmux_q_7_;
wire n_391;
wire delay_add_ln22_unr5_stage3_stallmux_q_18_;
wire n_16744;
wire n_30592;
wire n_36805;
wire n_23807;
wire n_17755;
wire n_5035;
wire n_435;
wire n_4012;
wire n_29250;
wire n_9825;
wire n_12325;
wire delay_xor_ln21_unr9_stage4_stallmux_q_22_;
wire n_22788;
wire n_39773;
wire n_2063;
wire n_41477;
wire FE_OCP_DRV_N1600_n_21493;
wire n_34198;
wire n_47244;
wire n_15363;
wire n_28837;
wire n_2725;
wire n_36688;
wire n_3593;
wire n_26523;
wire n_18975;
wire n_22473;
wire n_15672;
wire n_4238;
wire n_21905;
wire newNet_1075;
wire FE_RN_890_0;
wire n_8306;
wire n_24962;
wire n_36489;
wire n_41215;
wire FE_OCPN1257_n_13831;
wire newNet_914;
wire n_39120;
wire n_7738;
wire n_23334;
wire n_3737;
wire n_25660;
wire n_16017;
wire n_11351;
wire n_26131;
wire newNet_3085;
wire n_26861;
wire n_14149;
wire n_30113;
wire n_234;
wire n_38335;
wire n_27755;
wire n_14759;
wire n_11345;
wire n_34788;
wire n_20527;
wire n_42790;
wire n_31895;
wire newNet_474;
wire n_10115;
wire n_6030;
wire n_36947;
wire newNet_121;
wire FE_RN_555_0;
wire n_15091;
wire newNet_2146;
wire n_14997;
wire FE_RN_956_0;
wire newNet_1536;
wire delay_xor_ln21_unr15_stage6_stallmux_q_11_;
wire n_37502;
wire FE_OCP_RBN2324_n_13616;
wire delay_add_ln22_unr17_stage7_stallmux_q_21_;
wire newNet_392;
wire n_20743;
wire n_18323;
wire n_34135;
wire n_24615;
wire FE_OCP_RBN1173_n_13858;
wire n_21018;
wire n_731;
wire n_1270;
wire n_23760;
wire n_11922;
wire newNet_1329;
wire n_36108;
wire n_12685;
wire n_15974;
wire n_14463;
wire n_8819;
wire n_30064;
wire n_15763;
wire n_39207;
wire n_27655;
wire n_5980;
wire n_16536;
wire n_29975;
wire n_29318;
wire newNet_2316;
wire n_18079;
wire FE_RN_990_0;
wire FE_OCPN3749_n_34296;
wire n_21461;
wire n_34283;
wire FE_OCPN3761_n_2466;
wire n_14358;
wire n_33905;
wire FE_RN_1571_0;
wire delay_xor_ln21_unr18_stage7_stallmux_q_6_;
wire n_1996;
wire n_5805;
wire n_20980;
wire FE_OCP_RBN2527_n_3421;
wire n_37854;
wire n_37874;
wire n_10430;
wire n_42264;
wire n_7548;
wire n_25542;
wire n_27361;
wire n_7813;
wire n_20885;
wire newNet_2068;
wire n_15559;
wire FE_RN_195_0;
wire n_22154;
wire n_21074;
wire n_16706;
wire n_42483;
wire n_41856;
wire n_21645;
wire n_8236;
wire n_40829;
wire n_7598;
wire n_19712;
wire newNet_2811;
wire n_33921;
wire FE_OCP_RBN2435_n_14072;
wire n_5240;
wire n_10089;
wire n_31609;
wire FE_RN_621_0;
wire n_26271;
wire n_9665;
wire n_15187;
wire FE_OCPN1490_n_30823;
wire n_46223;
wire FE_OCP_RBN2715_n_14982;
wire n_25923;
wire FE_OCP_DRV_N1544_n_18854;
wire n_18533;
wire n_10369;
wire n_5544;
wire newNet_17;
wire n_18854;
wire n_31745;
wire n_23452;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_20_;
wire n_26195;
wire n_18400;
wire newNet_2490;
wire n_4105;
wire n_36387;
wire n_37424;
wire n_15417;
wire n_25534;
wire n_11085;
wire n_20929;
wire n_45026;
wire delay_add_ln22_unr27_stage10_stallmux_q_6_;
wire n_138;
wire n_8004;
wire FE_OCPN1436_n_19855;
wire n_2507;
wire n_9475;
wire n_13095;
wire newNet_1612;
wire n_6124;
wire n_10702;
wire FE_OCPN1736_n_37877;
wire n_28742;
wire n_12251;
wire FE_RN_667_0;
wire n_30588;
wire n_14633;
wire n_24370;
wire n_39757;
wire n_330;
wire n_16663;
wire n_11883;
wire n_30812;
wire n_40864;
wire n_34075;
wire FE_OCP_RBN3438_n_33750;
wire n_14306;
wire n_14514;
wire newNet_2298;
wire n_20924;
wire n_29384;
wire n_40757;
wire n_21826;
wire n_2427;
wire n_14906;
wire n_16076;
wire newNet_1752;
wire newNet_1282;
wire n_3867;
wire n_44826;
wire n_209;
wire n_42;
wire newNet_1235;
wire n_2683;
wire n_8423;
wire n_27439;
wire newNet_1352;
wire n_4025;
wire delay_add_ln22_unr23_stage9_stallmux_q_17_;
wire n_1760;
wire n_20872;
wire n_41596;
wire n_38985;
wire newNet_1798;
wire n_25454;
wire newNet_2398;
wire n_9644;
wire n_3626;
wire n_32441;
wire n_36562;
wire FE_RN_1716_0;
wire n_36256;
wire n_37563;
wire FE_OCPN1462_n_23759;
wire n_34577;
wire n_6816;
wire n_19130;
wire n_5517;
wire delay_xor_ln22_unr3_stage2_stallmux_q_10_;
wire n_25745;
wire n_29573;
wire FE_OCP_RBN2269_n_33803;
wire n_15163;
wire n_43905;
wire n_5125;
wire n_28204;
wire n_20042;
wire n_4466;
wire n_39105;
wire n_40245;
wire n_29174;
wire n_25578;
wire n_6412;
wire n_43282;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_12_;
wire n_44059;
wire n_23717;
wire n_36654;
wire n_11813;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_14_;
wire n_15422;
wire n_20967;
wire newNet_1723;
wire n_35442;
wire n_41500;
wire n_10445;
wire n_11601;
wire n_39822;
wire n_34938;
wire newNet_646;
wire newNet_605;
wire n_16624;
wire n_18023;
wire n_27161;
wire n_36261;
wire n_42957;
wire n_10399;
wire n_22700;
wire newNet_2886;
wire n_4911;
wire n_24210;
wire n_17050;
wire n_4212;
wire n_10970;
wire FE_RN_1337_0;
wire FE_OCP_RBN2451_n_34278;
wire n_34988;
wire n_41149;
wire n_26875;
wire n_38114;
wire FE_RN_482_0;
wire n_21633;
wire delay_add_ln22_unr23_stage9_stallmux_q_31_;
wire newNet_3018;
wire n_36290;
wire n_22288;
wire n_28405;
wire n_9057;
wire n_570;
wire FE_RN_332_0;
wire n_31787;
wire n_47251;
wire n_6646;
wire n_43128;
wire n_41786;
wire n_45808;
wire n_6986;
wire n_36867;
wire n_20285;
wire n_15541;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_15_;
wire n_13055;
wire n_25501;
wire n_28660;
wire FE_OCP_RBN2975_n_5531;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_16_;
wire newNet_2737;
wire n_30925;
wire n_20416;
wire n_4226;
wire FE_OCP_RBN3077_FE_OFN807_n_46195;
wire n_15989;
wire n_25176;
wire n_5504;
wire FE_RN_594_0;
wire n_42685;
wire n_46254;
wire FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire n_38436;
wire n_39350;
wire FE_OCP_RBN1060_n_24473;
wire newNet_1853;
wire n_31652;
wire n_39987;
wire n_6998;
wire n_14803;
wire n_20072;
wire n_10957;
wire FE_OCPN962_n_28506;
wire FE_RN_311_0;
wire n_24225;
wire FE_OCP_RBN2571_n_29922;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_25_;
wire n_21535;
wire n_6248;
wire n_2391;
wire n_19198;
wire n_12573;
wire n_42626;
wire n_26842;
wire FE_OCPN1228_n_46101;
wire n_17518;
wire n_7059;
wire n_23778;
wire newNet_638;
wire n_42435;
wire n_9527;
wire newNet_2450;
wire n_1630;
wire n_31418;
wire n_14265;
wire FE_OCP_RBN3313_delay_xor_ln22_unr18_stage7_stallmux_q_2_;
wire FE_RN_895_0;
wire n_5884;
wire n_26998;
wire newNet_3722;
wire n_15460;
wire n_18382;
wire n_7833;
wire FE_OCPN3777_n_43019;
wire n_15581;
wire n_8907;
wire n_44859;
wire n_22449;
wire FE_RN_1628_0;
wire FE_RN_164_0;
wire n_7259;
wire n_26643;
wire n_18589;
wire n_15009;
wire newNet_1461;
wire newNet_3513;
wire newNet_1668;
wire n_17619;
wire newNet_1313;
wire n_40002;
wire n_8492;
wire n_26675;
wire n_14056;
wire n_29113;
wire newNet_1263;
wire n_30454;
wire n_37213;
wire n_17638;
wire newNet_486;
wire n_28314;
wire n_30323;
wire n_28222;
wire delay_xor_ln22_unr18_stage7_stallmux_q_10_;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_11_;
wire n_2613;
wire newNet_3424;
wire newNet_1898;
wire n_20802;
wire n_874;
wire n_20704;
wire n_18163;
wire FE_RN_1470_0;
wire n_15623;
wire n_18265;
wire n_28572;
wire FE_OCP_RBN3703_n_26231;
wire newNet_997;
wire n_10091;
wire newNet_978;
wire n_42989;
wire n_33183;
wire n_41707;
wire newNet_1006;
wire n_7698;
wire n_11277;
wire FE_RN_189_0;
wire n_24665;
wire n_6364;
wire n_1608;
wire n_37785;
wire n_21776;
wire n_21326;
wire n_3333;
wire n_3025;
wire n_33603;
wire n_26823;
wire n_6658;
wire n_8728;
wire n_11236;
wire delay_xor_ln21_unr28_stage10_stallmux_q_1_;
wire n_6968;
wire n_3394;
wire n_23313;
wire n_24031;
wire newNet_2656;
wire n_26103;
wire n_8024;
wire n_36173;
wire n_7558;
wire n_46170;
wire n_34419;
wire n_28908;
wire newNet_551;
wire n_17523;
wire n_30977;
wire n_29565;
wire n_16192;
wire n_36642;
wire FE_OCP_RBN2869_n_10480;
wire n_6389;
wire newNet_1595;
wire newNet_795;
wire n_20535;
wire n_43393;
wire FE_OCP_DRV_N3155_n_15342;
wire n_27609;
wire newNet_85;
wire n_20947;
wire n_43406;
wire n_31426;
wire n_11919;
wire n_2164;
wire n_15042;
wire n_4789;
wire n_18295;
wire n_35892;
wire n_1231;
wire n_33945;
wire n_23033;
wire n_8488;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_29_;
wire n_28914;
wire FE_OCP_RBN3266_n_45224;
wire n_22229;
wire FE_OCPN1737_n_19052;
wire n_1539;
wire n_38481;
wire n_28156;
wire FE_RN_936_0;
wire n_24891;
wire n_10755;
wire n_27551;
wire n_10905;
wire FE_OCPN1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_18375;
wire newNet_2920;
wire n_27292;
wire newNet_2864;
wire n_18713;
wire n_27673;
wire n_24106;
wire n_155;
wire n_5405;
wire n_18317;
wire n_25720;
wire FE_RN_1497_0;
wire FE_OCPN3748_n_34296;
wire n_15855;
wire n_32808;
wire n_7198;
wire delay_xor_ln21_unr15_stage6_stallmux_q_2_;
wire n_26918;
wire n_35917;
wire newNet_2955;
wire FE_OCP_RBN3634_n_47260;
wire n_14096;
wire newNet_2648;
wire n_1799;
wire FE_OCP_RBN1195_n_22542;
wire n_33697;
wire n_11680;
wire n_8791;
wire n_31544;
wire n_30709;
wire n_943;
wire n_37435;
wire n_42192;
wire n_31635;
wire n_38130;
wire FE_OCP_RBN2300_n_7817;
wire FE_OCP_RBN2183_FE_RN_464_0;
wire n_14011;
wire n_20478;
wire newNet_2400;
wire n_532;
wire n_8670;
wire n_40953;
wire newNet_168;
wire newNet_2933;
wire n_29312;
wire n_37284;
wire FE_OCP_DRV_N3741_n_29576;
wire n_36616;
wire delay_add_ln22_unr20_stage8_stallmux_q_15_;
wire n_6155;
wire n_42564;
wire n_43061;
wire FE_RN_1695_0;
wire n_18494;
wire n_42140;
wire n_4296;
wire n_15832;
wire n_40845;
wire n_43687;
wire n_46934;
wire n_33313;
wire n_28531;
wire n_20085;
wire FE_OCPN1402_n_9642;
wire n_36405;
wire n_32745;
wire delay_sub_ln21_unr24_stage9_stallmux_q_2_;
wire n_2299;
wire n_41631;
wire n_38463;
wire newNet_2117;
wire n_31708;
wire delay_add_ln22_unr14_stage6_stallmux_q_26_;
wire n_13775;
wire n_37757;
wire newNet_2821;
wire n_39557;
wire n_44887;
wire n_28962;
wire n_20190;
wire n_3843;
wire n_40517;
wire n_19219;
wire n_39009;
wire FE_OCP_RBN3338_n_44610;
wire n_42581;
wire n_36130;
wire n_23856;
wire n_27958;
wire n_1444;
wire n_27223;
wire FE_OCP_RBN3503_n_38592;
wire n_16834;
wire n_9388;
wire n_33450;
wire n_6720;
wire n_30303;
wire n_37262;
wire FE_RN_291_0;
wire n_39242;
wire n_17207;
wire newNet_3155;
wire n_1843;
wire n_7238;
wire n_38180;
wire n_27241;
wire n_39690;
wire n_36165;
wire n_16375;
wire n_37299;
wire n_41869;
wire newNet_2277;
wire n_41164;
wire n_26547;
wire n_21124;
wire n_18730;
wire n_30736;
wire n_38038;
wire n_14865;
wire n_999;
wire n_29765;
wire n_32576;
wire n_5831;
wire n_9958;
wire n_35309;
wire n_23823;
wire n_28522;
wire n_17313;
wire n_30166;
wire n_37197;
wire n_6743;
wire n_37483;
wire n_35470;
wire n_1243;
wire n_29504;
wire n_13739;
wire n_35684;
wire n_19638;
wire n_12207;
wire n_45149;
wire n_31361;
wire n_4100;
wire n_21621;
wire n_19567;
wire newNet_905;
wire n_30759;
wire n_6106;
wire n_31978;
wire n_14882;
wire n_18829;
wire n_34563;
wire n_22903;
wire FE_OCP_RBN2510_n_13896;
wire newNet_1086;
wire newNet_2707;
wire newNet_63;
wire n_43720;
wire n_35665;
wire n_7386;
wire n_42299;
wire n_14352;
wire n_41590;
wire n_7722;
wire n_33519;
wire n_15921;
wire n_46386;
wire n_7312;
wire n_8800;
wire n_652;
wire n_10784;
wire n_36712;
wire n_32781;
wire n_33288;
wire n_22487;
wire newNet_1590;
wire n_7529;
wire n_45497;
wire n_35886;
wire n_20378;
wire newNet_3608;
wire n_41511;
wire FE_RN_1821_0;
wire n_15031;
wire n_3098;
wire n_41140;
wire n_33143;
wire n_12055;
wire n_27894;
wire n_20445;
wire n_39841;
wire n_41112;
wire n_27309;
wire n_40422;
wire n_16392;
wire newNet_1871;
wire newNet_2426;
wire n_24853;
wire n_2645;
wire n_20714;
wire n_8313;
wire n_30229;
wire n_27097;
wire n_32701;
wire n_32530;
wire n_23794;
wire n_10322;
wire n_45153;
wire newNet_2690;
wire n_40704;
wire n_7866;
wire n_26400;
wire FE_RN_353_0;
wire n_34168;
wire n_1387;
wire delay_sub_ln21_0_unr23_stage9_stallmux_q_16_;
wire n_38456;
wire n_33776;
wire n_19927;
wire n_21709;
wire n_12117;
wire n_42715;
wire FE_RN_8_0;
wire n_7401;
wire n_26003;
wire newNet_2387;
wire n_42768;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_2_;
wire n_26788;
wire n_11578;
wire FE_OCP_RBN2828_n_30731;
wire n_32810;
wire n_31199;
wire FE_RN_1520_0;
wire n_18477;
wire n_1145;
wire n_30055;
wire n_13593;
wire n_47021;
wire n_3699;
wire n_24958;
wire n_27175;
wire n_43328;
wire n_37444;
wire n_18916;
wire n_11746;
wire FE_RN_1412_0;
wire delay_add_ln22_unr17_stage7_stallmux_q_25_;
wire n_37492;
wire n_23204;
wire n_43790;
wire n_24882;
wire n_23660;
wire n_28505;
wire n_1260;
wire n_39069;
wire newNet_3655;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_5_;
wire newNet_1733;
wire n_43802;
wire FE_OCP_RBN2112_n_22650;
wire FE_OCP_RBN2697_n_14814;
wire n_34759;
wire FE_OCP_RBN1927_cordic_combinational_sub_ln23_0_unr12_z_0__;
wire n_35517;
wire n_40469;
wire n_32358;
wire n_23022;
wire newNet_2389;
wire n_24131;
wire FE_RN_652_0;
wire n_16128;
wire n_2269;
wire n_7159;
wire n_10690;
wire n_32288;
wire n_29136;
wire n_6910;
wire n_7106;
wire n_38813;
wire n_27203;
wire n_14122;
wire newNet_2175;
wire n_13156;
wire newNet_3204;
wire n_44764;
wire n_27574;
wire n_27036;
wire n_18005;
wire n_6001;
wire n_4134;
wire n_19752;
wire n_35657;
wire n_17925;
wire n_41853;
wire FE_RN_336_0;
wire n_18789;
wire newNet_109;
wire n_38516;
wire FE_OCP_RBN1730_n_22492;
wire n_31765;
wire n_21294;
wire n_16646;
wire n_2326;
wire n_1722;
wire n_17825;
wire n_39786;
wire n_1557;
wire n_20789;
wire newNet_3238;
wire n_31488;
wire n_1253;
wire n_35534;
wire n_24308;
wire n_21435;
wire n_40087;
wire delay_add_ln22_unr20_stage8_stallmux_q_27_;
wire n_15264;
wire n_14298;
wire FE_OFN787_n_25834;
wire n_40375;
wire n_42455;
wire n_21975;
wire n_24332;
wire n_13444;
wire n_40353;
wire n_33457;
wire n_21441;
wire n_15829;
wire FE_OFN803_n_46285;
wire n_35469;
wire n_19985;
wire n_4723;
wire n_6236;
wire newNet_923;
wire n_983;
wire n_4753;
wire n_42841;
wire n_19865;
wire n_26364;
wire n_31444;
wire n_14100;
wire n_16854;
wire n_9917;
wire n_31780;
wire n_36460;
wire n_42046;
wire n_25614;
wire n_42016;
wire n_4412;
wire n_14845;
wire n_11232;
wire n_17462;
wire n_29733;
wire delay_add_ln22_unr27_stage10_stallmux_q_0_;
wire newNet_1517;
wire n_3057;
wire n_28725;
wire n_46961;
wire n_21957;
wire n_19485;
wire n_26940;
wire n_40642;
wire n_34173;
wire n_36117;
wire FE_RN_59_0;
wire n_35146;
wire n_28415;
wire n_41774;
wire n_40047;
wire n_20504;
wire n_31327;
wire n_39681;
wire n_28360;
wire n_12731;
wire n_9130;
wire n_23883;
wire n_15709;
wire n_27371;
wire n_12287;
wire n_5097;
wire n_5329;
wire n_43371;
wire n_8248;
wire n_7749;
wire n_3310;
wire n_20866;
wire n_17792;
wire n_41343;
wire n_41931;
wire newNet_2623;
wire n_3922;
wire FE_RN_1802_0;
wire n_28495;
wire newNet_3475;
wire n_11669;
wire n_10362;
wire n_22584;
wire newNet_1366;
wire n_18684;
wire n_17983;
wire n_41564;
wire n_31887;
wire newNet_729;
wire n_29062;
wire n_25293;
wire n_27381;
wire n_24026;
wire n_22264;
wire n_12599;
wire n_24711;
wire n_9489;
wire n_30952;
wire n_9042;
wire n_7984;
wire FE_RN_681_0;
wire n_37657;
wire n_12787;
wire FE_OCPN1853_n_13366;
wire n_28550;
wire n_8030;
wire n_45200;
wire beta_30;
wire n_12317;
wire n_39375;
wire newNet_2680;
wire n_26602;
wire n_2253;
wire n_13932;
wire n_717;
wire n_382;
wire n_4714;
wire n_37465;
wire n_23394;
wire n_13114;
wire newNet_1472;
wire n_2995;
wire n_27108;
wire newNet_2814;
wire newNet_580;
wire FE_RN_1835_0;
wire FE_OCP_RBN2584_n_3858;
wire n_8452;
wire n_4804;
wire n_16764;
wire FE_OCPN1396_n_7881;
wire n_42276;
wire FE_RN_1486_0;
wire n_13074;
wire n_39833;
wire n_32960;
wire newNet_301;
wire n_1489;
wire n_5290;
wire n_41461;
wire n_23476;
wire FE_RN_624_0;
wire n_36882;
wire n_17036;
wire n_31041;
wire n_32901;
wire n_19946;
wire n_1392;
wire n_37037;
wire newNet_2503;
wire n_40318;
wire n_22760;
wire n_12900;
wire n_16881;
wire n_21402;
wire n_5080;
wire n_26493;
wire n_29963;
wire n_3055;
wire n_28354;
wire n_34585;
wire n_20817;
wire n_23371;
wire n_32486;
wire n_15393;
wire n_29590;
wire n_29481;
wire FE_RN_950_0;
wire n_41424;
wire n_36089;
wire n_38045;
wire n_13917;
wire newNet_362;
wire newNet_3272;
wire FE_OCP_RBN2139_n_17547;
wire n_32860;
wire n_33162;
wire n_6772;
wire n_18152;
wire n_476;
wire n_11853;
wire n_1346;
wire n_33931;
wire n_43553;
wire n_23141;
wire n_3473;
wire n_20482;
wire n_23327;
wire newNet_1916;
wire n_31303;
wire n_768;
wire n_16904;
wire n_7991;
wire n_10849;
wire FE_OCPN1481_n_22207;
wire n_19522;
wire n_30559;
wire n_22273;
wire n_4905;
wire n_41488;
wire n_22385;
wire n_17771;
wire n_16515;
wire n_37415;
wire n_4761;
wire FE_OCP_RBN3691_n_10567;
wire newNet_711;
wire n_29674;
wire FE_OCP_RBN2301_n_7817;
wire n_23971;
wire n_29536;
wire newNet_397;
wire n_27888;
wire n_20970;
wire n_16656;
wire n_7031;
wire FE_OCP_DRV_N1605_n_31445;
wire n_35410;
wire n_37049;
wire n_34593;
wire n_46179;
wire n_24498;
wire newNet_2923;
wire n_27102;
wire n_21323;
wire newNet_753;
wire n_32075;
wire n_21842;
wire n_38227;
wire n_710;
wire n_39353;
wire n_8274;
wire n_10350;
wire n_19126;
wire FE_RN_1419_0;
wire n_42779;
wire n_14270;
wire FE_OCPN3780_n_16440;
wire n_3778;
wire n_35326;
wire n_23252;
wire n_14256;
wire n_667;
wire n_4069;
wire n_33471;
wire newNet_2589;
wire n_42826;
wire n_13422;
wire n_22792;
wire n_5052;
wire n_21044;
wire n_3781;
wire n_1333;
wire n_32183;
wire n_14507;
wire n_40192;
wire n_37760;
wire n_26180;
wire n_42702;
wire n_30145;
wire n_19820;
wire FE_RN_1026_0;
wire n_35023;
wire n_39918;
wire n_10207;
wire FE_OCP_RBN2296_n_2438;
wire n_37704;
wire FE_OCP_RBN2436_n_14072;
wire n_38441;
wire n_12290;
wire n_10086;
wire n_40445;
wire newNet_2196;
wire FE_RN_600_0;
wire n_5729;
wire n_33793;
wire newNet_2207;
wire n_27524;
wire n_24940;
wire n_14140;
wire n_40057;
wire n_33688;
wire n_1702;
wire n_33386;
wire n_42056;
wire n_37770;
wire n_38187;
wire n_29862;
wire n_42137;
wire newNet_1401;
wire n_7629;
wire n_923;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_14_;
wire n_9603;
wire n_8016;
wire n_31993;
wire newNet_1575;
wire n_43818;
wire n_1525;
wire n_27928;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_16_;
wire newNet_3756;
wire n_34852;
wire n_4662;
wire n_2522;
wire n_41384;
wire n_32590;
wire n_17815;
wire n_19293;
wire n_15443;
wire n_31698;
wire n_22605;
wire n_22209;
wire n_9229;
wire n_2441;
wire FE_OCP_RBN3432_n_33664;
wire n_3231;
wire FE_RN_1195_0;
wire n_28994;
wire n_27298;
wire n_46243;
wire FE_OCPN1500_n_26125;
wire n_32697;
wire n_1818;
wire delay_add_ln22_unr17_stage7_stallmux_q_24_;
wire n_25013;
wire n_21768;
wire n_29237;
wire n_5810;
wire FE_RN_1155_0;
wire n_21672;
wire n_21457;
wire n_44322;
wire n_26374;
wire n_23683;
wire n_41490;
wire n_31473;
wire n_4049;
wire n_3809;
wire n_4395;
wire n_21296;
wire n_17451;
wire FE_RN_941_0;
wire n_21276;
wire n_34522;
wire FE_OCP_RBN2973_n_5531;
wire n_2574;
wire n_25422;
wire n_13382;
wire n_21230;
wire n_14583;
wire n_13897;
wire n_43361;
wire FE_RN_141_0;
wire n_21287;
wire n_33005;
wire n_603;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_21_;
wire n_41624;
wire newNet_807;
wire n_42962;
wire n_13838;
wire n_12520;
wire n_29852;
wire n_26898;
wire n_7513;
wire n_38590;
wire n_4657;
wire n_40922;
wire n_41057;
wire n_43834;
wire n_6208;
wire n_33550;
wire n_13184;
wire n_42922;
wire n_3460;
wire FE_RN_323_0;
wire n_14649;
wire FE_OCP_RBN3627_n_38870;
wire n_10609;
wire n_6780;
wire FE_OFN221_n_35655;
wire n_41647;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_5_;
wire newNet_3744;
wire n_33663;
wire n_6640;
wire n_39035;
wire delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire n_36793;
wire newNet_2558;
wire n_16582;
wire n_25382;
wire newNet_944;
wire n_7669;
wire FE_OCP_RBN3360_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire n_30549;
wire n_13065;
wire n_27532;
wire FE_OCP_RBN3658_n_15314;
wire delay_xor_ln21_unr12_stage5_stallmux_q_19_;
wire FE_RN_965_0;
wire n_22118;
wire n_28437;
wire n_21375;
wire n_31203;
wire n_40728;
wire n_37204;
wire n_15717;
wire delay_xor_ln21_unr12_stage5_stallmux_q_17_;
wire n_34624;
wire n_2152;
wire n_33655;
wire n_25162;
wire n_18462;
wire FE_OCP_RBN3358_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire n_4383;
wire n_28637;
wire n_17736;
wire n_17943;
wire n_11687;
wire n_1857;
wire n_9549;
wire n_29034;
wire n_1811;
wire n_23246;
wire n_1308;
wire n_22374;
wire n_32200;
wire n_34913;
wire n_17288;
wire n_1097;
wire n_11242;
wire FE_OCP_RBN2211_n_37720;
wire n_9342;
wire n_46958;
wire n_8871;
wire n_22313;
wire n_1059;
wire n_17769;
wire n_23892;
wire n_9832;
wire n_26964;
wire n_30876;
wire FE_RN_841_0;
wire n_13015;
wire n_40399;
wire n_42724;
wire n_41176;
wire n_32779;
wire n_42641;
wire n_20433;
wire newNet_425;
wire n_40200;
wire n_41846;
wire newNet_1272;
wire n_3903;
wire n_684;
wire FE_OCPN1771_n_26801;
wire FE_OCP_RBN2896_n_39575;
wire n_31187;
wire n_12221;
wire newNet_1956;
wire newNet_2033;
wire n_23167;
wire n_34630;
wire n_17917;
wire n_38323;
wire n_35434;
wire n_19642;
wire n_10684;
wire n_9212;
wire n_18042;
wire n_9189;
wire n_17410;
wire n_43912;
wire n_39436;
wire n_36094;
wire n_28489;
wire n_10585;
wire sin_out_15;
wire n_31512;
wire n_32585;
wire n_27599;
wire n_32423;
wire newNet_3547;
wire n_32290;
wire newNet_2832;
wire n_40022;
wire n_41699;
wire FE_OCP_RBN2254_n_33729;
wire n_15017;
wire n_8733;
wire n_14746;
wire n_27275;
wire n_40100;
wire n_22259;
wire n_4649;
wire n_29915;
wire n_30576;
wire n_13496;
wire n_4941;
wire n_7818;
wire n_3456;
wire delay_add_ln22_unr20_stage8_stallmux_q_28_;
wire n_38075;
wire n_950;
wire newNet_3571;
wire n_38750;
wire n_27010;
wire n_28678;
wire n_24621;
wire n_27681;
wire n_41888;
wire n_44150;
wire n_25388;
wire newNet_3186;
wire n_1509;
wire n_16548;
wire n_6012;
wire n_40456;
wire n_8914;
wire n_6790;
wire n_25730;
wire n_20916;
wire n_9860;
wire n_2005;
wire n_6762;
wire delay_xor_ln21_unr15_stage6_stallmux_q_7_;
wire n_3642;
wire n_8820;
wire n_38801;
wire n_23788;
wire n_3545;
wire FE_OCPN1530_n_26090;
wire n_2584;
wire FE_RN_857_0;
wire n_42460;
wire n_37065;
wire n_3196;
wire n_37144;
wire n_1219;
wire newNet_2501;
wire n_12458;
wire n_1010;
wire n_1102;
wire n_38628;
wire n_38543;
wire n_526;
wire n_20266;
wire newNet_341;
wire n_13171;
wire n_8052;
wire newNet_166;
wire FE_RN_1857_0;
wire n_26428;
wire FE_OCP_RBN3433_n_33664;
wire n_4690;
wire n_12886;
wire n_37282;
wire n_22098;
wire n_9553;
wire FE_OCPN1426_n_18099;
wire n_12544;
wire n_31070;
wire newNet_342;
wire n_25473;
wire n_61;
wire n_37493;
wire n_16702;
wire n_40514;
wire n_38217;
wire n_41698;
wire n_5915;
wire n_22305;
wire n_4115;
wire FE_RN_391_0;
wire n_26700;
wire n_10082;
wire n_17492;
wire n_19061;
wire n_11484;
wire n_4959;
wire n_20014;
wire n_43693;
wire n_40091;
wire n_7153;
wire n_36735;
wire n_37839;
wire n_44996;
wire FE_OCP_RBN3669_n_46982;
wire n_30012;
wire n_42740;
wire n_5965;
wire n_30949;
wire n_39081;
wire n_1519;
wire cos_out_8;
wire n_37027;
wire n_28247;
wire n_8393;
wire n_9268;
wire n_42908;
wire n_10498;
wire n_41191;
wire newNet_1685;
wire n_6771;
wire n_25928;
wire newNet_3237;
wire n_15882;
wire FE_OCP_RBN2877_n_10354;
wire n_3044;
wire FE_OCP_RBN1349_n_19270;
wire FE_OCP_RBN2847_n_39479;
wire n_16402;
wire n_41058;
wire newNet_662;
wire FE_OCP_RBN2817_n_4458;
wire n_32421;
wire n_811;
wire n_629;
wire newNet_1641;
wire n_21016;
wire n_42232;
wire n_18545;
wire n_33531;
wire n_28984;
wire newNet_3742;
wire n_37316;
wire FE_RN_530_0;
wire n_37782;
wire n_35579;
wire newNet_2516;
wire n_33166;
wire n_4864;
wire FE_RN_446_0;
wire n_36151;
wire n_937;
wire n_27494;
wire n_22247;
wire n_14793;
wire n_25147;
wire n_10825;
wire n_30969;
wire n_10463;
wire n_29604;
wire n_35170;
wire n_15792;
wire newNet_689;
wire n_10562;
wire n_26392;
wire n_14353;
wire n_47012;
wire n_22212;
wire FE_OCP_RBN1991_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire newNet_2564;
wire n_35025;
wire FE_OCP_RBN3247_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire FE_RN_628_0;
wire n_27402;
wire n_43523;
wire sin_out_29;
wire FE_OCPN1002_n_45660;
wire n_37755;
wire n_30808;
wire n_18061;
wire n_28391;
wire n_10145;
wire FE_RN_1822_0;
wire n_39326;
wire n_4267;
wire FE_OCPN3183_n_22294;
wire n_32456;
wire newNet_3262;
wire n_17439;
wire n_41839;
wire n_40299;
wire n_40181;
wire FE_RN_1347_0;
wire n_6521;
wire n_23894;
wire n_4097;
wire n_32292;
wire n_222;
wire n_40073;
wire n_33728;
wire n_27812;
wire n_2777;
wire n_506;
wire n_4582;
wire n_32485;
wire n_15567;
wire n_16682;
wire n_37361;
wire n_27247;
wire n_38058;
wire n_11416;
wire n_17487;
wire n_10238;
wire n_42334;
wire n_42470;
wire n_42663;
wire n_34187;
wire n_37205;
wire n_12064;
wire n_35238;
wire n_28262;
wire n_29506;
wire newNet_3416;
wire n_25555;
wire delay_add_ln22_unr27_stage10_stallmux_q_9_;
wire FE_OCP_RBN2545_n_44944;
wire newNet_3042;
wire delay_xor_ln22_unr3_stage2_stallmux_q_7_;
wire n_28960;
wire n_1005;
wire n_12162;
wire n_24816;
wire n_11244;
wire FE_OCP_RBN2319_n_2367;
wire newNet_3577;
wire n_12288;
wire n_28254;
wire n_37817;
wire n_18246;
wire n_38790;
wire newNet_3187;
wire n_6939;
wire n_43237;
wire newNet_3100;
wire n_6836;
wire n_19826;
wire n_43528;
wire n_36558;
wire FE_OCP_RBN3715_n_39913;
wire newNet_648;
wire n_7775;
wire newNet_509;
wire n_36542;
wire FE_RN_742_0;
wire n_15105;
wire n_6823;
wire n_41453;
wire n_41863;
wire n_15118;
wire n_2847;
wire n_26773;
wire n_43819;
wire n_41399;
wire n_3116;
wire FE_OCP_RBN2394_n_8288;
wire n_10903;
wire n_40553;
wire n_31294;
wire n_6929;
wire n_33554;
wire n_2884;
wire n_35281;
wire n_41852;
wire FE_RN_133_0;
wire FE_OFN794_n_45813;
wire n_954;
wire n_15656;
wire n_34181;
wire FE_RN_492_0;
wire n_2141;
wire n_15910;
wire newNet_2238;
wire n_37109;
wire n_32929;
wire n_33588;
wire n_43126;
wire n_2041;
wire n_11393;
wire FE_RN_1185_0;
wire n_25353;
wire n_5454;
wire n_45812;
wire FE_OCP_RBN3530_n_13765;
wire delay_add_ln22_unr17_stage7_stallmux_q_0_;
wire n_10731;
wire FE_OCPN1016_n_23307;
wire n_597;
wire n_1666;
wire delay_add_ln22_unr8_stage4_stallmux_q_2_;
wire n_8613;
wire n_23192;
wire n_8638;
wire n_7057;
wire n_11635;
wire n_43085;
wire n_21974;
wire n_95;
wire n_42600;
wire n_34376;
wire n_38857;
wire n_17456;
wire n_15277;
wire n_11166;
wire n_22689;
wire n_4210;
wire n_7344;
wire n_27000;
wire n_14718;
wire n_46145;
wire newNet_1482;
wire n_42923;
wire n_30029;
wire n_19841;
wire n_32491;
wire n_2375;
wire n_17223;
wire n_1124;
wire n_27628;
wire FE_RN_1088_0;
wire n_29230;
wire FE_RN_1071_0;
wire n_13999;
wire n_40151;
wire n_22307;
wire n_6843;
wire n_3026;
wire FE_OCPN992_n_22249;
wire n_29535;
wire n_36608;
wire n_39576;
wire FE_OCP_RBN2663_n_20333;
wire n_35159;
wire newNet_1577;
wire n_14177;
wire n_19177;
wire n_23676;
wire n_19690;
wire n_26352;
wire newNet_1969;
wire n_39007;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_14_;
wire n_2357;
wire n_41183;
wire n_18428;
wire n_25011;
wire n_25693;
wire n_23234;
wire n_7399;
wire n_42344;
wire n_17748;
wire newNet_1887;
wire FE_OCP_RBN3420_n_12739;
wire n_3458;
wire newNet_412;
wire n_5101;
wire newNet_870;
wire n_26389;
wire n_13645;
wire n_43782;
wire newNet_1494;
wire FE_RN_876_0;
wire n_15205;
wire n_22387;
wire n_27685;
wire n_27154;
wire n_19357;
wire n_10967;
wire n_23919;
wire n_21678;
wire n_422;
wire n_26718;
wire newNet_806;
wire n_7071;
wire n_42377;
wire n_16134;
wire n_40655;
wire n_34700;
wire newNet_1037;
wire n_10716;
wire FE_OCP_RBN2535_n_47018;
wire n_26633;
wire n_21258;
wire n_33056;
wire newNet_1265;
wire n_18380;
wire n_40242;
wire newNet_2195;
wire n_7650;
wire n_7795;
wire n_30452;
wire n_38997;
wire FE_OCP_RBN2800_n_15706;
wire n_18587;
wire n_17816;
wire newNet_2367;
wire n_42383;
wire n_9357;
wire n_8010;
wire n_11233;
wire FE_OCP_RBN2309_n_29298;
wire n_14585;
wire n_29675;
wire n_35123;
wire n_12415;
wire n_44831;
wire n_27263;
wire FE_RN_889_0;
wire n_12294;
wire n_38164;
wire FE_RN_1785_0;
wire n_17686;
wire n_25038;
wire n_33021;
wire n_1546;
wire n_13440;
wire n_43788;
wire n_24044;
wire n_32584;
wire n_34538;
wire n_16169;
wire n_3485;
wire n_40790;
wire n_12328;
wire FE_RN_562_0;
wire n_42176;
wire n_24531;
wire n_38802;
wire n_17356;
wire newNet_2073;
wire n_19146;
wire FE_OCPN1482_n_22207;
wire n_12097;
wire n_21065;
wire n_20842;
wire n_20850;
wire n_24119;
wire n_9071;
wire n_24656;
wire newNet_1348;
wire FE_OCP_RBN2748_n_9584;
wire FE_OCP_RBN1143_n_29292;
wire n_30472;
wire n_27269;
wire n_46366;
wire n_17037;
wire n_16855;
wire n_35435;
wire n_15779;
wire n_40376;
wire n_43148;
wire n_39548;
wire newNet_952;
wire n_3873;
wire n_13746;
wire n_35876;
wire n_33775;
wire n_16455;
wire n_15529;
wire n_43511;
wire n_39016;
wire newNet_2015;
wire n_1881;
wire FE_OCP_RBN3411_n_33547;
wire FE_RN_1753_0;
wire n_36217;
wire n_38754;
wire n_37110;
wire n_27939;
wire n_6082;
wire delay_xor_ln21_unr9_stage4_stallmux_q_10_;
wire n_37892;
wire n_29877;
wire n_32847;
wire n_20379;
wire n_2803;
wire newNet_3280;
wire newNet_3011;
wire n_193;
wire n_9406;
wire n_39262;
wire n_18930;
wire newNet_3286;
wire n_33434;
wire n_19858;
wire n_39222;
wire n_38401;
wire n_33100;
wire n_41127;
wire n_3739;
wire FE_RN_677_0;
wire n_13321;
wire n_4306;
wire n_9831;
wire n_18809;
wire newNet_1378;
wire n_21108;
wire n_40691;
wire newNet_2090;
wire n_8421;
wire n_13473;
wire n_35821;
wire FE_OCP_RBN2492_n_8508;
wire n_26303;
wire n_9314;
wire n_13487;
wire newNet_2123;
wire n_42802;
wire n_32532;
wire n_19173;
wire n_655;
wire n_5742;
wire n_35147;
wire n_8379;
wire FE_OCPN1395_n_7881;
wire n_13822;
wire n_4341;
wire n_28202;
wire newNet_2528;
wire n_42351;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_18_;
wire FE_RN_1149_0;
wire n_5727;
wire n_5477;
wire FE_RN_806_0;
wire newNet_1385;
wire n_1756;
wire n_12690;
wire n_783;
wire FE_OCP_RBN3731_n_31819;
wire n_41428;
wire n_16825;
wire newNet_34;
wire n_16619;
wire n_15699;
wire n_43860;
wire n_117;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_5_;
wire FE_OCPN1796_n_30546;
wire n_10886;
wire n_38987;
wire newNet_2792;
wire n_25232;
wire n_15300;
wire delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire n_42205;
wire newNet_907;
wire n_36465;
wire n_1135;
wire n_39534;
wire n_42959;
wire n_12788;
wire FE_OCP_RBN2215_FE_OCPN950_n_28595;
wire n_5398;
wire n_8370;
wire n_32743;
wire n_26385;
wire n_24314;
wire n_9006;
wire FE_OCP_RBN2966_n_26231;
wire n_38695;
wire n_41940;
wire n_11897;
wire n_31186;
wire n_27598;
wire n_27126;
wire n_22653;
wire n_36301;
wire n_24639;
wire newNet_2817;
wire n_20668;
wire n_32098;
wire n_15788;
wire n_30098;
wire n_24698;
wire n_26060;
wire n_39638;
wire n_13594;
wire n_36039;
wire n_26832;
wire n_10241;
wire n_38258;
wire n_11619;
wire n_20338;
wire n_22770;
wire n_39566;
wire n_22135;
wire newNet_3404;
wire n_14567;
wire n_26686;
wire n_2211;
wire n_5611;
wire n_18771;
wire FE_OCP_RBN2668_n_4158;
wire n_449;
wire FE_RN_1450_0;
wire n_30996;
wire n_41011;
wire n_39411;
wire FE_OCP_RBN2295_n_2438;
wire n_23838;
wire n_37718;
wire n_18506;
wire n_26500;
wire n_23288;
wire n_22791;
wire n_39820;
wire n_27907;
wire n_4426;
wire n_37005;
wire FE_OCP_RBN2489_n_3338;
wire n_30288;
wire n_11580;
wire n_23601;
wire n_13759;
wire n_24368;
wire n_40811;
wire n_16203;
wire n_13265;
wire n_37370;
wire delay_add_ln22_unr23_stage9_stallmux_q_0_;
wire FE_RN_1567_0;
wire FE_RN_520_0;
wire n_35565;
wire n_18973;
wire n_40762;
wire n_43250;
wire n_31930;
wire FE_OCP_RBN2791_n_9910;
wire n_21388;
wire n_25331;
wire n_36349;
wire n_13231;
wire n_22076;
wire n_10676;
wire newNet_875;
wire n_25731;
wire n_27896;
wire n_4508;
wire n_38885;
wire n_18749;
wire n_18479;
wire n_36111;
wire newNet_3653;
wire n_16743;
wire n_43660;
wire n_28490;
wire FE_RN_1395_0;
wire n_26802;
wire n_28824;
wire FE_RN_153_0;
wire n_21030;
wire n_18639;
wire n_30243;
wire n_1103;
wire n_33807;
wire n_29;
wire newNet_1309;
wire n_20904;
wire n_2505;
wire n_27329;
wire newNet_3140;
wire n_9890;
wire n_16210;
wire n_42045;
wire n_39763;
wire newNet_3353;
wire n_1204;
wire n_19112;
wire n_18194;
wire n_39967;
wire n_17798;
wire FE_RN_610_0;
wire FE_OFN76_n_5397;
wire n_7444;
wire FE_OCP_RBN2431_n_14018;
wire n_22471;
wire n_29001;
wire n_42659;
wire n_21078;
wire n_14590;
wire n_17471;
wire n_14271;
wire n_28744;
wire newNet_3145;
wire newNet_931;
wire FE_RN_251_0;
wire n_4954;
wire FE_OCP_RBN2699_n_4238;
wire n_37632;
wire newNet_2963;
wire n_40193;
wire n_32471;
wire n_18397;
wire newNet_3666;
wire n_42085;
wire n_28453;
wire n_7527;
wire n_23972;
wire n_6309;
wire n_9810;
wire n_36863;
wire n_16677;
wire n_22973;
wire n_18230;
wire n_37856;
wire newNet_2927;
wire n_22379;
wire n_36644;
wire newNet_3458;
wire n_10860;
wire n_32436;
wire n_6158;
wire n_17973;
wire n_17280;
wire n_25096;
wire n_25440;
wire n_21508;
wire n_13869;
wire newNet_1933;
wire n_37446;
wire FE_OCPN3784_FE_OCP_RBN2831_n_10198;
wire FE_RN_1744_0;
wire n_29610;
wire n_11504;
wire n_19623;
wire newNet_1147;
wire n_31381;
wire n_29823;
wire n_42112;
wire n_17944;
wire n_31677;
wire n_9091;
wire n_36221;
wire n_7294;
wire n_23472;
wire n_40676;
wire newNet_2588;
wire delay_add_ln22_unr14_stage6_stallmux_q_20_;
wire n_21592;
wire newNet_1088;
wire n_929;
wire FE_RN_840_0;
wire n_31915;
wire n_27059;
wire n_32616;
wire n_4074;
wire n_41319;
wire n_37292;
wire n_19526;
wire n_14656;
wire n_6879;
wire FE_OCP_RBN1094_n_45224;
wire n_21242;
wire n_41265;
wire n_28364;
wire n_33843;
wire n_8970;
wire n_12988;
wire n_20949;
wire n_19901;
wire n_16183;
wire n_16132;
wire n_34626;
wire n_23888;
wire n_24229;
wire n_40574;
wire n_34223;
wire n_9021;
wire n_30125;
wire newNet_2144;
wire n_24675;
wire n_10382;
wire n_8102;
wire n_35884;
wire n_10786;
wire n_42689;
wire n_41159;
wire n_26658;
wire n_10942;
wire n_11685;
wire n_16259;
wire n_9587;
wire FE_RN_1370_0;
wire FE_RN_411_0;
wire n_25581;
wire newNet_1456;
wire n_15857;
wire n_3844;
wire n_484;
wire n_14028;
wire n_1691;
wire n_5315;
wire n_11427;
wire n_22002;
wire n_36219;
wire n_40337;
wire n_12442;
wire n_28976;
wire n_39957;
wire n_26471;
wire n_6760;
wire n_35366;
wire n_2239;
wire n_10980;
wire n_38809;
wire n_24776;
wire n_9595;
wire newNet_1829;
wire n_7554;
wire n_26104;
wire n_14964;
wire n_35556;
wire FE_OCP_RBN3009_n_31117;
wire n_42051;
wire newNet_2522;
wire n_4966;
wire n_38170;
wire n_32025;
wire n_12014;
wire n_4094;
wire n_42443;
wire n_35331;
wire n_21892;
wire n_30162;
wire newNet_1659;
wire n_42770;
wire newNet_845;
wire cordic_combinational_sub_ln23_0_unr20_z_0_;
wire FE_OCP_RBN1702_n_19560;
wire n_33372;
wire n_13497;
wire n_28215;
wire n_22586;
wire n_13172;
wire newNet_2944;
wire delay_add_ln22_unr17_stage7_stallmux_q_19_;
wire n_31779;
wire FE_OCP_RBN1921_n_22476;
wire n_27644;
wire n_42169;
wire n_18731;
wire FE_RN_1583_0;
wire n_37905;
wire newNet_3397;
wire n_30157;
wire n_2279;
wire n_42034;
wire n_33486;
wire FE_OCP_RBN3674_FE_RN_1581_0;
wire n_21884;
wire n_35857;
wire n_8905;
wire n_38472;
wire FE_OCP_RBN2447_n_14114;
wire n_34854;
wire n_25824;
wire FE_OCP_RBN2808_n_35285;
wire n_26763;
wire FE_OCP_RBN3733_n_31819;
wire newNet_3270;
wire n_37198;
wire n_3774;
wire FE_OCP_RBN1847_n_22068;
wire n_8716;
wire n_11057;
wire n_32817;
wire n_24661;
wire n_44030;
wire FE_OCP_RBN3587_n_47016;
wire n_29985;
wire n_17287;
wire n_13326;
wire n_32163;
wire n_19972;
wire n_35084;
wire FE_RN_1637_0;
wire n_4131;
wire newNet_2402;
wire n_14430;
wire n_19206;
wire n_13267;
wire n_18280;
wire n_19223;
wire n_32852;
wire n_26252;
wire n_26159;
wire n_15047;
wire n_14610;
wire n_3805;
wire n_26093;
wire FE_RN_1259_0;
wire newNet_1159;
wire n_38200;
wire newNet_320;
wire n_6593;
wire n_27054;
wire newNet_3122;
wire n_24932;
wire n_7605;
wire n_15504;
wire n_36284;
wire n_31130;
wire n_23325;
wire FE_RN_1872_0;
wire n_34921;
wire n_28085;
wire n_3883;
wire n_36329;
wire n_8078;
wire n_27362;
wire FE_OCP_RBN3081_n_16977;
wire n_38367;
wire n_6996;
wire n_24390;
wire delay_xor_ln22_unr21_stage8_stallmux_q_5_;
wire n_36687;
wire newNet_3363;
wire n_2834;
wire n_5910;
wire n_27428;
wire n_19569;
wire n_15133;
wire n_4915;
wire n_20029;
wire FE_RN_392_0;
wire n_35865;
wire n_30772;
wire n_27250;
wire newNet_1067;
wire n_37597;
wire n_39487;
wire FE_OCP_RBN2542_n_38721;
wire n_15683;
wire n_36069;
wire n_35575;
wire FE_OCP_RBN2501_n_13896;
wire newNet_819;
wire n_3780;
wire FE_RN_1659_0;
wire n_7788;
wire newNet_143;
wire n_4396;
wire n_20791;
wire FE_OCPN1025_n_25481;
wire n_27869;
wire n_31680;
wire n_13255;
wire newNet_915;
wire n_12614;
wire n_21538;
wire n_2053;
wire FE_OCP_RBN3022_n_39942;
wire FE_OCP_RBN2227_n_7598;
wire n_31172;
wire n_10071;
wire n_27426;
wire n_8119;
wire n_22732;
wire n_14505;
wire n_3397;
wire n_42987;
wire n_18780;
wire FE_RN_145_0;
wire FE_OCP_RBN3588_n_9408;
wire n_31457;
wire n_43609;
wire n_42222;
wire n_37673;
wire n_17869;
wire n_15621;
wire n_5045;
wire n_45844;
wire n_8980;
wire n_7798;
wire n_21778;
wire n_40660;
wire n_10248;
wire n_36323;
wire n_29071;
wire n_33173;
wire n_30065;
wire FE_OCP_RBN2687_n_38870;
wire n_15934;
wire n_20065;
wire n_44356;
wire delay_add_ln22_unr27_stage10_stallmux_q_29_;
wire n_38319;
wire n_14216;
wire n_12336;
wire n_29757;
wire FE_RN_214_0;
wire n_24048;
wire n_27450;
wire FE_OCPN1384_n_18345;
wire newNet_2331;
wire newNet_93;
wire n_13958;
wire n_24456;
wire newNet_296;
wire n_2908;
wire n_26909;
wire n_15984;
wire n_6722;
wire n_19936;
wire n_17140;
wire FE_RN_1222_0;
wire n_23314;
wire n_13927;
wire n_19204;
wire n_35543;
wire n_4604;
wire n_16005;
wire n_39040;
wire n_12203;
wire n_1997;
wire n_39232;
wire n_30937;
wire n_38553;
wire n_39807;
wire FE_OCP_RBN2442_n_8402;
wire FE_RN_99_0;
wire n_32824;
wire n_38915;
wire newNet_1760;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_17_;
wire n_8159;
wire n_16425;
wire n_24215;
wire n_16823;
wire n_33130;
wire n_31589;
wire n_34467;
wire newNet_1018;
wire n_1626;
wire n_42252;
wire n_43497;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_12_;
wire FE_OCP_RBN2330_n_9003;
wire n_36412;
wire n_32678;
wire FE_RN_1301_0;
wire newNet_2855;
wire newNet_478;
wire FE_OCP_RBN3415_n_12739;
wire n_23028;
wire n_19661;
wire FE_RN_1589_0;
wire n_45659;
wire n_530;
wire n_17783;
wire n_33645;
wire n_27968;
wire newNet_2478;
wire n_41133;
wire n_19294;
wire n_6824;
wire n_23645;
wire n_36237;
wire n_2635;
wire delay_sub_ln21_0_unr5_stage3_stallmux_q_3_;
wire n_45887;
wire n_8163;
wire n_2392;
wire n_4739;
wire n_21899;
wire n_34479;
wire n_16562;
wire n_1724;
wire n_3331;
wire n_14447;
wire n_37177;
wire n_34513;
wire n_15722;
wire n_23643;
wire n_22443;
wire n_1872;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_20_;
wire n_31461;
wire n_46183;
wire n_27356;
wire n_34304;
wire n_24161;
wire n_41214;
wire n_18035;
wire n_5411;
wire n_9897;
wire n_19956;
wire n_12963;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_19_;
wire n_31788;
wire FE_OCPUNCON1803_n_18111;
wire n_23124;
wire n_17674;
wire n_8863;
wire n_33346;
wire n_20086;
wire FE_OCP_RBN3572_n_44563;
wire n_38592;
wire n_27237;
wire n_3960;
wire n_40;
wire n_36759;
wire n_17950;
wire n_17852;
wire n_17504;
wire n_16552;
wire n_34146;
wire n_42018;
wire n_27449;
wire FE_OCP_RBN3364_n_44722;
wire n_23860;
wire FE_OCP_RBN3368_n_32436;
wire n_39306;
wire n_29437;
wire n_34004;
wire n_34749;
wire n_18449;
wire newNet_2785;
wire n_3222;
wire n_8833;
wire n_43838;
wire n_39161;
wire n_35056;
wire n_20173;
wire newNet_16;
wire cos_out_23;
wire n_14631;
wire n_22341;
wire n_13146;
wire n_17985;
wire n_9915;
wire n_43573;
wire newNet_2753;
wire n_39106;
wire n_27624;
wire n_29443;
wire newNet_3614;
wire n_7882;
wire n_11434;
wire FE_RN_1211_0;
wire FE_OCPN1503_n_47257;
wire n_41800;
wire FE_RN_1685_0;
wire n_34152;
wire n_27080;
wire n_20831;
wire n_26478;
wire n_2555;
wire n_25310;
wire n_17325;
wire n_41152;
wire newNet_3028;
wire n_12396;
wire n_46215;
wire n_14249;
wire n_37405;
wire n_28090;
wire n_9365;
wire n_43443;
wire n_24246;
wire n_8543;
wire newNet_2432;
wire n_35459;
wire n_15430;
wire n_24549;
wire n_912;
wire n_10836;
wire FE_OCP_RBN2623_n_3631;
wire n_46230;
wire n_23656;
wire n_18623;
wire n_34070;
wire n_1712;
wire n_1091;
wire n_42832;
wire n_43615;
wire FE_OCP_RBN2126_n_44734;
wire n_3758;
wire n_368;
wire n_46940;
wire FE_OCP_RBN2134_n_45508;
wire n_18605;
wire n_4314;
wire n_35471;
wire n_42527;
wire n_1178;
wire n_24553;
wire n_31906;
wire n_37188;
wire n_12677;
wire n_25747;
wire n_8404;
wire newNet_3025;
wire n_14927;
wire n_17339;
wire n_3989;
wire n_480;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_17_;
wire n_28160;
wire n_26698;
wire n_2425;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_24_;
wire n_1613;
wire n_9503;
wire n_10529;
wire n_13023;
wire n_26132;
wire n_24177;
wire n_5546;
wire n_8029;
wire n_34109;
wire n_17421;
wire n_2416;
wire newNet_1070;
wire n_22832;
wire n_34316;
wire n_20638;
wire n_755;
wire n_5595;
wire FE_OCP_RBN2990_n_35539;
wire newNet_282;
wire n_7982;
wire n_14414;
wire n_28835;
wire n_2188;
wire n_3130;
wire n_41320;
wire n_43569;
wire delay_xor_ln22_unr12_stage5_stallmux_q_16_;
wire n_4497;
wire n_4457;
wire n_42644;
wire n_1900;
wire n_23816;
wire n_1714;
wire n_37398;
wire n_30911;
wire n_15868;
wire n_15645;
wire n_30403;
wire n_25502;
wire n_23344;
wire newNet_3469;
wire n_9462;
wire n_12507;
wire n_46163;
wire n_1487;
wire n_16283;
wire n_14712;
wire n_38338;
wire n_9520;
wire n_21874;
wire n_18241;
wire FE_RN_264_0;
wire n_31617;
wire sin_out_20;
wire FE_RN_1582_0;
wire n_43219;
wire n_1294;
wire n_278;
wire n_35089;
wire FE_OCP_RBN3114_n_6379;
wire n_32958;
wire n_24352;
wire n_36007;
wire n_12822;
wire n_36832;
wire newNet_2714;
wire n_21988;
wire n_26562;
wire n_10764;
wire n_36930;
wire n_5566;
wire n_2308;
wire newNet_1143;
wire n_12448;
wire n_6259;
wire n_12357;
wire n_5225;
wire n_22894;
wire FE_OCP_RBN2146_FE_OCPN861_n_45450;
wire n_36335;
wire n_10582;
wire n_32716;
wire n_12627;
wire FE_OCP_RBN3400_n_37670;
wire n_29884;
wire n_46962;
wire n_35624;
wire n_786;
wire n_14327;
wire n_39556;
wire FE_RN_1831_0;
wire FE_RN_964_0;
wire n_32008;
wire n_30049;
wire FE_OCP_RBN1851_n_22556;
wire n_17193;
wire n_3949;
wire n_14993;
wire newNet_1999;
wire FE_RN_991_0;
wire n_25548;
wire n_40032;
wire n_34857;
wire n_27648;
wire n_11908;
wire n_21606;
wire n_20076;
wire newNet_3436;
wire FE_OCP_RBN1713_FE_RN_664_0;
wire n_34944;
wire newNet_1796;
wire n_37157;
wire n_29094;
wire n_12432;
wire newNet_3413;
wire n_43646;
wire n_11062;
wire n_21512;
wire n_7764;
wire n_31339;
wire n_40424;
wire n_8919;
wire n_37540;
wire n_29422;
wire FE_OCP_RBN3524_n_8242;
wire n_2280;
wire n_29168;
wire n_38730;
wire newNet_3425;
wire n_34496;
wire n_17165;
wire n_43633;
wire n_12121;
wire n_6969;
wire n_5114;
wire FE_RN_1214_0;
wire n_34364;
wire n_33019;
wire n_7410;
wire n_13840;
wire n_28422;
wire n_27436;
wire n_13000;
wire n_12460;
wire FE_RN_871_0;
wire n_41973;
wire n_19626;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_20_;
wire n_4871;
wire n_9906;
wire n_40253;
wire n_28866;
wire n_29974;
wire n_308;
wire n_1971;
wire n_10433;
wire delay_xor_ln22_unr12_stage5_stallmux_q_6_;
wire n_21832;
wire n_8629;
wire n_1753;
wire n_21856;
wire n_24738;
wire n_38811;
wire n_4449;
wire newNet_1099;
wire n_26276;
wire n_18217;
wire n_30874;
wire n_37452;
wire n_42598;
wire n_4419;
wire FE_RN_1163_0;
wire n_6299;
wire n_13533;
wire n_37351;
wire n_2133;
wire n_36310;
wire n_41679;
wire n_29564;
wire FE_RN_269_0;
wire n_16763;
wire n_36998;
wire n_43809;
wire FE_OCP_RBN2448_n_14114;
wire n_1460;
wire n_24895;
wire n_18722;
wire n_23389;
wire n_12153;
wire n_31536;
wire FE_OCP_RBN1155_n_18375;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_11_;
wire n_26852;
wire newNet_179;
wire FE_RN_120_0;
wire FE_RN_1165_0;
wire n_13129;
wire n_27038;
wire FE_OCPUNCON1805_n_19801;
wire n_7450;
wire n_39876;
wire n_35048;
wire n_6122;
wire n_29696;
wire n_40419;
wire n_37120;
wire n_4372;
wire n_19472;
wire n_3370;
wire n_3973;
wire n_10258;
wire n_16759;
wire n_39913;
wire n_27590;
wire newNet_1341;
wire n_23604;
wire n_26681;
wire n_26934;
wire n_8973;
wire n_39851;
wire n_6890;
wire n_14304;
wire n_9019;
wire n_43389;
wire n_7950;
wire n_39689;
wire n_156;
wire n_32088;
wire n_31559;
wire FE_OCP_RBN3543_n_44575;
wire delay_add_ln22_unr2_stage2_stallmux_q_14_;
wire n_39431;
wire n_6160;
wire n_26896;
wire n_19552;
wire FE_RN_396_0;
wire n_8512;
wire n_2348;
wire FE_OCP_RBN2661_n_9292;
wire n_16928;
wire n_13850;
wire n_34344;
wire n_37087;
wire n_40283;
wire n_15228;
wire n_38655;
wire n_2612;
wire FE_OCPUNCON1802_n_29375;
wire FE_OCP_RBN1332_n_20249;
wire n_26879;
wire n_24976;
wire newNet_2575;
wire n_29251;
wire newNet_3540;
wire newNet_1239;
wire n_19169;
wire n_7227;
wire n_30511;
wire n_2863;
wire n_27566;
wire n_25934;
wire n_3521;
wire n_32998;
wire n_24823;
wire n_41102;
wire n_35220;
wire n_43610;
wire n_25840;
wire n_29039;
wire FE_OCP_RBN2614_n_35005;
wire n_40601;
wire n_25086;
wire n_41051;
wire newNet_946;
wire n_6953;
wire n_35644;
wire n_3582;
wire n_40089;
wire n_9012;
wire n_28620;
wire n_5165;
wire sin_out_4;
wire n_10626;
wire n_10673;
wire n_10364;
wire n_7065;
wire n_33995;
wire n_26333;
wire newNet_3107;
wire n_33310;
wire n_35179;
wire n_27334;
wire n_17526;
wire n_28327;
wire newNet_483;
wire n_18179;
wire n_28350;
wire n_1561;
wire n_38650;
wire newNet_3223;
wire n_38526;
wire n_611;
wire n_44325;
wire n_43845;
wire n_26740;
wire n_43151;
wire n_18226;
wire n_26786;
wire n_20691;
wire n_14838;
wire n_24666;
wire n_22099;
wire newNet_3539;
wire n_30231;
wire n_18919;
wire n_28720;
wire n_40933;
wire FE_OCP_RBN2113_n_45224;
wire n_37826;
wire n_31764;
wire n_19828;
wire n_5173;
wire n_34529;
wire n_36391;
wire n_46248;
wire n_550;
wire n_32692;
wire n_20835;
wire n_23702;
wire n_26001;
wire n_13198;
wire FE_OCP_RBN3431_n_33664;
wire n_2461;
wire FE_OCP_RBN3453_FE_OCPN1240_n_7721;
wire n_14762;
wire n_38783;
wire FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_;
wire n_24519;
wire FE_RN_1221_0;
wire n_14392;
wire FE_RN_1574_0;
wire n_13529;
wire n_12958;
wire n_36666;
wire n_14774;
wire n_12229;
wire n_2562;
wire n_10178;
wire newNet_2035;
wire n_5104;
wire n_32605;
wire n_22441;
wire n_39358;
wire n_21046;
wire n_39030;
wire n_16867;
wire n_25920;
wire n_33532;
wire n_22316;
wire n_37568;
wire newNet_3735;
wire n_27726;
wire FE_OCP_RBN2572_n_29922;
wire n_26136;
wire n_16506;
wire n_32197;
wire n_22666;
wire n_1008;
wire n_33038;
wire n_43358;
wire FE_OCP_RBN1990_delay_xor_ln23_unr6_stage3_stallmux_q;
wire n_20587;
wire n_262;
wire n_3824;
wire n_27015;
wire delay_add_ln22_unr23_stage9_stallmux_q_1_;
wire n_42577;
wire n_9515;
wire FE_RN_713_0;
wire n_30152;
wire FE_RN_829_0;
wire FE_RN_1128_0;
wire n_40428;
wire n_30050;
wire n_28579;
wire n_17465;
wire n_41896;
wire n_26796;
wire FE_OCP_RBN1849_n_22639;
wire FE_OCP_RBN2946_n_5428;
wire n_30091;
wire n_39921;
wire n_39675;
wire n_13894;
wire n_14519;
wire n_183;
wire n_11592;
wire n_17562;
wire n_39740;
wire n_1325;
wire n_1437;
wire n_11974;
wire n_27246;
wire n_22318;
wire n_8231;
wire n_4823;
wire n_12077;
wire n_20895;
wire n_20973;
wire FE_OCP_DRV_N3738_n_29439;
wire n_32599;
wire n_39302;
wire FE_OCP_RBN2814_n_25817;
wire n_11620;
wire n_29218;
wire newNet_832;
wire n_4366;
wire n_715;
wire FE_RN_1733_0;
wire n_21071;
wire n_38037;
wire n_43919;
wire n_33045;
wire n_17703;
wire newNet_1260;
wire FE_OCP_RBN2916_n_10644;
wire n_8911;
wire n_27143;
wire n_40265;
wire newNet_0;
wire delay_xor_ln21_unr6_stage3_stallmux_q_24_;
wire n_1886;
wire n_1528;
wire n_15434;
wire n_24593;
wire n_1904;
wire n_22031;
wire n_19327;
wire n_21142;
wire n_21024;
wire n_15695;
wire n_45740;
wire n_31281;
wire n_13389;
wire n_37418;
wire n_15535;
wire n_17321;
wire n_2177;
wire n_41667;
wire n_46174;
wire FE_OCP_RBN2104_delay_sub_ln23_unr9_stage4_stallmux_q_3_;
wire n_15631;
wire n_10127;
wire newNet_1977;
wire n_38212;
wire n_135;
wire FE_OCP_RBN3390_n_33108;
wire n_27210;
wire n_37843;
wire n_6490;
wire n_29785;
wire n_21795;
wire newNet_1077;
wire n_40807;
wire n_36097;
wire n_13325;
wire n_26324;
wire n_33672;
wire n_21470;
wire n_36139;
wire n_15835;
wire n_43637;
wire n_1016;
wire n_17949;
wire newNet_1369;
wire n_20917;
wire n_2787;
wire n_23176;
wire n_26201;
wire n_23535;
wire n_23259;
wire n_22049;
wire n_5582;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_11_;
wire n_3732;
wire n_3940;
wire n_8872;
wire n_2994;
wire n_25026;
wire n_35716;
wire n_27119;
wire n_21185;
wire newNet_2979;
wire n_13587;
wire n_8001;
wire n_31804;
wire n_17931;
wire n_2094;
wire n_23533;
wire n_34560;
wire n_20203;
wire n_41843;
wire n_21052;
wire n_28359;
wire n_6517;
wire n_6167;
wire FE_OCP_RBN2312_n_41420;
wire n_12455;
wire n_20144;
wire n_10376;
wire FE_RN_554_0;
wire n_38021;
wire n_26247;
wire delay_xor_ln21_unr15_stage6_stallmux_q_6_;
wire n_41830;
wire n_9783;
wire n_41534;
wire n_35970;
wire n_2421;
wire n_6178;
wire n_1338;
wire newNet_3751;
wire n_12453;
wire n_37281;
wire n_23612;
wire n_13454;
wire n_45527;
wire n_34590;
wire newNet_2215;
wire n_38535;
wire n_42584;
wire FE_RN_92_0;
wire n_28675;
wire n_27322;
wire n_30773;
wire n_14454;
wire FE_OCP_RBN2048_delay_sub_ln23_unr17_stage6_stallmux_q_1_;
wire newNet_2540;
wire newNet_556;
wire newNet_3215;
wire n_38939;
wire FE_RN_1271_0;
wire n_16768;
wire n_13522;
wire n_40107;
wire FE_OCP_DRV_N1548_n_17643;
wire n_2184;
wire n_23302;
wire n_19931;
wire n_43801;
wire n_759;
wire n_42145;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_7_;
wire n_37384;
wire n_2114;
wire n_13062;
wire n_5032;
wire n_23520;
wire n_9302;
wire n_37342;
wire n_26264;
wire n_12146;
wire n_16649;
wire n_37536;
wire n_26458;
wire FE_RN_957_0;
wire n_38007;
wire n_16578;
wire n_6651;
wire n_32349;
wire n_32236;
wire n_33344;
wire n_28063;
wire newNet_667;
wire n_34826;
wire n_15799;
wire n_42461;
wire n_33542;
wire n_35359;
wire n_16564;
wire n_41258;
wire FE_OCP_RBN3561_n_29857;
wire FE_OCP_RBN3427_n_44881;
wire n_30089;
wire newNet_1780;
wire n_28975;
wire n_37910;
wire n_26768;
wire n_28840;
wire newNet_3444;
wire n_14209;
wire n_2157;
wire FE_RN_801_0;
wire n_27737;
wire n_10032;
wire n_13361;
wire n_37986;
wire n_21951;
wire n_7509;
wire n_17229;
wire newNet_1119;
wire n_23872;
wire n_11702;
wire delay_sub_ln21_unr24_stage9_stallmux_q_1_;
wire newNet_1411;
wire n_26692;
wire n_1669;
wire newNet_2718;
wire n_34730;
wire n_16629;
wire n_21896;
wire n_396;
wire FE_OCPN974_n_46956;
wire n_42639;
wire n_10608;
wire n_31580;
wire n_19776;
wire newNet_2993;
wire n_11375;
wire n_38841;
wire n_38418;
wire FE_RN_1001_0;
wire n_22417;
wire n_20748;
wire FE_OCPN3792_n_31804;
wire n_22205;
wire n_13943;
wire n_20022;
wire delay_add_ln22_unr11_stage5_stallmux_q_7_;
wire n_9220;
wire n_1483;
wire n_12089;
wire n_24567;
wire FE_RN_626_0;
wire FE_OCP_RBN2899_n_44853;
wire n_41877;
wire n_13176;
wire n_224;
wire n_7281;
wire n_46377;
wire n_5487;
wire n_24630;
wire newNet_1300;
wire n_6893;
wire sin_out_18;
wire n_21454;
wire n_39261;
wire n_31919;
wire n_29177;
wire n_4665;
wire n_34177;
wire FE_OCPN1745_n_29420;
wire n_28859;
wire newNet_1438;
wire n_8707;
wire n_25831;
wire newNet_2675;
wire n_9202;
wire n_39273;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_7_;
wire n_2406;
wire n_16967;
wire newNet_2593;
wire n_25210;
wire n_22184;
wire n_32150;
wire n_31738;
wire n_34777;
wire n_8585;
wire n_41949;
wire n_34067;
wire FE_OCP_RBN3557_n_8687;
wire n_33270;
wire n_28447;
wire n_3638;
wire n_16084;
wire n_214;
wire n_31196;
wire n_20350;
wire FE_RN_339_0;
wire n_43556;
wire n_13079;
wire n_13577;
wire n_18859;
wire n_5575;
wire newNet_1673;
wire n_3147;
wire n_3556;
wire n_26851;
wire n_23833;
wire FE_OCP_RBN2829_n_30731;
wire n_38807;
wire n_43374;
wire newNet_1560;
wire n_12270;
wire n_850;
wire n_32765;
wire delay_add_ln22_unr5_stage3_stallmux_q_9_;
wire newNet_263;
wire n_21253;
wire n_23748;
wire FE_OCP_RBN3798_delay_xor_ln22_unr12_stage5_stallmux_q_0_;
wire n_15939;
wire n_42505;
wire delay_xor_ln21_unr18_stage7_stallmux_q_10_;
wire n_20372;
wire n_805;
wire n_14827;
wire beta_19;
wire newNet_3599;
wire n_12409;
wire n_12653;
wire n_35769;
wire n_40166;
wire n_40198;
wire FE_OCP_RBN2750_n_9629;
wire n_32417;
wire n_27095;
wire n_11294;
wire n_18874;
wire newNet_793;
wire n_41968;
wire n_17318;
wire newNet_3512;
wire delay_add_ln22_unr17_stage7_stallmux_q_3_;
wire n_35378;
wire n_2060;
wire n_2655;
wire FE_RN_690_0;
wire n_32100;
wire n_36889;
wire n_6015;
wire n_18459;
wire n_35436;
wire n_23944;
wire n_26868;
wire newNet_2922;
wire n_18472;
wire newNet_3005;
wire n_43768;
wire n_23512;
wire n_7389;
wire n_6667;
wire n_4538;
wire n_4265;
wire FE_OCP_RBN1369_n_20763;
wire newNet_685;
wire n_16010;
wire n_29855;
wire n_12804;
wire n_27823;
wire n_5986;
wire n_7662;
wire FE_RN_1608_0;
wire n_32539;
wire newNet_2161;
wire n_5168;
wire n_55;
wire n_31937;
wire FE_RN_1363_0;
wire n_33581;
wire n_40228;
wire n_38093;
wire n_38451;
wire n_28024;
wire n_5720;
wire n_7306;
wire n_36752;
wire n_19790;
wire n_2871;
wire n_13474;
wire n_7188;
wire n_12402;
wire FE_RN_119_0;
wire n_40028;
wire n_16755;
wire n_32773;
wire n_5522;
wire n_30150;
wire n_17715;
wire n_16322;
wire newNet_641;
wire FE_RN_329_0;
wire n_38797;
wire n_19218;
wire n_36470;
wire n_35612;
wire n_24234;
wire n_13547;
wire n_4875;
wire n_9571;
wire n_31577;
wire n_13540;
wire n_44516;
wire FE_RN_1300_0;
wire n_11864;
wire n_19006;
wire n_8760;
wire n_29671;
wire n_20516;
wire n_2232;
wire n_29649;
wire n_22721;
wire n_11987;
wire n_31377;
wire n_29461;
wire n_46987;
wire n_21282;
wire n_19314;
wire FE_OCP_RBN3610_FE_OCPN1797_n_20333;
wire n_27619;
wire n_34918;
wire n_38684;
wire n_42296;
wire FE_OCP_RBN3605_n_8981;
wire n_22790;
wire newNet_1618;
wire n_46220;
wire n_25003;
wire n_26571;
wire n_16612;
wire n_544;
wire newNet_750;
wire n_11025;
wire n_35257;
wire n_5253;
wire n_22847;
wire n_20047;
wire n_26073;
wire n_34322;
wire n_12995;
wire n_24513;
wire FE_OCP_RBN2995_n_35539;
wire delay_xor_ln21_unr21_stage8_stallmux_q_8_;
wire n_43813;
wire n_34491;
wire n_19641;
wire FE_RN_29_0;
wire FE_OCP_RBN1216_n_20595;
wire n_14172;
wire newNet_1807;
wire n_24102;
wire n_1022;
wire FE_OCP_RBN3825_n_18951;
wire n_35508;
wire n_24508;
wire newNet_2242;
wire n_42978;
wire n_32258;
wire n_15930;
wire n_43143;
wire n_32269;
wire n_31372;
wire n_43222;
wire newNet_2744;
wire n_13098;
wire n_39150;
wire n_19362;
wire n_45155;
wire n_19547;
wire n_44819;
wire newNet_1485;
wire n_17392;
wire n_21275;
wire n_43604;
wire n_23397;
wire n_294;
wire n_17298;
wire n_41330;
wire n_29599;
wire n_31485;
wire FE_OCPN953_n_41540;
wire n_11850;
wire delay_xor_ln21_unr3_stage2_stallmux_q_28_;
wire FE_RN_1557_0;
wire FE_RN_362_0;
wire n_7729;
wire n_14808;
wire n_43722;
wire n_12379;
wire n_29308;
wire n_41608;
wire n_33852;
wire n_19011;
wire newNet_1738;
wire n_38458;
wire newNet_1342;
wire delay_xor_ln22_unr21_stage8_stallmux_q_0_;
wire n_30267;
wire n_4492;
wire FE_OCP_RBN3687_n_5105;
wire n_16367;
wire n_20162;
wire n_15753;
wire n_16176;
wire n_30868;
wire n_14669;
wire n_42933;
wire n_29110;
wire n_27273;
wire n_6312;
wire n_35531;
wire n_19872;
wire n_24452;
wire n_8094;
wire n_22709;
wire n_4145;
wire n_34608;
wire n_27538;
wire n_7090;
wire n_36416;
wire n_36547;
wire n_12150;
wire n_6369;
wire n_25447;
wire newNet_528;
wire n_32137;
wire n_2504;
wire n_46353;
wire n_7633;
wire n_2384;
wire n_29491;
wire FE_RN_1606_0;
wire n_37409;
wire n_4908;
wire n_11575;
wire n_16885;
wire n_47007;
wire n_42207;
wire n_27384;
wire FE_OCP_RBN2009_n_45622;
wire n_18912;
wire n_15735;
wire n_7750;
wire n_41222;
wire n_23924;
wire FE_RN_672_0;
wire n_11890;
wire FE_OCPN1527_n_26296;
wire n_36792;
wire n_29300;
wire n_29960;
wire n_40356;
wire n_27531;
wire n_31211;
wire newNet_3472;
wire newNet_2845;
wire n_46187;
wire n_38596;
wire n_39383;
wire n_22117;
wire n_14560;
wire n_27447;
wire n_19672;
wire n_5295;
wire FE_OCP_RBN2167_n_32892;
wire n_23466;
wire n_17256;
wire n_16439;
wire newNet_2877;
wire n_8125;
wire n_19518;
wire n_46141;
wire FE_OCP_RBN1365_n_29444;
wire n_4382;
wire FE_RN_1805_0;
wire n_46251;
wire delay_xor_ln22_unr6_stage3_stallmux_q_18_;
wire n_30416;
wire n_39500;
wire FE_OCP_RBN2533_n_47018;
wire n_7996;
wire n_35547;
wire n_18725;
wire n_29164;
wire n_18816;
wire n_27026;
wire n_1603;
wire n_38261;
wire n_11304;
wire newNet_1051;
wire n_15449;
wire n_38113;
wire n_26468;
wire n_41348;
wire n_25186;
wire n_11599;
wire newNet_3706;
wire newNet_84;
wire n_26125;
wire n_14127;
wire n_16988;
wire n_31438;
wire n_7987;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_31_;
wire newNet_1946;
wire n_39684;
wire n_46211;
wire n_33752;
wire n_986;
wire n_34767;
wire n_12980;
wire newNet_3687;
wire n_2225;
wire newNet_1592;
wire n_7404;
wire n_13862;
wire n_20215;
wire n_20413;
wire n_13801;
wire n_7177;
wire n_38356;
wire n_43064;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_24_;
wire n_28287;
wire n_4122;
wire newNet_2247;
wire FE_RN_278_0;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_1_;
wire n_4222;
wire n_29417;
wire newNet_1663;
wire FE_RN_173_0;
wire n_28198;
wire n_26880;
wire delay_add_ln22_unr27_stage10_stallmux_q_11_;
wire n_35860;
wire n_16673;
wire n_3064;
wire n_28559;
wire n_31423;
wire n_43772;
wire n_24937;
wire n_29224;
wire newNet_1850;
wire n_12620;
wire n_36915;
wire n_25727;
wire n_5979;
wire n_20267;
wire n_14771;
wire n_40883;
wire n_24018;
wire newNet_938;
wire n_33065;
wire n_24471;
wire n_22804;
wire newNet_2393;
wire n_21378;
wire newNet_2199;
wire n_42062;
wire n_16537;
wire n_32375;
wire n_36265;
wire n_19041;
wire n_10633;
wire newNet_277;
wire n_6561;
wire n_9689;
wire n_32518;
wire n_30260;
wire FE_OCP_RBN2188_n_37686;
wire n_15354;
wire n_1743;
wire n_3309;
wire n_9112;
wire n_855;
wire n_9993;
wire delay_add_ln22_unr27_stage10_stallmux_q_31_;
wire n_2104;
wire n_28831;
wire n_609;
wire n_40638;
wire n_40581;
wire n_36123;
wire n_42073;
wire n_38241;
wire n_29333;
wire n_31463;
wire n_29124;
wire n_3857;
wire n_42982;
wire n_31076;
wire n_43731;
wire newNet_2644;
wire n_1570;
wire n_127;
wire n_12141;
wire n_4101;
wire n_35347;
wire FE_OCP_RBN2415_n_8219;
wire n_24968;
wire n_10270;
wire n_41368;
wire n_42680;
wire n_44687;
wire n_43045;
wire n_37421;
wire n_31815;
wire n_21462;
wire newNet_2253;
wire n_11711;
wire n_9083;
wire n_5808;
wire n_21702;
wire FE_RN_1386_0;
wire n_28270;
wire n_33020;
wire n_17545;
wire n_41530;
wire FE_OCP_RBN2530_n_9044;
wire n_10220;
wire n_13223;
wire n_24961;
wire n_2722;
wire n_19424;
wire FE_RN_589_0;
wire newNet_3695;
wire n_19279;
wire n_32113;
wire n_20680;
wire n_20532;
wire n_10614;
wire delay_add_ln22_unr11_stage5_stallmux_q_16_;
wire n_24318;
wire n_38017;
wire n_4844;
wire n_26057;
wire n_12734;
wire n_38334;
wire n_32051;
wire n_20069;
wire newNet_3015;
wire n_491;
wire n_23517;
wire n_6287;
wire n_34989;
wire n_37207;
wire n_11741;
wire n_28077;
wire n_33932;
wire n_25341;
wire n_12600;
wire n_14858;
wire n_42514;
wire n_41476;
wire n_3436;
wire newNet_1001;
wire n_32969;
wire n_15392;
wire n_30908;
wire n_43004;
wire n_35581;
wire n_40616;
wire FE_RN_462_0;
wire n_12027;
wire n_8698;
wire newNet_2287;
wire newNet_2274;
wire n_29626;
wire n_6767;
wire n_8087;
wire FE_OCP_RBN2930_n_5221;
wire n_2594;
wire n_12976;
wire n_32378;
wire FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire n_31725;
wire n_14138;
wire n_26407;
wire n_21825;
wire n_21365;
wire n_20288;
wire n_24929;
wire n_37636;
wire n_31121;
wire n_16569;
wire n_8507;
wire n_40451;
wire n_35316;
wire n_27378;
wire n_43311;
wire newNet_2861;
wire n_31722;
wire newNet_325;
wire n_25115;
wire newNet_565;
wire n_18665;
wire n_3413;
wire n_19104;
wire n_14402;
wire n_4008;
wire FE_RN_404_0;
wire n_19033;
wire FE_RN_485_0;
wire n_31139;
wire n_26162;
wire n_4293;
wire n_21628;
wire n_40938;
wire n_26520;
wire n_18468;
wire n_32638;
wire n_31837;
wire n_39289;
wire n_15598;
wire newNet_587;
wire n_3938;
wire n_19565;
wire n_32399;
wire FE_OCP_RBN3734_n_31819;
wire newNet_469;
wire n_40111;
wire n_21762;
wire n_18497;
wire n_4320;
wire FE_RN_1027_0;
wire FE_OCPN1449_n_20443;
wire delay_xor_ln21_unr3_stage2_stallmux_q_7_;
wire n_24844;
wire n_32054;
wire n_33724;
wire n_16376;
wire n_37079;
wire n_34228;
wire n_24635;
wire n_15410;
wire n_581;
wire FE_RN_1427_0;
wire n_29072;
wire n_27555;
wire n_505;
wire n_40248;
wire n_23824;
wire FE_OCP_RBN3307_n_44722;
wire n_37896;
wire n_11218;
wire n_4026;
wire n_32294;
wire n_30883;
wire n_2898;
wire n_17388;
wire n_39091;
wire n_35424;
wire n_5648;
wire newNet_1856;
wire n_3186;
wire n_5769;
wire n_25370;
wire n_37276;
wire FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_16344;
wire n_30178;
wire n_26113;
wire n_25962;
wire n_35415;
wire n_539;
wire n_42193;
wire newNet_2904;
wire n_32805;
wire n_16171;
wire newNet_3298;
wire n_7426;
wire n_38053;
wire FE_OCP_DRV_N1591_n_34327;
wire FE_OCPN870_n_2737;
wire n_5285;
wire n_17017;
wire n_20095;
wire newNet_679;
wire n_23277;
wire newNet_186;
wire n_21969;
wire FE_OCP_RBN3564_n_29857;
wire n_24899;
wire n_36534;
wire n_18198;
wire n_47261;
wire n_12523;
wire n_33715;
wire FE_OCP_RBN2918_n_16084;
wire n_1447;
wire n_35481;
wire n_25303;
wire n_5637;
wire n_32867;
wire FE_OCP_RBN2726_n_4219;
wire n_7791;
wire n_17310;
wire newNet_861;
wire FE_OCP_RBN3142_n_32395;
wire n_6233;
wire FE_OCPN1397_n_21973;
wire n_10037;
wire FE_OCPN1465_n_13014;
wire n_40037;
wire n_25601;
wire n_22128;
wire newNet_2493;
wire n_24798;
wire n_8497;
wire n_924;
wire n_32926;
wire n_411;
wire n_7998;
wire n_32951;
wire n_36400;
wire n_10773;
wire n_38427;
wire newNet_1716;
wire n_12102;
wire n_17616;
wire n_25066;
wire n_24785;
wire n_30735;
wire n_9924;
wire n_9424;
wire n_30136;
wire n_18059;
wire n_36592;
wire n_9875;
wire n_2853;
wire n_12748;
wire n_15850;
wire n_23225;
wire FE_OCP_RBN2382_n_3502;
wire n_38213;
wire n_39177;
wire n_14018;
wire FE_OCP_RBN2558_n_44576;
wire n_27862;
wire n_2585;
wire n_43908;
wire n_31624;
wire newNet_725;
wire n_15677;
wire n_3579;
wire n_25898;
wire n_24100;
wire n_438;
wire n_40471;
wire n_35294;
wire n_28788;
wire newNet_3463;
wire n_11098;
wire n_5736;
wire newNet_2030;
wire n_33395;
wire newNet_1959;
wire n_3762;
wire n_28778;
wire n_28436;
wire n_3980;
wire n_12500;
wire newNet_1326;
wire n_3717;
wire newNet_2206;
wire FE_OCP_RBN2444_n_42051;
wire n_18088;
wire newNet_3116;
wire FE_OCP_RBN2994_n_35539;
wire n_40777;
wire n_7895;
wire delay_xor_ln21_unr3_stage2_stallmux_q_16_;
wire n_16029;
wire newNet_3621;
wire n_5092;
wire FE_OCP_RBN2141_FE_OCPN861_n_45450;
wire n_36105;
wire n_37871;
wire n_27414;
wire n_7632;
wire FE_RN_1867_0;
wire n_23030;
wire n_11;
wire n_40547;
wire n_43740;
wire n_11759;
wire n_30373;
wire FE_RN_946_0;
wire n_6035;
wire n_15373;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_15_;
wire n_21901;
wire n_10471;
wire n_23331;
wire n_15812;
wire delay_xor_ln22_unr3_stage2_stallmux_q_8_;
wire n_6328;
wire newNet_2082;
wire newNet_422;
wire n_39322;
wire n_37574;
wire n_11631;
wire n_29639;
wire n_1795;
wire n_19922;
wire n_16059;
wire n_10467;
wire n_37494;
wire n_25818;
wire n_22170;
wire n_7848;
wire n_45144;
wire n_15784;
wire n_3661;
wire n_5933;
wire n_26006;
wire n_2759;
wire n_24414;
wire n_1213;
wire n_7235;
wire n_14443;
wire n_13430;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_8_;
wire FE_RN_924_0;
wire n_30974;
wire n_15461;
wire n_24107;
wire n_17841;
wire n_12136;
wire n_13103;
wire n_31630;
wire newNet_28;
wire n_963;
wire n_12514;
wire n_30246;
wire n_6297;
wire FE_OCP_RBN2631_n_29947;
wire FE_OCP_RBN1923_cordic_combinational_sub_ln23_0_unr12_z_0__;
wire FE_OCP_RBN1210_n_16814;
wire n_13492;
wire n_24748;
wire n_328;
wire n_4516;
wire n_46937;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_4_;
wire FE_OCP_RBN1223_n_22914;
wire n_14071;
wire n_5370;
wire n_26791;
wire n_9660;
wire n_24153;
wire n_13902;
wire n_25140;
wire n_252;
wire n_16363;
wire FE_OCP_RBN3282_n_44365;
wire n_19127;
wire n_30499;
wire newNet_12;
wire FE_RN_1372_0;
wire n_648;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_29_;
wire n_6809;
wire n_31666;
wire FE_OCP_RBN2862_n_5024;
wire n_12178;
wire n_1830;
wire FE_RN_309_0;
wire FE_OCP_RBN2980_n_5656;
wire n_23345;
wire n_31742;
wire n_43480;
wire delay_xor_ln21_unr9_stage4_stallmux_q_6_;
wire n_9705;
wire FE_OCP_RBN2610_n_3718;
wire n_15552;
wire n_27652;
wire n_28079;
wire n_30399;
wire newNet_1980;
wire n_31953;
wire n_39221;
wire n_7298;
wire n_20812;
wire n_5064;
wire n_32168;
wire n_10023;
wire n_34451;
wire n_29664;
wire n_3377;
wire n_39984;
wire n_4235;
wire sin_out_25;
wire n_38645;
wire n_7712;
wire beta_11;
wire n_38051;
wire n_2904;
wire n_30306;
wire n_11810;
wire n_15513;
wire n_3040;
wire n_17170;
wire n_23855;
wire n_6330;
wire n_25772;
wire n_14741;
wire n_14615;
wire n_25591;
wire FE_RN_772_0;
wire n_25743;
wire n_33873;
wire n_25869;
wire n_23039;
wire n_19148;
wire newNet_2972;
wire n_39202;
wire n_33296;
wire n_7971;
wire n_41901;
wire FE_OCP_RBN3074_n_43230;
wire n_41314;
wire n_15164;
wire n_7578;
wire n_31877;
wire n_8318;
wire n_41077;
wire n_28653;
wire n_10403;
wire n_15151;
wire n_5321;
wire n_41097;
wire FE_RN_1303_0;
wire n_15949;
wire n_34247;
wire n_13705;
wire n_26220;
wire n_17091;
wire n_12704;
wire n_20928;
wire cos_out_13;
wire n_7203;
wire n_29570;
wire n_45616;
wire n_32489;
wire n_355;
wire newNet_2799;
wire n_38310;
wire n_3276;
wire n_4055;
wire n_42936;
wire n_27031;
wire n_20106;
wire newNet_1883;
wire n_3108;
wire n_22088;
wire n_1369;
wire n_34648;
wire n_29389;
wire n_1982;
wire n_36253;
wire n_1698;
wire FE_RN_1799_0;
wire n_10722;
wire n_18108;
wire n_6371;
wire n_40308;
wire n_1071;
wire delay_xor_ln21_unr18_stage7_stallmux_q_12_;
wire n_6746;
wire delay_add_ln22_unr5_stage3_stallmux_q_28_;
wire n_16471;
wire newNet_3530;
wire n_38569;
wire newNet_2776;
wire n_13244;
wire n_28528;
wire FE_OCP_RBN3576_n_4528;
wire n_4089;
wire n_25849;
wire n_12648;
wire delay_add_ln22_unr17_stage7_stallmux_q_11_;
wire n_7877;
wire n_34704;
wire n_10355;
wire n_24760;
wire n_8471;
wire n_43471;
wire n_30518;
wire newNet_764;
wire newNet_740;
wire n_15609;
wire n_39112;
wire n_32831;
wire newNet_2932;
wire n_41324;
wire n_27521;
wire n_39551;
wire n_30714;
wire n_28730;
wire delay_xor_ln21_unr6_stage3_stallmux_q_19_;
wire n_14836;
wire n_12496;
wire n_38586;
wire n_27752;
wire n_10094;
wire n_17272;
wire n_5071;
wire FE_OCP_RBN1347_n_19270;
wire n_36567;
wire n_7016;
wire newNet_1254;
wire n_21573;
wire n_4066;
wire n_38761;
wire n_34049;
wire newNet_3443;
wire FE_OCP_RBN3486_n_2438;
wire n_5057;
wire n_18583;
wire n_12790;
wire n_9800;
wire n_34138;
wire n_14638;
wire n_39462;
wire n_10835;
wire n_34256;
wire n_20528;
wire n_18184;
wire n_42022;
wire n_20509;
wire n_202;
wire FE_OCP_RBN2958_n_26231;
wire n_16297;
wire n_21088;
wire newNet_1558;
wire newNet_955;
wire n_4379;
wire n_35399;
wire FE_RN_1306_0;
wire n_33929;
wire n_3726;
wire n_21481;
wire n_18041;
wire n_7838;
wire n_28165;
wire n_22054;
wire n_34509;
wire n_13009;
wire n_30615;
wire n_3028;
wire n_43337;
wire n_8580;
wire FE_OCP_RBN3018_n_31117;
wire FE_RN_1286_0;
wire n_378;
wire n_9103;
wire n_29368;
wire n_10219;
wire n_31970;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_3_;
wire newNet_1728;
wire n_11856;
wire n_2558;
wire n_12316;
wire n_20774;
wire n_42996;
wire n_15706;
wire n_20305;
wire FE_RN_1459_0;
wire n_42703;
wire n_18846;
wire n_8528;
wire n_34877;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_6_;
wire delay_add_ln22_unr2_stage2_stallmux_q_10_;
wire n_75;
wire n_12985;
wire n_17228;
wire delay_add_ln22_unr2_stage2_stallmux_q_29_;
wire n_37774;
wire n_18355;
wire n_16332;
wire n_5761;
wire n_41485;
wire n_29408;
wire n_21403;
wire delay_sub_ln21_0_unr20_stage8_stallmux_q_19_;
wire n_43171;
wire n_5750;
wire n_17299;
wire n_38341;
wire n_24007;
wire n_28136;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_13_;
wire n_8269;
wire n_43814;
wire n_14125;
wire n_43429;
wire n_14715;
wire n_20858;
wire n_3250;
wire n_15108;
wire n_36248;
wire n_23733;
wire n_36883;
wire FE_OCP_RBN2350_n_38515;
wire n_36987;
wire n_8353;
wire n_14709;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_21_;
wire delay_sub_ln23_0_unr16_stage6_stallmux_q_29_;
wire newNet_731;
wire n_20577;
wire n_4542;
wire FE_RN_227_0;
wire newNet_3452;
wire n_7196;
wire newNet_3563;
wire n_14817;
wire FE_RN_149_0;
wire n_20851;
wire FE_OCPN1531_n_21790;
wire n_29390;
wire n_15498;
wire n_5081;
wire n_2687;
wire n_32093;
wire n_14881;
wire n_43396;
wire n_28656;
wire newNet_1334;
wire n_43130;
wire n_42429;
wire n_12848;
wire n_1721;
wire FE_OCPN3776_n_43019;
wire n_27720;
wire newNet_433;
wire n_3354;
wire n_249;
wire n_19716;
wire n_15086;
wire n_37461;
wire n_6989;
wire n_29791;
wire n_3741;
wire n_10929;
wire n_13077;
wire n_42418;
wire n_27135;
wire n_19170;
wire newNet_1926;
wire delay_xor_ln21_unr3_stage2_stallmux_q_26_;
wire FE_RN_65_0;
wire n_12693;
wire n_35995;
wire n_29480;
wire n_15665;
wire newNet_1917;
wire n_21322;
wire n_43370;
wire n_10257;
wire n_1232;
wire n_32527;
wire FE_OCP_RBN2813_n_25817;
wire n_40654;
wire n_21428;
wire n_38067;
wire n_35653;
wire n_16553;
wire FE_RN_1008_0;
wire n_42356;
wire n_1228;
wire n_12660;
wire n_28259;
wire n_29684;
wire n_42115;
wire n_34618;
wire n_38119;
wire n_30479;
wire n_26268;
wire n_26666;
wire n_35336;
wire n_13827;
wire n_5854;
wire n_23884;
wire n_42303;
wire n_12212;
wire n_24047;
wire n_16211;
wire n_41514;
wire n_22112;
wire n_31414;
wire n_39612;
wire FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_;
wire n_7613;
wire n_39360;
wire n_42629;
wire n_1055;
wire n_19796;
wire n_28647;
wire n_27487;
wire n_7505;
wire n_19818;
wire n_13795;
wire newNet_271;
wire n_25119;
wire n_27096;
wire n_19530;
wire FE_OCP_RBN2764_n_25732;
wire FE_RN_1494_0;
wire n_25517;
wire n_7590;
wire n_9001;
wire n_15771;
wire n_4247;
wire n_21821;
wire n_18932;
wire newNet_3711;
wire n_2677;
wire n_7937;
wire newNet_2945;
wire n_39768;
wire delay_add_ln22_unr20_stage8_stallmux_q_23_;
wire FE_OCP_RBN2251_n_13017;
wire n_45188;
wire n_16929;
wire n_40954;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_18_;
wire n_10783;
wire newNet_3021;
wire n_19099;
wire FE_OCPN878_n_44734;
wire FE_OCPN847_n_3597;
wire n_31672;
wire n_11463;
wire n_34953;
wire n_25093;
wire n_15338;
wire n_20849;
wire n_45884;
wire n_39181;
wire delay_add_ln22_unr17_stage7_stallmux_q_23_;
wire n_19580;
wire n_17158;
wire n_26002;
wire newNet_1582;
wire n_39335;
wire newNet_2633;
wire n_3449;
wire n_30955;
wire n_39830;
wire n_13115;
wire FE_RN_866_0;
wire n_34849;
wire n_38880;
wire newNet_1532;
wire n_26294;
wire n_15653;
wire n_43587;
wire n_8669;
wire newNet_3409;
wire n_36384;
wire n_38091;
wire FE_OCPN850_n_2306;
wire FE_OCP_RBN1146_n_13098;
wire n_3409;
wire n_4831;
wire n_20426;
wire n_11069;
wire FE_OCP_RBN3015_n_31117;
wire n_28450;
wire n_23227;
wire n_4540;
wire n_36421;
wire n_35845;
wire n_16164;
wire newNet_1063;
wire n_1084;
wire n_11999;
wire n_19708;
wire n_23543;
wire n_15442;
wire n_13711;
wire n_18719;
wire n_30080;
wire n_11400;
wire n_32289;
wire n_22448;
wire n_21855;
wire n_23173;
wire n_37647;
wire n_17867;
wire n_36777;
wire n_19650;
wire n_43686;
wire newNet_2691;
wire n_42492;
wire n_10090;
wire n_3225;
wire n_24852;
wire FE_OCP_RBN3847_FE_RN_1548_0;
wire n_35285;
wire n_9763;
wire delay_xor_ln22_unr6_stage3_stallmux_q_6_;
wire FE_RN_241_0;
wire n_38154;
wire n_2636;
wire n_31572;
wire n_42510;
wire n_4922;
wire n_42721;
wire n_26899;
wire n_13447;
wire n_32248;
wire n_23430;
wire newNet_316;
wire n_8898;
wire n_26747;
wire n_34106;
wire n_27916;
wire n_40493;
wire n_25076;
wire n_22165;
wire n_38882;
wire newNet_922;
wire n_18945;
wire newNet_2704;
wire n_43516;
wire n_41310;
wire n_18433;
wire n_19113;
wire n_24307;
wire n_39635;
wire n_27895;
wire n_17826;
wire n_3495;
wire n_16162;
wire FE_OCP_DRV_N1550_n_19053;
wire n_37584;
wire n_23684;
wire n_269;
wire n_31057;
wire n_29135;
wire n_7387;
wire n_12477;
wire n_24216;
wire n_23423;
wire n_7566;
wire n_4709;
wire n_445;
wire n_43054;
wire n_38776;
wire n_11730;
wire n_35947;
wire n_16725;
wire n_23879;
wire n_16727;
wire FE_OCP_RBN2459_n_13765;
wire n_34147;
wire n_29016;
wire FE_OCP_DRV_N3147_n_33225;
wire n_30357;
wire n_35350;
wire newNet_2513;
wire newNet_1695;
wire n_6874;
wire n_22366;
wire n_20936;
wire n_42341;
wire n_11678;
wire n_12185;
wire n_34061;
wire n_24116;
wire n_18235;
wire newNet_1872;
wire n_8688;
wire n_37255;
wire n_17495;
wire newNet_543;
wire n_44659;
wire n_40120;
wire FE_OCP_DRV_N1561_n_19562;
wire n_24768;
wire n_8229;
wire newNet_2483;
wire FE_RN_1759_0;
wire n_16944;
wire newNet_902;
wire n_7449;
wire n_5026;
wire newNet_598;
wire FE_OCP_RBN2336_n_8269;
wire newNet_49;
wire delay_add_ln22_unr20_stage8_stallmux_q_19_;
wire n_29745;
wire n_22198;
wire FE_RN_20_0;
wire n_29271;
wire n_42654;
wire n_21466;
wire n_23777;
wire n_16228;
wire n_25636;
wire newNet_1031;
wire FE_OCP_RBN3458_n_33872;
wire n_21638;
wire n_46203;
wire n_32625;
wire n_25812;
wire n_9127;
wire n_36544;
wire n_1144;
wire n_17483;
wire n_43304;
wire delay_xor_ln22_unr3_stage2_stallmux_q_19_;
wire newNet_1055;
wire n_30739;
wire n_16464;
wire n_1088;
wire newNet_2227;
wire n_8153;
wire FE_OCP_DRV_N1612_n_21706;
wire n_34566;
wire n_21743;
wire n_39892;
wire n_18889;
wire n_30180;
wire n_8513;
wire n_32748;
wire FE_OCP_RBN3014_n_31117;
wire n_28464;
wire FE_RN_1510_0;
wire n_42778;
wire n_15920;
wire newNet_2824;
wire n_12929;
wire FE_OCP_RBN2341_n_29470;
wire n_43578;
wire FE_OCP_RBN2854_n_45462;
wire beta_3;
wire n_25455;
wire n_18540;
wire n_18488;
wire n_40104;
wire n_34031;
wire n_18115;
wire n_30611;
wire n_36683;
wire n_42107;
wire FE_OCP_RBN1989_delay_xor_ln23_unr6_stage3_stallmux_q;
wire n_7932;
wire n_11359;
wire n_10156;
wire n_35619;
wire n_7817;
wire n_13385;
wire n_10313;
wire n_12389;
wire n_38326;
wire n_41996;
wire newNet_3257;
wire beta_31;
wire FE_OCP_RBN1145_n_13098;
wire n_21120;
wire n_22258;
wire n_40157;
wire n_28988;
wire n_20038;
wire newNet_3572;
wire n_39992;
wire n_13334;
wire FE_RN_1593_0;
wire newNet_2833;
wire n_41423;
wire n_40913;
wire FE_RN_1735_0;
wire FE_RN_1243_0;
wire n_39555;
wire n_14982;
wire n_34658;
wire n_34026;
wire n_1194;
wire n_41963;
wire n_37312;
wire n_24408;
wire n_20219;
wire n_42840;
wire n_40800;
wire FE_OCP_RBN3481_n_13667;
wire n_41695;
wire n_37150;
wire n_37129;
wire n_41744;
wire delay_xor_ln21_unr9_stage4_stallmux_q_21_;
wire n_14582;
wire n_15149;
wire n_1518;
wire n_40222;
wire n_35787;
wire n_32426;
wire n_16910;
wire n_8362;
wire n_28510;
wire FE_RN_1698_0;
wire n_11426;
wire newNet_1373;
wire n_14790;
wire n_29317;
wire newNet_1892;
wire newNet_2485;
wire n_2566;
wire n_34843;
wire n_37428;
wire newNet_963;
wire n_15889;
wire n_271;
wire n_17549;
wire n_28245;
wire newNet_701;
wire n_34808;
wire n_41736;
wire newNet_1312;
wire n_11095;
wire n_1654;
wire n_5204;
wire n_15819;
wire n_34715;
wire n_6209;
wire n_10387;
wire n_37366;
wire n_36392;
wire n_5948;
wire n_23790;
wire delay_xor_ln21_unr9_stage4_stallmux_q_14_;
wire n_19808;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_20_;
wire n_24393;
wire n_29523;
wire n_30751;
wire n_4656;
wire n_1291;
wire n_33831;
wire newNet_3745;
wire n_42119;
wire n_29430;
wire n_14288;
wire n_31253;
wire n_23891;
wire n_9213;
wire n_42616;
wire FE_OCP_RBN2932_n_5307;
wire newNet_1789;
wire n_18634;
wire n_5154;
wire n_9717;
wire FE_OFN790_n_8981;
wire n_1589;
wire delay_add_ln22_unr14_stage6_stallmux_q_29_;
wire newNet_2898;
wire n_7658;
wire n_8267;
wire n_3286;
wire n_16984;
wire n_39026;
wire FE_OCP_RBN3377_n_1675;
wire n_46193;
wire n_6456;
wire FE_RN_209_0;
wire n_402;
wire n_2428;
wire n_37814;
wire FE_OFN27_n_1142;
wire FE_RN_1559_0;
wire n_41001;
wire cos_out_9;
wire n_6383;
wire n_26766;
wire n_15186;
wire n_21344;
wire n_23958;
wire n_33549;
wire n_516;
wire FE_OCP_RBN2746_n_47011;
wire n_23987;
wire FE_OCP_DRV_N3152_n_13264;
wire n_10518;
wire n_30072;
wire n_3650;
wire n_17510;
wire n_858;
wire n_44296;
wire n_37332;
wire n_35325;
wire n_33792;
wire n_14261;
wire FE_OCP_RBN2986_n_35539;
wire n_22308;
wire n_43388;
wire n_23806;
wire n_39758;
wire n_29439;
wire n_14077;
wire n_41574;
wire newNet_1815;
wire n_30605;
wire n_14110;
wire n_2611;
wire newNet_2230;
wire n_14191;
wire n_33115;
wire n_33662;
wire n_4591;
wire n_21971;
wire n_35806;
wire newNet_493;
wire n_230;
wire n_2523;
wire n_39803;
wire n_5864;
wire n_9621;
wire n_12765;
wire n_11815;
wire n_13695;
wire n_34088;
wire n_18565;
wire n_12864;
wire newNet_844;
wire n_10391;
wire n_12883;
wire n_44213;
wire n_36756;
wire newNet_583;
wire n_1556;
wire FE_RN_883_0;
wire n_21946;
wire n_31491;
wire n_24191;
wire n_3160;
wire n_27833;
wire FE_RN_1017_0;
wire n_9541;
wire n_37201;
wire n_37064;
wire n_1495;
wire n_9965;
wire FE_OCP_RBN3110_n_43711;
wire n_26590;
wire n_43661;
wire n_37092;
wire n_7514;
wire FE_OCP_RBN2851_n_46982;
wire n_33648;
wire n_11961;
wire n_45514;
wire n_4144;
wire n_40448;
wire n_22522;
wire n_23554;
wire n_4861;
wire n_21958;
wire n_26739;
wire newNet_3170;
wire n_42305;
wire newNet_3133;
wire n_26425;
wire n_29109;
wire n_27910;
wire n_23787;
wire n_25286;
wire n_36102;
wire n_31752;
wire n_1952;
wire n_19496;
wire n_16354;
wire n_45533;
wire n_38872;
wire n_5471;
wire n_3538;
wire FE_OCPN1750_n_27223;
wire n_22824;
wire n_25629;
wire n_1165;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_3_;
wire n_24480;
wire newNet_212;
wire FE_RN_1812_0;
wire newNet_2163;
wire n_40405;
wire delay_xor_ln21_unr6_stage3_stallmux_q_13_;
wire n_36574;
wire n_43446;
wire n_6801;
wire n_47212;
wire n_7969;
wire n_46375;
wire n_4880;
wire n_41126;
wire sin_out_3;
wire newNet_744;
wire n_33018;
wire n_24497;
wire n_17238;
wire n_29654;
wire n_15649;
wire n_17376;
wire n_31299;
wire n_9155;
wire n_18750;
wire n_15960;
wire n_42632;
wire n_19766;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_2_;
wire n_32059;
wire n_40421;
wire newNet_3254;
wire n_21554;
wire n_41009;
wire FE_OCP_RBN3511_n_19599;
wire newNet_3597;
wire n_19523;
wire n_26337;
wire n_19821;
wire n_21338;
wire n_7407;
wire n_5423;
wire n_23541;
wire newNet_3721;
wire n_12037;
wire n_18242;
wire n_27121;
wire newNet_3635;
wire newNet_1298;
wire newNet_2728;
wire FE_OCPN3175_n_31125;
wire newNet_3292;
wire n_19323;
wire n_1595;
wire n_4889;
wire n_37688;
wire n_5966;
wire n_34853;
wire n_12611;
wire n_13423;
wire n_24449;
wire n_26944;
wire n_32310;
wire n_17566;
wire n_13672;
wire newNet_440;
wire n_12581;
wire n_22885;
wire n_21053;
wire n_4034;
wire n_34367;
wire n_29550;
wire n_5344;
wire n_36377;
wire n_13185;
wire n_26175;
wire n_31981;
wire n_16482;
wire n_30276;
wire n_31269;
wire newNet_2929;
wire n_41190;
wire n_41199;
wire n_37291;
wire n_5433;
wire n_25685;
wire delay_add_ln22_unr11_stage5_stallmux_q_29_;
wire n_6379;
wire n_40550;
wire n_2438;
wire n_4942;
wire n_17834;
wire n_4044;
wire n_23270;
wire n_42710;
wire n_34278;
wire n_16816;
wire n_23818;
wire n_28703;
wire n_14528;
wire n_12799;
wire n_23815;
wire n_8764;
wire n_13020;
wire n_24467;
wire FE_OCP_RBN2179_FE_RN_526_0;
wire n_12939;
wire FE_OCP_RBN2502_n_13896;
wire FE_OCPN1783_n_26801;
wire n_189;
wire n_18837;
wire n_41804;
wire n_19970;
wire n_36706;
wire n_25670;
wire n_15336;
wire n_21598;
wire n_46965;
wire n_15381;
wire FE_RN_867_0;
wire n_42096;
wire n_42227;
wire n_3489;
wire n_14909;
wire n_37742;
wire n_41970;
wire n_16839;
wire n_19895;
wire n_16304;
wire n_13876;
wire n_39524;
wire n_38206;
wire newNet_2457;
wire n_5117;
wire n_39686;
wire n_1779;
wire FE_RN_692_0;
wire FE_OCP_RBN1992_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_;
wire n_25401;
wire n_23449;
wire n_5464;
wire n_35430;
wire n_4201;
wire n_15303;
wire n_42212;
wire n_17343;
wire n_19072;
wire n_30007;
wire n_39717;
wire newNet_1886;
wire FE_OCP_RBN2662_n_20333;
wire n_21695;
wire n_5516;
wire n_27279;
wire n_25744;
wire n_13853;
wire n_42162;
wire n_41329;
wire n_34497;
wire n_30670;
wire n_28006;
wire n_42181;
wire newNet_789;
wire n_11829;
wire n_3902;
wire n_41797;
wire n_2749;
wire n_13043;
wire n_5331;
wire n_34282;
wire n_42878;
wire n_8250;
wire n_7881;
wire FE_RN_1390_0;
wire n_22690;
wire newNet_3419;
wire n_21983;
wire n_21734;
wire n_300;
wire n_28140;
wire n_20611;
wire n_4767;
wire n_45070;
wire n_29584;
wire n_36222;
wire n_32081;
wire n_5367;
wire n_39469;
wire n_43544;
wire n_32408;
wire n_11481;
wire n_3757;
wire n_29630;
wire n_42265;
wire n_32250;
wire FE_RN_1345_0;
wire n_28921;
wire n_19416;
wire n_19713;
wire n_44723;
wire n_12711;
wire newNet_1495;
wire n_21307;
wire n_17368;
wire FE_RN_614_0;
wire n_16662;
wire n_19555;
wire n_5730;
wire n_17006;
wire n_8942;
wire n_39345;
wire n_30076;
wire n_2134;
wire n_30765;
wire n_43611;
wire n_34104;
wire n_18867;
wire n_35456;
wire n_16683;
wire n_8868;
wire n_41298;
wire FE_RN_1236_0;
wire n_29374;
wire n_4740;
wire n_29446;
wire newNet_1941;
wire n_2241;
wire n_8717;
wire FE_OCPN3757_n_13889;
wire newNet_1507;
wire n_8601;
wire n_16574;
wire n_4521;
wire n_21642;
wire FE_OCP_RBN3137_n_32380;
wire n_5788;
wire n_23990;
wire FE_OCP_RBN3828_n_19204;
wire n_23720;
wire newNet_1160;
wire n_17721;
wire n_13807;
wire n_38671;
wire FE_OCP_RBN3339_n_44610;
wire n_24636;
wire newNet_781;
wire n_7769;
wire n_22344;
wire FE_RN_976_0;
wire n_16405;
wire n_30835;
wire n_9458;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_20_;
wire newNet_1071;
wire n_24703;
wire newNet_2149;
wire n_30729;
wire n_35010;
wire n_19151;
wire n_4847;
wire n_6586;
wire n_146;
wire n_26818;
wire n_364;
wire n_32178;
wire newNet_2315;
wire n_22377;
wire n_45137;
wire n_17937;
wire newNet_3698;
wire n_10766;
wire n_8252;
wire FE_RN_815_0;
wire n_3005;
wire n_35244;
wire n_24011;
wire newNet_1236;
wire FE_RN_152_0;
wire newNet_1574;
wire n_41107;
wire n_16781;
wire n_9419;
wire FE_OCP_RBN1374_n_35275;
wire n_23333;
wire n_41268;
wire n_43757;
wire n_2077;
wire n_27677;
wire n_46229;
wire n_28514;
wire n_3643;
wire n_4335;
wire FE_RN_14_0;
wire n_43875;
wire n_24690;
wire n_11110;
wire n_28838;
wire FE_OCP_RBN1335_n_20941;
wire n_15299;
wire newNet_2873;
wire n_2974;
wire n_24035;
wire n_40780;
wire n_29928;
wire n_14154;
wire n_1862;
wire n_3242;
wire n_12488;
wire n_38235;
wire FE_OCP_RBN3409_n_45120;
wire n_20176;
wire n_28853;
wire n_14490;
wire n_27713;
wire n_9944;
wire n_31228;
wire n_33463;
wire n_17072;
wire n_1111;
wire delay_xor_ln22_unr9_stage4_stallmux_q_11_;
wire n_24695;
wire newNet_656;
wire n_41919;
wire n_35280;
wire n_15973;
wire n_19054;
wire newNet_1539;
wire n_3817;
wire newNet_1148;
wire n_6840;
wire n_41648;
wire n_1477;
wire n_23235;
wire n_27763;
wire newNet_1996;
wire n_23866;
wire n_15642;
wire n_30279;
wire n_21019;
wire n_14726;
wire n_22930;
wire n_2643;
wire n_3305;
wire n_42816;
wire FE_RN_849_0;
wire n_30255;
wire n_26647;
wire n_31799;
wire n_19935;
wire n_44056;
wire FE_RN_783_0;
wire n_18169;
wire FE_RN_1242_0;
wire n_18710;
wire n_29544;
wire n_6907;
wire n_29569;
wire n_18507;
wire n_29693;
wire FE_OCPN1248_n_44267;
wire n_30505;
wire n_40235;
wire n_31968;
wire n_16289;
wire n_9378;
wire n_43855;
wire newNet_1741;
wire n_29660;
wire n_8959;
wire n_19666;
wire n_19572;
wire n_10893;
wire n_40168;
wire n_22868;
wire n_10851;
wire n_32402;
wire n_42459;
wire n_22566;
wire n_24896;
wire n_13953;
wire n_12852;
wire n_20868;
wire FE_RN_937_0;
wire FE_RN_1119_0;
wire FE_OCPN1036_n_28288;
wire n_29141;
wire n_19837;
wire n_34839;
wire n_16807;
wire n_27157;
wire n_36025;
wire n_16188;
wire n_30541;
wire n_22631;
wire n_7462;
wire n_22494;
wire n_36313;
wire n_41723;
wire n_37054;
wire n_42649;
wire n_40370;
wire n_14996;
wire n_43104;
wire n_38072;
wire n_25209;
wire n_16605;
wire n_19181;
wire n_10317;
wire n_16099;
wire n_34388;
wire FE_OFN774_n_46137;
wire n_33224;
wire n_23648;
wire n_22677;
wire n_17756;
wire n_43258;
wire n_43851;
wire FE_RN_1103_0;
wire n_43369;
wire n_20907;
wire n_42007;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_28_;
wire n_18510;
wire n_30946;
wire n_43178;
wire FE_OCP_RBN2364_n_24372;
wire n_94;
wire n_41978;
wire n_22012;
wire n_9090;
wire n_22291;
wire FE_OCPN1507_n_23414;
wire n_12743;
wire newNet_311;
wire n_41283;
wire n_28749;
wire n_1311;
wire n_9829;
wire FE_RN_1804_0;
wire newNet_3039;
wire n_11303;
wire n_12560;
wire n_30493;
wire FE_RN_1115_0;
wire n_41672;
wire n_38651;
wire n_2508;
wire n_11750;
wire n_26958;
wire newNet_3141;
wire FE_OCP_RBN3832_n_19204;
wire n_39774;
wire FE_RN_360_0;
wire n_4019;
wire n_35647;
wire n_8548;
wire n_39214;
wire n_31851;
wire n_22084;
wire n_19733;
wire n_6616;
wire n_38274;
wire n_7535;
wire n_37480;
wire n_3880;
wire n_40043;
wire n_41130;
wire n_28963;
wire n_30235;
wire n_37803;
wire n_9869;
wire n_33489;
wire FE_OCP_RBN3686_n_16074;
wire n_13352;
wire n_29080;
wire n_2298;
wire FE_OCP_RBN2149_FE_OCPN861_n_45450;
wire FE_OCP_RBN2657_FE_RN_1288_0;
wire n_14020;
wire n_42909;
wire n_43;
wire n_14467;
wire n_27748;
wire n_17639;
wire n_33503;
wire n_21815;
wire n_26117;
wire n_1940;
wire FE_RN_1469_0;
wire n_33755;
wire n_18528;
wire newNet_3360;
wire n_6085;
wire n_36359;
wire n_32017;
wire n_14435;
wire n_36319;
wire newNet_2527;
wire newNet_3371;
wire n_7901;
wire n_29716;
wire n_7070;
wire FE_OFN361_n_9391;
wire n_14698;
wire n_30302;
wire n_47020;
wire n_18347;
wire FE_OCP_RBN1716_n_20734;
wire n_40332;
wire n_28571;
wire n_41401;
wire n_873;
wire n_1306;
wire n_34395;
wire n_31077;
wire n_163;
wire n_15793;
wire newNet_1278;
wire n_27421;
wire n_34127;
wire n_39455;
wire n_23556;
wire newNet_2655;
wire n_468;
wire FE_RN_25_0;
wire n_1050;
wire n_44853;
wire n_29429;
wire n_2222;
wire n_27466;
wire n_7992;
wire n_37635;
wire delay_xor_ln21_unr12_stage5_stallmux_q_14_;
wire n_18666;
wire n_18990;
wire n_38576;
wire FE_RN_678_0;
wire n_30320;
wire newNet_1462;
wire FE_RN_23_0;
wire n_35604;
wire n_34549;
wire n_18700;
wire n_8815;
wire n_22758;
wire newNet_1210;
wire n_38026;
wire n_38348;
wire n_17645;
wire n_24779;
wire n_31142;
wire n_8487;
wire n_13094;
wire n_2007;
wire n_10754;
wire n_42104;
wire n_34603;
wire newNet_196;
wire n_34613;
wire n_11252;
wire n_10042;
wire n_24208;
wire n_25043;
wire newNet_2072;
wire FE_OCP_RBN2741_n_15206;
wire delay_add_ln22_unr20_stage8_stallmux_q_9_;
wire n_11476;
wire FE_OCP_RBN2906_n_16230;
wire newNet_2740;
wire newNet_1218;
wire n_18038;
wire n_8036;
wire n_5849;
wire n_283;
wire n_697;
wire n_43147;
wire n_29512;
wire n_35520;
wire n_39671;
wire FE_OCPN3788_n_15708;
wire n_16443;
wire n_18785;
wire n_28547;
wire FE_RN_349_0;
wire FE_OCP_DRV_N1539_n_35427;
wire n_30747;
wire n_43896;
wire n_20043;
wire n_6186;
wire n_15826;
wire n_6512;
wire n_18316;
wire n_20007;
wire n_14183;
wire n_16912;
wire n_18033;
wire FE_RN_930_0;
wire n_12598;
wire n_37214;
wire n_38608;
wire n_7496;
wire newNet_699;
wire delay_sub_ln23_0_unr29_stage10_stallmux_q;
wire n_32844;
wire newNet_1492;
wire FE_OCP_RBN2130_n_32647;
wire FE_RN_1846_0;
wire n_28753;
wire n_2341;
wire n_41550;
wire n_9569;
wire n_23715;
wire n_39068;
wire n_39954;
wire n_32360;
wire FE_OCP_RBN2981_n_26591;
wire n_4416;
wire n_37436;
wire n_14673;
wire newNet_3156;
wire n_9070;
wire n_10943;
wire delay_sub_ln21_0_unr8_stage4_stallmux_q_9_;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_29_;
wire n_38359;
wire n_40681;
wire n_36442;
wire n_1473;
wire n_34233;
wire n_46417;
wire n_12350;
wire newNet_2297;
wire newNet_458;
wire n_42368;
wire n_11222;
wire n_37622;
wire n_5826;
wire n_23694;
wire n_118;
wire n_27107;
wire n_25470;
wire n_14222;
wire FE_OCPN1432_n_29504;
wire n_12019;
wire n_26351;
wire n_12911;
wire n_2951;
wire n_4114;
wire n_39314;
wire n_22841;
wire n_18920;
wire n_17120;
wire n_8795;
wire n_23620;
wire n_13624;
wire n_489;
wire delay_add_ln22_unr8_stage4_stallmux_q_21_;
wire n_4501;
wire n_6054;
wire n_19207;
wire newNet_616;
wire n_5076;
wire n_19566;
wire n_4077;
wire newNet_6;
wire n_9034;
wire n_35516;
wire n_26234;
wire n_29829;
wire n_21580;
wire n_18264;
wire n_4774;
wire n_5680;
wire FE_OCP_RBN3425_n_44881;
wire n_14497;
wire n_21591;
wire n_37848;
wire n_17803;
wire n_7940;
wire delay_add_ln22_unr5_stage3_stallmux_q_17_;
wire n_11503;
wire FE_OCP_RBN1706_n_20616;
wire n_2621;
wire n_1665;
wire newNet_2401;
wire n_11923;
wire newNet_475;
wire n_33057;
wire n_32893;
wire n_4329;
wire n_33872;
wire FE_OCP_RBN2629_n_14590;
wire n_29851;
wire n_40528;
wire n_31061;
wire n_42580;
wire n_24750;
wire n_36624;
wire n_28152;
wire n_28771;
wire n_25060;
wire n_15178;
wire n_24919;
wire FE_RN_1321_0;
wire n_27234;
wire n_19082;
wire n_32761;
wire n_23187;
wire n_9145;
wire n_25580;
wire n_22107;
wire delay_xor_ln22_unr12_stage5_stallmux_q_11_;
wire n_32577;
wire n_1403;
wire FE_RN_1673_0;
wire FE_RN_1806_0;
wire delay_xor_ln22_unr6_stage3_stallmux_q_4_;
wire n_42684;
wire n_25586;
wire n_37765;
wire n_29764;
wire n_25059;
wire n_29723;
wire n_8730;
wire n_39421;
wire n_9847;
wire n_40010;
wire n_43833;
wire n_39484;
wire n_32026;
wire n_20801;
wire FE_OCP_RBN3838_n_19513;
wire n_18390;
wire n_31390;
wire n_39712;
wire n_27130;
wire newNet_1136;
wire n_28945;
wire n_1132;
wire n_7557;
wire n_242;
wire n_30978;
wire n_2020;
wire n_4601;
wire n_41232;
wire n_29002;
wire n_31783;
wire n_30722;
wire n_4350;
wire n_20672;
wire FE_OCP_RBN1708_n_22150;
wire n_28112;
wire newNet_2257;
wire n_39412;
wire n_42374;
wire n_33825;
wire newNet_3230;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_27_;
wire n_17384;
wire n_36262;
wire delay_add_ln22_unr27_stage10_stallmux_q_30_;
wire newNet_2736;
wire n_22005;
wire n_14646;
wire FE_RN_738_0;
wire n_7432;
wire n_36280;
wire n_28909;
wire n_20548;
wire newNet_2320;
wire n_20401;
wire n_15252;
wire n_15074;
wire n_33256;
wire n_24550;
wire n_12029;
wire n_25192;
wire n_35587;
wire newNet_839;
wire n_5669;
wire n_23079;
wire n_18999;
wire n_45685;
wire n_35000;
wire n_5356;
wire delay_add_ln22_unr23_stage9_stallmux_q_7_;
wire n_37712;
wire n_4429;
wire n_35793;
wire n_40705;
wire n_36179;
wire n_28542;
wire n_19136;
wire n_26486;
wire FE_OCPN1749_n_27223;
wire n_29779;
wire newNet_403;
wire n_31683;
wire n_20081;
wire n_28939;
wire newNet_535;
wire n_23042;
wire n_2735;
wire n_38437;
wire n_35156;
wire n_29734;
wire newNet_663;
wire n_5505;
wire n_13214;
wire n_11561;
wire n_32634;
wire n_16131;
wire n_36294;
wire n_938;
wire n_36928;
wire n_10274;
wire n_35107;
wire n_6625;
wire n_12669;
wire n_34760;
wire n_41379;
wire n_23353;
wire n_29212;
wire n_6851;
wire n_33896;
wire n_22590;
wire n_29349;
wire n_16067;
wire n_23379;
wire n_18882;
wire n_23530;
wire newNet_684;
wire n_38572;
wire n_38743;
wire n_6319;
wire delay_add_ln22_unr5_stage3_stallmux_q_31_;
wire n_2285;
wire n_35033;
wire FE_OCP_RBN3697_n_35543;
wire n_40136;
wire n_35961;
wire n_22853;
wire FE_OCP_RBN3835_n_19241;
wire n_21039;
wire n_39382;
wire n_29477;
wire delay_add_ln22_unr20_stage8_stallmux_q_12_;
wire FE_OCP_RBN2669_n_4158;
wire n_10520;
wire n_2499;
wire n_584;
wire n_35561;
wire newNet_2427;
wire newNet_3676;
wire n_39792;
wire newNet_1269;
wire n_37730;
wire FE_OFN805_n_46196;
wire n_22983;
wire n_40720;
wire n_39290;
wire FE_RN_140_0;
wire n_1577;
wire n_1244;
wire n_41227;
wire n_16020;
wire n_39451;
wire n_14886;
wire n_27901;
wire n_17905;
wire FE_RN_981_0;
wire n_11788;
wire newNet_374;
wire n_2870;
wire n_15450;
wire n_30828;
wire n_3854;
wire n_14399;
wire n_44277;
wire n_22844;
wire n_31346;
wire delay_add_ln22_unr14_stage6_stallmux_q_18_;
wire n_42422;
wire n_28060;
wire newNet_2837;
wire n_32243;
wire n_31073;
wire n_21501;
wire n_34797;
wire n_3833;
wire n_10668;
wire n_39724;
wire n_37058;
wire FE_OCP_RBN3531_n_13765;
wire n_11326;
wire n_8516;
wire n_5498;
wire n_23307;
wire n_23844;
wire n_32350;
wire n_14987;
wire n_6552;
wire n_511;
wire newNet_3694;
wire n_28672;
wire n_24873;
wire n_20488;
wire n_28968;
wire n_46381;
wire n_34825;
wire n_11846;
wire n_42497;
wire n_19436;
wire n_2032;
wire n_42156;
wire n_35493;
wire n_33816;
wire newNet_158;
wire n_14545;
wire n_42905;
wire n_46351;
wire FE_RN_56_0;
wire n_16325;
wire n_33779;
wire n_29880;
wire n_31633;
wire n_853;
wire n_7308;
wire n_1748;
wire n_16634;
wire n_2551;
wire n_33121;
wire n_16590;
wire n_360;
wire n_40670;
wire n_31273;
wire n_29420;
wire n_26980;
wire n_27342;
wire newNet_625;
wire n_25047;
wire n_12503;
wire n_44563;
wire n_4531;
wire newNet_1547;
wire n_42855;
wire n_8884;
wire n_39583;
wire n_34325;
wire FE_RN_167_0;
wire n_37102;
wire n_27100;
wire n_13741;
wire n_39474;
wire n_11378;
wire n_32706;
wire n_35094;
wire n_26625;
wire n_37033;
wire n_20781;
wire n_42241;
wire newNet_1229;
wire n_39226;
wire FE_OCP_RBN2953_n_21538;
wire n_20648;
wire n_41796;
wire newNet_2243;
wire n_25031;
wire n_12112;
wire n_37790;
wire n_4533;
wire n_11507;
wire n_9722;
wire n_34399;
wire n_24577;
wire newNet_461;
wire FE_OCP_RBN2187_n_37686;
wire n_9066;
wire n_12999;
wire n_19686;
wire n_20910;
wire n_1981;
wire n_6091;
wire n_39628;
wire n_23797;
wire FE_OCP_RBN3242_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_;
wire n_20367;
wire newNet_1521;
wire n_20679;
wire n_3282;
wire n_22063;
wire n_28775;
wire n_24039;
wire n_18223;
wire n_28401;
wire n_15488;
wire n_5840;
wire n_43880;
wire n_14005;
wire FE_OCP_RBN2180_FE_RN_526_0;
wire n_3933;
wire n_19398;
wire newNet_1563;
wire n_39607;
wire n_27722;
wire n_2434;
wire n_7423;
wire n_8704;
wire n_34267;
wire n_29489;
wire n_10414;
wire n_1782;
wire newNet_1128;
wire FE_RN_1323_0;
wire n_3323;
wire n_13208;
wire n_9878;
wire n_15613;
wire n_30639;
wire n_23564;
wire n_9294;
wire n_41311;
wire n_22269;
wire n_34123;
wire n_33190;
wire n_4845;
wire n_19702;
wire FE_RN_305_0;
wire n_1706;
wire n_35215;
wire n_43286;
wire n_25101;
wire FE_OCP_DRV_N1567_n_19751;
wire FE_RN_1552_0;
wire FE_OCP_RBN1721_n_21004;
wire n_36270;
wire mux_while_ln12_psv_q_7_;
wire n_8568;
wire newNet_367;
wire delay_sub_ln23_0_unr26_stage9_stallmux_q_1_;
wire n_39147;
wire n_3173;
wire n_19884;
wire n_8336;
wire n_40310;
wire n_41756;
wire n_39840;
wire n_14873;
wire n_35706;
wire delay_sub_ln22_unr24_stage9_stallmux_q_4_;
wire n_23289;
wire n_39865;
wire n_26228;
wire n_10874;
wire n_11407;
wire n_33306;
wire n_17574;
wire n_24079;
wire newNet_3334;
wire n_33889;
wire n_26212;
wire n_23880;
wire delay_sub_ln21_0_unr17_stage7_stallmux_q_9_;
wire n_23015;
wire n_11037;
wire n_12656;
wire n_44218;
wire newNet_1636;
wire n_7802;
wire n_31012;
wire n_41518;
wire n_38759;
wire n_29951;
wire n_16117;
wire n_9939;
wire n_16336;
wire FE_OCP_RBN2306_n_24288;
wire newNet_239;
wire n_17910;
wire n_7474;
wire n_19677;
wire n_211;
wire n_9492;
wire n_32885;
wire n_16957;
wire n_20838;
wire n_2248;
wire n_16119;
wire newNet_3624;
wire newNet_2773;
wire n_9394;
wire n_10260;
wire n_26263;
wire n_3690;
wire n_18681;
wire n_30227;
wire n_39733;
wire n_29401;
wire newNet_3336;
wire n_8137;
wire n_43841;
wire n_6229;
wire n_33325;
wire n_38301;
wire n_28565;
wire n_7676;
wire newNet_755;
wire n_42041;
wire n_4834;
wire n_44334;
wire n_1929;
wire n_42620;
wire n_13161;
wire n_10254;
wire n_5288;
wire delay_sub_ln21_0_unr2_stage2_stallmux_q_25_;
wire n_21196;
wire n_26574;
wire n_15804;
wire n_2527;
wire n_44570;
wire newNet_2083;
wire delay_xor_ln21_unr3_stage2_stallmux_q_12_;
wire n_17400;
wire FE_OCP_RBN3831_n_19204;
wire n_10441;
wire n_36722;
wire newNet_254;
wire n_36584;
wire n_44112;
wire n_9025;
wire n_18360;
wire n_3318;
wire n_37928;
wire n_20229;
wire n_20136;
wire n_27970;
wire n_4345;
wire FE_RN_1352_0;
wire n_37385;
wire n_41205;
wire n_7197;
wire n_26465;
wire n_40023;
wire n_30609;
wire n_22562;
wire n_41583;
wire n_38283;
wire n_6265;
wire n_36446;
wire n_41540;
wire n_25334;
wire n_44637;
wire delay_xor_ln23_unr3_stage2_stallmux_q;
wire n_21477;
wire n_7374;
wire FE_OCP_RBN3381_n_1732;
wire n_36229;
wire FE_OCP_RBN2450_n_14114;
wire n_42508;
wire newNet_2789;
wire n_2363;
wire n_27029;
wire n_25938;
wire n_6322;
wire n_12737;
wire FE_RN_1227_0;
wire n_40632;
wire n_38311;
wire n_31088;
wire n_24489;
wire n_39443;
wire n_23051;
wire n_7208;
wire n_9111;
wire n_43247;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_3_;
wire n_21409;
wire newNet_3579;
wire newNet_2976;
wire n_2910;
wire n_15403;
wire n_33797;
wire n_11570;
wire n_12813;
wire n_38943;
wire n_4272;
wire n_3565;
wire n_33093;
wire n_30486;
wire n_4668;
wire n_7510;
wire n_36367;
wire newNet_2337;
wire FE_RN_838_0;
wire n_20723;
wire n_39658;
wire n_27920;
wire n_30413;
wire FE_RN_833_0;
wire n_38449;
wire n_21684;
wire n_3770;
wire n_1286;
wire FE_RN_1529_0;
wire n_21931;
wire n_13118;
wire n_44364;
wire n_10196;
wire n_10057;
wire n_39998;
wire n_17838;
wire n_34703;
wire n_24510;
wire n_4182;
wire n_34991;
wire n_40935;
wire FE_RN_1357_0;
wire n_19940;
wire n_33680;
wire n_38859;
wire n_26793;
wire n_41291;
wire n_29352;
wire FE_RN_136_0;
wire n_15033;
wire n_18125;
wire n_4173;
wire delay_sub_ln21_0_unr27_stage10_stallmux_q_8_;
wire n_38928;
wire n_17860;
wire n_14137;
wire n_29334;
wire n_40887;
wire n_663;
wire n_42519;
wire FE_OCP_RBN2804_n_30534;
wire n_20583;
wire n_5996;
wire n_36175;
wire n_14941;
wire newNet_1672;
wire n_17881;
wire newNet_569;
wire n_7621;
wire FE_OCP_RBN1926_cordic_combinational_sub_ln23_0_unr12_z_0__;
wire n_2351;
wire newNet_1421;
wire FE_OCP_RBN2162_n_12312;
wire n_42038;
wire n_33577;
wire n_29290;
wire n_17468;
wire n_4564;
wire n_23387;
wire n_8387;
wire n_25438;
wire n_42885;
wire FE_OCP_RBN2418_n_19601;
wire n_18408;
wire n_24945;
wire FE_OCP_RBN2936_n_10626;
wire n_7954;
wire delay_sub_ln23_0_unr24_stage8_stallmux_q_9_;
wire n_10394;
wire n_43182;
wire n_43355;
wire n_1127;
wire n_27863;
wire newNet_3328;
wire n_42378;
wire n_15313;
wire n_27442;
wire n_11473;
wire n_6672;
wire n_41618;
wire n_36481;
wire n_33511;
wire n_41480;
wire n_35418;
wire n_42466;
wire n_33765;
wire n_28089;
wire newNet_1182;
wire n_5170;
wire FE_OCPN3779_n_36126;
wire FE_OCP_RBN1700_n_19353;
wire n_18534;
wire n_25248;
wire n_45217;
wire n_25566;
wire newNet_3553;
wire n_29197;
wire n_7329;
wire n_43859;
wire n_25363;
wire newNet_3030;
wire n_33117;
wire newNet_265;
wire delay_sub_ln23_0_unr5_stage3_stallmux_q_10_;
wire n_23186;
wire newNet_1499;
wire FE_OCP_RBN3827_n_18951;
wire FE_OCPN973_n_15900;
wire n_29840;
wire n_553;
wire FE_OCP_RBN3270_n_45224;
wire n_45745;
wire n_5001;
wire n_13767;
wire n_13934;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_21_;
wire n_28145;
wire newNet_981;
wire n_2146;
wire n_11289;
wire n_15344;
wire FE_OFN745_n_23604;
wire n_22619;
wire n_39157;
wire n_27839;
wire n_20556;
wire n_33107;
wire n_27186;
wire n_24596;
wire n_29378;
wire n_35583;
wire n_46980;
wire n_26022;
wire n_19544;
wire n_19393;
wire n_10632;
wire n_16920;
wire delay_sub_ln23_0_unr28_stage9_stallmux_q_16_;
wire newNet_2672;
wire n_42916;
wire n_35267;
wire n_34865;
wire n_27320;
wire FE_OCP_RBN3673_n_30820;
wire n_15953;
wire n_9400;
wire FE_OCP_RBN3395_n_28651;
wire FE_RN_923_0;
wire FE_OCP_RBN1348_n_19270;
wire n_790;
wire n_3633;
wire n_17603;
wire n_36678;
wire n_36662;
wire n_40667;
wire n_42971;
wire n_29645;
wire n_5489;
wire n_21356;
wire n_7736;
wire n_1796;
wire n_15815;
wire n_25424;
wire n_30634;
wire n_22242;
wire n_37571;
wire newNet_3340;
wire n_11048;
wire n_10795;
wire n_10601;
wire n_7020;
wire n_39594;
wire n_122;
wire newNet_560;
wire FE_OCP_RBN1920_n_22476;
wire FE_RN_31_0;
wire n_5714;
wire n_41767;
wire n_19319;
wire n_34604;
wire FE_RN_1338_0;
wire n_14198;
wire n_24057;
wire n_8879;
wire n_16526;
wire n_37345;
wire n_33077;
wire n_42652;
wire n_37746;
wire n_2763;
wire n_39465;
wire n_41246;
wire FE_OFN782_delay_sub_ln23_0_unr15_stage6_stallmux_q;
wire newNet_3104;
wire n_23525;
wire n_23732;
wire n_32731;
wire n_25622;
wire n_19475;
wire n_37044;
wire n_4644;
wire FE_RN_1701_0;
wire n_12898;
wire n_23572;
wire n_1186;
wire n_10289;
wire n_5675;
wire cos_out_2;
wire n_38842;
wire n_31690;
wire n_22460;
wire n_6862;
wire n_25738;
wire n_39546;
wire n_34735;
wire n_37095;
wire n_19370;
wire FE_RN_388_0;
wire n_5209;
wire n_39804;
wire n_2595;
wire n_28322;
wire n_19899;
wire n_27828;
wire n_17556;
wire n_13413;
wire n_11073;
wire n_41835;
wire newNet_2321;
wire newNet_136;
wire newNet_2188;
wire n_18964;
wire n_11805;
wire n_5776;
wire n_18517;
wire FE_OCP_RBN2196_n_2103;
wire n_36243;
wire newNet_2911;
wire n_3468;
wire newNet_125;
wire n_25415;
wire n_112;
wire FE_OCP_RBN2925_n_10525;
wire n_1365;
wire n_8851;
wire n_18384;
wire n_21547;
wire n_9813;
wire n_35536;
wire n_17241;
wire n_27537;
wire n_31757;
wire n_1315;
wire FE_RN_105_0;
wire n_14524;
wire newNet_2472;
wire n_35675;
wire n_28106;
wire n_19441;
wire n_3479;
wire n_12564;
wire n_35126;
wire n_21753;
wire n_15692;
wire n_3990;
wire n_3293;
wire n_6797;
wire n_18655;
wire n_37510;
wire n_29579;
wire n_7396;
wire n_5446;
wire n_43156;
wire n_33032;
wire n_28440;
wire FE_RN_1400_0;
wire n_18794;
wire n_35989;
wire n_12038;
wire n_26742;
wire n_21557;
wire n_42719;
wire n_2464;
wire n_32770;
wire FE_OCP_RBN1682_n_33491;
wire FE_OCP_RBN2197_n_12830;
wire n_26652;
wire n_27128;
wire n_25042;
wire n_35372;
wire n_17273;
wire n_18056;
wire n_14734;
wire n_30305;
wire n_27018;
wire n_37517;
wire n_32594;
wire n_21300;
wire n_17425;
wire n_1051;
wire n_16873;
wire n_832;
wire FE_RN_363_0;
wire n_1033;
wire n_19784;
wire n_39401;
wire FE_OCP_RBN2368_n_38545;
wire n_13669;
wire FE_OCP_RBN2832_n_26081;
wire n_11822;
wire n_30470;
wire n_67;
wire n_41261;
wire n_13339;
wire n_8920;
wire n_14283;
wire n_23707;
wire n_21138;
wire n_39113;
wire n_10120;
wire n_33786;
wire FE_OCPN3781_n_16440;
wire n_7277;
wire n_9225;
wire newNet_3263;
wire FE_OCP_RBN2845_n_10326;
wire n_18173;
wire n_6370;
wire n_14278;
wire n_38791;
wire FE_RN_807_0;
wire n_16513;
wire n_7082;
wire n_26371;
wire n_33379;
wire n_4818;
wire n_4140;
wire n_42891;
wire newNet_3217;
wire n_37655;
wire n_43203;
wire n_7358;
wire n_1850;
wire n_8955;
wire n_37837;
wire n_6237;
wire n_30942;
wire n_23986;
wire n_5484;
wire n_8441;
wire n_21663;
wire newNet_707;
wire n_12610;
wire n_34751;
wire n_41639;
wire n_32394;
wire n_17342;
wire n_15517;
wire newNet_2849;
wire n_1328;
wire n_25154;
wire n_14065;
wire n_16144;
wire n_42384;
wire n_25655;
wire n_40274;
wire newNet_1601;
wire n_29076;
wire n_37987;
wire n_4487;
wire n_33691;
wire n_3654;
wire n_5300;
wire FE_OCP_RBN2362_n_13785;
wire n_13541;
wire n_4937;
wire n_44445;
wire n_43889;
wire n_11215;
wire newNet_2106;
wire n_46197;
wire n_35406;
wire n_36494;
wire n_34242;
wire n_11776;
wire n_46986;
wire n_15741;
wire n_12847;
wire n_2015;
wire n_31257;
wire n_6479;
wire n_22746;
wire n_8216;
wire n_40304;
wire sin_out_17;
wire n_15175;
wire FE_OCP_RBN2541_n_8800;
wire n_11102;
wire n_10553;
wire n_18500;
wire n_10007;
wire n_32972;
wire n_40329;
wire newNet_1703;
wire FE_OCP_RBN2259_n_18899;
wire n_23503;
wire n_10771;
wire n_40960;
wire n_26110;
wire n_24170;
wire n_21361;
wire n_17829;
wire n_2193;
wire n_645;
wire n_27150;
wire n_18571;
wire n_4727;
wire n_19300;
wire n_797;
wire n_8067;
wire n_38001;
wire n_28904;
wire n_37556;
wire n_10699;
wire n_22937;
wire newNet_3094;
wire newNet_1103;
wire newNet_1974;
wire n_22782;
wire n_24468;
wire n_622;
wire FE_OCP_RBN2142_FE_OCPN861_n_45450;
wire n_5312;
wire n_41668;
wire n_24967;
wire n_34386;
wire n_46173;
wire n_20491;
wire n_14751;
wire n_45196;
wire n_23501;
wire n_19592;
wire n_41988;
wire FE_RN_1262_0;
wire n_19914;
wire n_34141;
wire n_15026;
wire newNet_3564;
wire newNet_1358;
wire n_16472;
wire n_32279;
wire n_1918;
wire n_11800;
wire n_1868;
wire n_2756;
wire n_16752;
wire n_36434;
wire n_2988;
wire FE_OCPN1775_n_18263;
wire n_25509;
wire n_38950;
wire n_32006;
wire n_33616;
wire n_33044;
wire n_32410;
wire n_2600;
wire n_30299;
wire FE_OCP_RBN1057_n_18267;
wire FE_OCP_RBN1701_n_19353;
wire n_24294;
wire newNet_2870;
wire n_35465;
wire n_32665;
wire n_22675;
wire n_13405;
wire n_29055;
wire n_21265;
wire newNet_652;
wire n_12642;
wire n_42502;
wire FE_OCP_RBN3336_n_44610;
wire FE_RN_885_0;
wire n_15099;
wire FE_RN_1656_0;
wire n_36636;
wire n_8283;
wire FE_RN_533_0;
wire FE_OCP_RBN2534_n_47018;
wire FE_OCP_RBN2833_n_26081;
wire n_26139;
wire n_29028;
wire n_1804;
wire n_19998;
wire n_23058;
wire FE_OCP_RBN3359_delay_sub_ln23_unr13_stage5_stallmux_q_1_;
wire delay_xor_ln21_unr12_stage5_stallmux_q_13_;
wire n_38609;
wire newNet_50;
wire n_1812;
wire n_9207;
wire FE_OCPN1533_n_29842;
wire n_39192;
wire n_6962;
wire n_34507;
wire n_4781;
wire n_17897;
wire n_25067;
wire n_10761;
wire n_17624;
wire n_15745;
wire n_919;
wire n_12411;
wire n_37240;
wire n_9097;
wire n_2888;
wire n_7829;
wire n_38407;
wire n_32391;
wire n_16291;
wire n_37945;
wire n_23758;
wire newNet_1905;
wire n_32225;
wire delay_sub_ln21_0_unr14_stage6_stallmux_q_29_;
wire n_35392;
wire n_28162;
wire n_31315;
wire n_1739;
wire n_35814;
wire n_29990;
wire n_11643;
wire FE_OCP_RBN3471_n_7886;
wire n_39303;
wire n_7645;
wire n_20034;
wire n_3156;
wire n_3767;
wire n_40295;
wire newNet_216;
wire newNet_2604;
wire n_25800;
wire n_21640;
wire n_30446;
wire n_16793;
wire n_12795;
wire n_17728;
wire n_21119;
wire n_35356;
wire n_27354;
wire n_7469;
wire newNet_2132;
wire n_15370;
wire n_7403;
wire n_39810;
wire newNet_2411;
wire n_1992;
wire n_21202;
wire n_11271;
wire n_1421;
wire n_16565;
wire n_5657;
wire n_17888;
wire n_1835;
wire n_27453;
wire n_3839;
wire n_32370;
wire n_31145;
wire newNet_2764;
wire n_11409;
wire n_40217;
wire newNet_720;
wire newNet_2495;
wire FE_OCP_RBN3000_n_42959;
wire FE_OFN775_n_46137;
wire n_18778;
wire n_4681;
wire n_6725;
wire n_17257;
wire n_12705;
wire n_18021;
wire n_34785;
wire n_5298;
wire n_22764;
wire n_26320;
wire n_36744;
wire n_20894;
wire n_20212;
wire n_41524;
wire FE_OCP_RBN3031_n_39942;
wire n_26830;
wire FE_OCPN875_n_44672;
wire n_40532;
wire FE_OCP_RBN3650_n_35169;
wire n_35169;
wire n_41071;
wire n_41414;
wire n_36193;
wire n_7015;
wire n_40474;
wire n_4148;
wire n_46188;
wire n_23010;
wire n_43795;
wire n_31348;
wire n_17098;
wire n_41046;
wire n_4163;
wire n_42014;
wire n_26090;
wire n_30858;
wire n_7690;
wire n_37604;
wire n_40434;
wire n_18984;
wire n_7577;
wire n_32342;
wire n_39814;
wire newNet_2620;
wire FE_OCP_RBN1727_FE_RN_1583_0;
wire n_43636;
wire n_24146;
wire delay_sub_ln23_0_unr12_stage5_stallmux_q_14_;
wire n_22996;
wire n_12481;
wire n_7925;
wire n_37898;
wire n_33719;
wire FE_OCPN1010_n_7802;
wire n_32448;
wire n_29634;
wire n_34957;
wire newNet_1834;
wire n_23636;
wire n_41706;
wire n_15437;
wire n_39135;
wire n_31794;
wire n_13369;
wire n_12981;
wire n_36599;
wire n_29245;
wire n_1599;
wire n_18594;
wire n_38379;
wire n_9040;
wire n_12615;
wire FE_OCPUNCON1806_n_19801;
wire n_1129;
wire FE_OCP_RBN2287_n_2268;
wire n_29899;
wire n_1889;
wire FE_OCP_RBN3310_n_44722;
wire FE_OCP_RBN2591_n_14460;
wire FE_RN_64_0;
wire n_26150;
wire FE_OCP_RBN2543_n_9082;
wire n_31601;
wire FE_RN_216_0;
wire n_26310;
wire n_3522;
wire n_31832;
wire n_8177;
wire n_31126;
wire n_8344;
wire n_28791;
wire n_24610;
wire n_43821;
wire newNet_2390;
wire n_31095;
wire n_27065;
wire FE_OCP_RBN2577_n_47017;
wire n_756;
wire n_44425;
wire n_6317;
wire n_43565;
wire n_28755;
wire n_38397;
wire n_33999;
wire n_39704;
wire n_30272;
wire FE_OCP_RBN3030_n_39942;
wire n_26198;
wire n_16199;
wire n_7537;
wire n_24683;
wire n_7540;
wire n_33855;
wire FE_OCPN1431_n_29504;
wire n_38125;
wire n_9380;
wire newNet_1405;
wire newNet_992;
wire n_43046;
wire FE_OFN760_n_45813;
wire n_3604;
wire n_804;
wire newNet_1116;
wire n_12047;
wire n_35394;
wire n_18458;
wire n_29770;
wire n_13709;
wire n_15532;
wire n_4255;
wire n_27243;
wire n_15349;
wire n_12362;
wire n_33152;
wire n_19274;
wire FE_RN_448_0;
wire n_35227;
wire n_40773;
wire n_11176;
wire FE_OCP_RBN1201_n_25763;
wire newNet_1173;
wire n_37268;
wire n_40320;
wire n_11726;
wire FE_OCPN897_n_44776;
wire n_24186;
wire n_16815;
wire n_24445;
wire n_21807;
wire n_25816;
wire newNet_355;
wire n_24455;
wire beta_14;
wire n_27502;
wire n_10494;
wire n_26027;
wire n_802;
wire n_17319;
wire n_29068;
wire n_12537;
wire FE_RN_469_0;
wire n_3668;
wire delay_add_ln22_unr2_stage2_stallmux_q_23_;
wire n_38363;
wire n_33357;
wire n_27948;
wire n_24755;
wire n_23763;
wire newNet_2264;
wire n_10052;
wire n_1269;
wire n_39174;
wire n_35444;
wire n_17696;
wire n_36918;
wire n_33958;
wire n_30234;
wire FE_OCPN3785_FE_OCP_RBN2831_n_10198;
wire newNet_773;
wire n_11337;
wire n_43069;
wire n_4890;
wire n_13686;
wire n_43418;
wire n_2533;
wire FE_OCP_RBN2216_FE_OCPN950_n_28595;
wire n_35374;
wire n_25528;
wire n_36370;
wire n_28610;
wire n_35063;
wire n_19211;
wire n_1551;
wire n_13657;
wire n_8460;
wire n_3034;
wire n_25846;
wire n_20343;
wire FE_OCP_RBN2737_n_15300;
wire n_15003;
wire newNet_497;
wire n_45840;
wire n_39254;
wire n_29795;
wire n_19921;
wire newNet_3137;
wire n_30094;
wire FE_OCP_DRV_N1581_n_35500;
wire delay_sub_ln23_0_unr8_stage4_stallmux_q_8_;
wire n_36618;
wire n_24647;
wire FE_OFN840_n_3500;
wire n_12068;
wire n_43314;
wire n_33291;
wire n_3081;
wire n_11265;
wire n_39292;
wire newNet_841;
wire delay_xor_ln22_unr15_stage6_stallmux_q_0_;
wire n_5260;
wire n_14182;
wire FE_OCP_RBN3096_n_43489;
wire newNet_3016;
wire n_33088;
wire n_11514;
wire n_36071;
wire n_4401;
wire FE_RN_1463_0;
wire newNet_1650;
wire n_31774;
wire n_889;
wire n_34176;
wire n_31221;
wire n_16104;
wire n_11609;
wire FE_OCP_RBN2307_n_24288;
wire FE_OFN824_n_3500;
wire n_14692;
wire n_14334;
wire delay_sub_ln23_0_unr2_stage2_stallmux_q_14_;
wire n_31668;
wire n_11693;
wire n_1600;
wire FE_OCP_RBN3398_n_37624;
wire n_10434;
wire n_2661;
wire n_34234;
wire FE_OCP_RBN2467_n_8767;
wire n_34078;
wire n_5069;
wire n_4517;
wire n_32187;
wire n_4434;
wire n_42913;
wire n_10912;
wire n_29151;
wire newNet_692;
wire n_32480;
wire FE_RN_70_0;
wire n_470;
wire FE_OCP_RBN3386_n_33108;
wire n_18936;
wire n_32169;
wire n_15874;
wire FE_RN_125_0;
wire n_21373;
wire n_20054;
wire n_33336;
wire n_22807;
wire n_14332;
wire newNet_970;
wire n_32523;
wire n_11520;
wire n_12807;
wire n_10198;
wire n_17655;
wire n_30420;
wire n_29045;
wire newNet_2040;
wire n_18200;
wire n_2101;
wire n_16278;
wire n_433;
wire n_24743;
wire n_7251;
wire FE_RN_1787_0;
wire n_4929;
wire n_19345;
wire newNet_2290;
wire n_178;
wire n_19762;
wire n_23365;
wire n_6977;
wire n_10301;
wire n_37457;
wire n_28735;
wire newNet_1232;
wire n_22237;
wire FE_RN_1064_0;
wire newNet_3246;
wire n_29418;
wire n_14555;
wire n_23156;
wire n_12721;
wire n_41305;
wire newNet_71;
wire n_36305;
wire n_17848;
wire n_24784;
wire FE_RN_954_0;
wire newNet_676;
wire n_2862;
wire n_6636;
wire n_41874;
wire n_14229;
wire n_13976;
wire n_3261;
wire n_27347;
wire delay_sub_ln21_0_unr11_stage5_stallmux_q_20_;
wire n_39076;
wire n_32046;
wire n_15189;
wire delay_xor_ln21_unr12_stage5_stallmux_q_11_;
wire n_27549;
wire n_40830;
wire n_25954;
wire n_43709;
wire delay_xor_ln22_unr9_stage4_stallmux_q_13_;
wire n_26293;
wire n_7896;
wire FE_OCP_RBN3596_FE_OCPN1243_n_44460;
wire n_38633;
wire n_43652;
wire n_32635;
wire n_20622;
wire n_32836;
wire FE_RN_618_0;
wire n_12022;
wire n_36146;
wire n_22643;
wire newNet_547;
wire n_24274;
wire n_9733;
wire n_14420;
wire n_14417;
wire n_59;
wire n_22048;
wire newNet_2062;
wire newNet_2894;
wire n_10995;
wire n_12181;
wire n_3229;
wire delay_add_ln22_unr17_stage7_stallmux_q_13_;
wire n_9954;
wire n_13857;
wire delay_xor_ln21_unr6_stage3_stallmux_q_1_;
wire n_43026;
wire n_42131;
wire n_3612;
wire n_43332;
wire newNet_2159;
wire n_42066;
wire n_2292;
wire n_34571;
wire n_10712;
wire n_42198;
wire n_10617;
wire n_8414;
wire FE_RN_1818_0;
wire n_19694;
wire n_3794;
wire n_28681;
wire n_25895;
wire n_26472;
wire n_5897;
wire n_3681;
wire FE_OFN814_n_18287;
wire n_8070;
wire newNet_1620;
wire n_46167;
wire n_39282;
wire n_32305;
wire n_15993;
wire n_5839;
wire n_26912;
wire n_32801;
wire n_30349;
wire n_11874;
wire newNet_2307;
wire FE_OCPN1859_n_35415;
wire n_23177;
wire n_40738;
wire n_37969;
wire n_4357;
wire n_21851;
wire n_35100;
wire n_27881;
wire n_27468;
wire n_13967;
wire n_6292;
wire n_20264;
wire n_10915;
wire n_10212;
wire n_40563;
wire n_28035;
wire n_4030;
wire n_44800;
wire n_38772;
wire n_17700;
wire n_9780;
wire newNet_60;
wire n_11735;
wire newNet_826;
wire n_30892;
wire n_24474;
wire n_106;
wire n_2838;
wire n_32136;
wire newNet_2747;
wire newNet_1660;
wire n_22816;
wire delay_add_ln22_unr8_stage4_stallmux_q_7_;
wire n_21882;
wire n_8025;
wire n_40718;
wire n_29024;
wire n_14214;
wire newNet_2609;
wire n_41506;
wire n_31401;
wire n_9422;
wire n_33966;
wire n_33337;
wire newNet_860;
wire n_40796;
wire FE_OCP_RBN1711_n_21087;
wire n_34016;
wire FE_RN_619_0;
wire n_38138;
wire FE_RN_1229_0;
wire n_1374;
wire n_47183;
wire n_18071;
wire n_17332;
wire n_12666;
wire n_42848;
wire n_21587;
wire n_2336;
wire n_30500;
wire n_32890;
wire n_40917;
wire newNet_2532;
wire n_8748;
wire n_1029;
wire n_4613;
wire n_37947;
wire n_28231;
wire delay_sub_ln23_0_unr20_stage7_stallmux_q_26_;
wire n_18333;
wire n_35155;
wire n_23036;
wire n_42734;
wire n_10991;
wire n_17396;
wire n_12552;
wire n_7437;
wire n_25598;
wire n_16432;
wire n_36784;
wire FE_RN_1018_0;
wire n_14019;
wire n_9445;

// Start cells
in01f80 g777999 ( .a(n_3086), .o(n_3165) );
na03f80 g742748 ( .a(n_37230), .b(n_37289), .c(n_36973), .o(n_37348) );
no02f80 g768800 ( .a(n_11958), .b(n_11924), .o(n_11925) );
na02f80 g747181 ( .a(n_32702), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(n_32701) );
na02f80 g756560 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_23_), .o(n_23757) );
no03m80 g774079 ( .a(n_6716), .b(FE_OCP_RBN3373_n_6745), .c(n_6715), .o(n_6775) );
ao12f80 g746110 ( .a(n_33731), .b(n_33777), .c(n_33830), .o(n_33877) );
no02f80 g776594 ( .a(n_4352), .b(n_4148), .o(n_4413) );
na02f80 g777331 ( .a(FE_OCP_RBN2731_n_4219), .b(FE_OFN820_n_4333), .o(n_4426) );
oa12f80 FE_RC_2608_0 ( .a(FE_RN_1083_0), .b(FE_RN_1084_0), .c(n_17954), .o(n_18056) );
na02f80 g782634 ( .a(n_40655), .b(n_40654), .o(n_44027) );
no02f80 g748388 ( .a(FE_OCPN1052_n_31674), .b(n_31502), .o(n_31791) );
in01f80 newInst_410 ( .a(newNet_409), .o(newNet_410) );
in01f80 g756638 ( .a(n_23651), .o(n_23652) );
in01f80 g754886 ( .a(n_25562), .o(n_25563) );
in01f80 g768902 ( .a(n_11777), .o(n_11823) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_4_ ( .ck(newNet_2351), .d(n_35474), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_) );
na02f80 g774726 ( .a(n_6329), .b(n_6348), .o(n_6393) );
ao12f80 g751080 ( .a(n_28507), .b(n_28852), .c(n_28532), .o(n_28894) );
in01f80 g740911 ( .a(n_39808), .o(n_39427) );
in01f80 newInst_3491 ( .a(newNet_3490), .o(newNet_3491) );
in01f80 g759966 ( .a(n_47175), .o(n_22036) );
in01f80 g751951 ( .a(n_28924), .o(n_28925) );
no02f80 g741334 ( .a(FE_OCP_RBN2553_n_44921), .b(n_38574), .o(n_38974) );
na02f80 g771260 ( .a(n_9353), .b(n_9318), .o(n_9495) );
no02f80 FE_RC_2319_0 ( .a(FE_RN_882_0), .b(n_36513), .o(n_36558) );
in01f80 g753147 ( .a(n_27457), .o(n_27458) );
no02f80 g740023 ( .a(n_40113), .b(n_40070), .o(n_40147) );
in01f80 g769764 ( .a(n_11169), .o(n_11170) );
na02f80 g762435 ( .a(n_18021), .b(n_17919), .o(n_18089) );
ao22s80 FE_RC_408_0 ( .a(FE_OCP_RBN3506_n_13860), .b(n_14286), .c(FE_OCP_RBN3507_n_13860), .d(n_14186), .o(n_14372) );
no02f80 g775134 ( .a(n_5827), .b(n_5839), .o(n_5921) );
no02f80 g762691 ( .a(FE_OCP_RBN2145_FE_OCPN861_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .o(n_17929) );
na02f80 g761079 ( .a(n_19168), .b(n_19056), .o(n_19273) );
no02f80 g753580 ( .a(n_26669), .b(n_26579), .o(n_26729) );
no02f80 g745651 ( .a(n_34166), .b(n_34135), .o(n_34208) );
no02f80 g777381 ( .a(n_3475), .b(n_3248), .o(n_3496) );
no02f80 g743131 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n_37038) );
no02f80 g756035 ( .a(n_24906), .b(n_23836), .o(n_24929) );
in01f80 g770719 ( .a(n_10305), .o(n_10306) );
ao12f80 g762953 ( .a(n_17963), .b(n_17962), .c(n_17961), .o(n_18416) );
ao22s80 FE_RC_3387_0 ( .a(FE_OCP_RBN1163_n_13726), .b(n_13840), .c(FE_OCP_RBN1164_n_13726), .d(n_13814), .o(n_14004) );
na02f80 g750513 ( .a(n_29559), .b(n_29558), .o(n_29560) );
in01f80 newInst_1465 ( .a(newNet_1464), .o(newNet_1465) );
in01f80 g748677 ( .a(n_32781), .o(n_32628) );
na02f80 g740617 ( .a(FE_OCP_RBN2872_n_39542), .b(n_45840), .o(n_39578) );
in01f80 FE_RC_2684_0 ( .a(FE_RN_1123_0), .o(n_8651) );
na02f80 g771747 ( .a(n_8879), .b(n_8189), .o(n_8971) );
in01f80 g761026 ( .a(n_19348), .o(n_19349) );
in01f80 g768945 ( .a(n_11787), .o(n_12088) );
in01f80 g750497 ( .a(n_29545), .o(n_29562) );
in01f80 FE_OCP_RBC2135_n_11780 ( .a(n_11780), .o(FE_OCP_RBN2135_n_11780) );
no02f80 g770335 ( .a(n_10707), .b(FE_OCP_RBN2586_n_9009), .o(n_10748) );
no02f80 g775583 ( .a(n_5284), .b(n_4606), .o(n_5293) );
in01f80 g771668 ( .a(n_9203), .o(n_9264) );
na02f80 g761497 ( .a(n_19787), .b(n_19928), .o(n_20220) );
in01f80 newInst_2576 ( .a(newNet_624), .o(newNet_2576) );
in01f80 g760944 ( .a(n_19497), .o(n_20124) );
na02f80 g737906 ( .a(FE_OCPN936_n_42192), .b(n_42191), .o(n_42403) );
in01f80 g737748 ( .a(n_43016), .o(n_42249) );
in01f80 g746695 ( .a(n_34359), .o(n_34300) );
oa22f80 g777227 ( .a(n_3705), .b(n_47341), .c(n_3604), .d(n_3240), .o(n_3751) );
in01f80 g761130 ( .a(n_19203), .o(n_19238) );
na02f80 g774828 ( .a(n_6228), .b(FE_OCP_RBN2975_n_5531), .o(n_6386) );
no02f80 g765619 ( .a(n_15105), .b(n_14192), .o(n_15099) );
in01f80 newInst_3310 ( .a(newNet_3309), .o(newNet_3310) );
no02f80 g784770 ( .a(n_14547), .b(FE_OCP_RBN3529_n_13765), .o(n_47256) );
no02f80 g780826 ( .a(n_414), .b(n_434), .o(n_435) );
oa12f80 g756673 ( .a(n_24107), .b(n_24064), .c(n_23803), .o(n_24132) );
in01f80 FE_OCP_RBC1058_n_18267 ( .a(FE_OCP_RBN1057_n_18267), .o(FE_OCP_RBN1058_n_18267) );
in01f80 g775549 ( .a(n_5681), .o(n_5702) );
in01f80 g754420 ( .a(n_25702), .o(n_25703) );
na02f80 g778023 ( .a(n_3000), .b(n_2247), .o(n_3009) );
no02f80 g736838 ( .a(n_43017), .b(n_43016), .o(n_43029) );
in01f80 newInst_644 ( .a(newNet_99), .o(newNet_644) );
in01f80 newInst_2169 ( .a(newNet_2168), .o(newNet_2169) );
no02f80 g766097 ( .a(n_14480), .b(n_14416), .o(n_14560) );
na02f80 FE_RC_2361_0 ( .a(FE_RN_912_0), .b(n_19191), .o(FE_RN_913_0) );
na02f80 g739001 ( .a(n_41144), .b(n_41143), .o(n_41145) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_0_ ( .ck(newNet_1656), .d(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_186) );
in01f80 g753289 ( .a(n_27463), .o(n_27373) );
oa12f80 g742700 ( .a(n_37481), .b(n_37480), .c(n_37479), .o(n_37544) );
in01f80 g742431 ( .a(n_38698), .o(n_38736) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_19_ ( .ck(newNet_1858), .d(n_16926), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_) );
oa12f80 g759447 ( .a(n_21111), .b(n_21110), .c(FE_OCP_RBN1729_n_20903), .o(n_21173) );
no02f80 g746169 ( .a(n_35089), .b(n_34700), .o(n_35127) );
oa22f80 g737646 ( .a(FE_OCPN887_n_42367), .b(n_42335), .c(n_42392), .d(n_42241), .o(n_42587) );
na02f80 g766797 ( .a(n_14525), .b(n_14562), .o(n_15575) );
in01f80 g780595 ( .a(n_732), .o(n_733) );
oa12f80 g755281 ( .a(n_24859), .b(n_24877), .c(n_24923), .o(n_24977) );
na02f80 g747982 ( .a(n_33030), .b(n_32723), .o(n_33119) );
no02f80 g740661 ( .a(n_39482), .b(n_39208), .o(n_39526) );
na02f80 g762333 ( .a(n_18008), .b(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_18060) );
in01f80 g739419 ( .a(n_40917), .o(n_40918) );
no02f80 g752975 ( .a(n_27931), .b(n_27923), .o(n_28195) );
in01f80 g778574 ( .a(n_2499), .o(n_2500) );
in01f80 g753844 ( .a(n_27079), .o(n_27080) );
na02f80 g766272 ( .a(n_14437), .b(n_14399), .o(n_14497) );
na02f80 g762735 ( .a(n_17826), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .o(n_17896) );
na02f80 g738403 ( .a(n_41414), .b(n_41433), .o(n_41434) );
in01f80 newInst_2658 ( .a(newNet_2657), .o(newNet_2658) );
in01f80 newInst_2019 ( .a(newNet_2018), .o(newNet_2019) );
in01f80 g763100 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n_18368) );
in01f80 FE_OCPC1789_n_18119 ( .a(n_18119), .o(FE_OCPN1789_n_18119) );
ao22s80 g776536 ( .a(n_4302), .b(n_4146), .c(n_4303), .d(n_4145), .o(n_4485) );
no02f80 g765203 ( .a(n_15771), .b(n_15300), .o(n_15408) );
in01f80 newInst_298 ( .a(newNet_297), .o(newNet_298) );
no02f80 g744580 ( .a(n_35376), .b(n_35361), .o(n_35438) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_10_ ( .ck(newNet_1653), .d(n_27016), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_) );
ao22s80 FE_RC_822_0 ( .a(n_19372), .b(n_19818), .c(FE_OCPN969_n_19342), .d(n_19819), .o(n_19922) );
oa22f80 FE_RC_3156_0 ( .a(n_17584), .b(n_17594), .c(n_16339), .d(n_17565), .o(n_17654) );
in01f80 newInst_2395 ( .a(newNet_56), .o(newNet_2395) );
na02f80 g780294 ( .a(n_1023), .b(FE_OFN50_n_1045), .o(n_1024) );
ao12f80 g740690 ( .a(n_39421), .b(n_39497), .c(n_39487), .o(n_39524) );
no02f80 g779791 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(n_1431) );
na02f80 g781298 ( .a(beta_31), .b(beta_17), .o(n_62) );
na02f80 g763866 ( .a(n_16590), .b(n_16534), .o(n_16643) );
no02f80 g760784 ( .a(n_20137), .b(n_20135), .o(n_20138) );
in01f80 g748612 ( .a(n_31334), .o(n_31335) );
in01f80 g759695 ( .a(FE_OCPN1502_n_20723), .o(n_20717) );
ms00f80 delay_sub_ln23_0_unr20_stage8_stallmux_q_reg ( .ck(newNet_1557), .d(n_28336), .o(n_44962) );
na02f80 g764177 ( .a(n_16469), .b(n_16445), .o(n_16532) );
ao22s80 g756530 ( .a(n_23572), .b(n_22858), .c(n_23678), .d(delay_add_ln22_unr14_stage6_stallmux_q_25_), .o(n_23914) );
in01f80 FE_OCPC3174_n_38799 ( .a(FE_OCPN3173_n_38799), .o(FE_OCPN3174_n_38799) );
na02f80 g776913 ( .a(n_3854), .b(n_3778), .o(n_3950) );
in01f80 g754531 ( .a(n_26351), .o(n_26352) );
na02f80 g776350 ( .a(n_4397), .b(n_4699), .o(n_4540) );
in01f80 g769135 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .o(n_11663) );
na02f80 g739577 ( .a(n_40638), .b(n_39737), .o(n_40645) );
in01f80 g744248 ( .a(n_36184), .o(n_36185) );
oa12f80 g762900 ( .a(n_17140), .b(n_17494), .c(n_17070), .o(n_17597) );
na02f80 g760131 ( .a(n_20537), .b(FE_OCP_RBN3511_n_19599), .o(n_20748) );
in01f80 FE_OCP_RBC2521_n_8951 ( .a(n_8951), .o(FE_OCP_RBN2521_n_8951) );
in01f80 g779189 ( .a(n_1894), .o(n_1895) );
in01f80 g752950 ( .a(n_27848), .o(n_27902) );
in01f80 g742518 ( .a(n_37601), .o(n_37602) );
in01f80 g780920 ( .a(n_369), .o(n_365) );
in01f80 g777040 ( .a(FE_OCP_RBN2611_n_3718), .o(n_4886) );
ao12f80 g761360 ( .a(n_18765), .b(n_19613), .c(n_18841), .o(n_19681) );
in01f80 FE_RC_2227_0 ( .a(n_37032), .o(FE_RN_809_0) );
na02f80 g753776 ( .a(n_26469), .b(n_26468), .o(n_26495) );
no02f80 g748696 ( .a(n_32557), .b(n_32536), .o(n_32607) );
oa12f80 g738089 ( .a(n_41875), .b(n_42105), .c(n_41532), .o(n_42133) );
in01f80 g763278 ( .a(n_17231), .o(n_17232) );
in01f80 g759939 ( .a(n_21624), .o(n_21697) );
na02f80 g739028 ( .a(n_41117), .b(n_41116), .o(n_41118) );
na02f80 FE_RC_4167_0 ( .a(n_18519), .b(FE_RN_1815_0), .o(FE_RN_1816_0) );
no03m80 g768386 ( .a(n_12416), .b(n_12401), .c(n_12402), .o(n_12417) );
in01f80 g763116 ( .a(n_17452), .o(n_17446) );
oa22f80 FE_RC_987_0 ( .a(n_26050), .b(n_25971), .c(n_26004), .d(n_26049), .o(n_26267) );
na02f80 g748289 ( .a(n_31522), .b(n_31501), .o(n_31523) );
in01f80 g740334 ( .a(n_40355), .o(n_40356) );
in01f80 newInst_2072 ( .a(newNet_2071), .o(newNet_2072) );
no02f80 g756822 ( .a(n_24063), .b(n_24076), .o(n_24064) );
in01f80 g771876 ( .a(n_8863), .o(n_8819) );
in01f80 g747559 ( .a(n_32471), .o(n_32429) );
no02f80 g739989 ( .a(n_40020), .b(n_40016), .o(n_40121) );
no02f80 g758778 ( .a(n_21765), .b(n_21787), .o(n_21897) );
ao22s80 FE_RC_1441_0 ( .a(n_31842), .b(n_32150), .c(n_31843), .d(n_32145), .o(n_32239) );
in01f80 newInst_2300 ( .a(newNet_2299), .o(newNet_2300) );
no02f80 g753807 ( .a(n_26327), .b(n_26208), .o(n_26375) );
na02f80 g738829 ( .a(n_44430), .b(n_41302), .o(n_41342) );
in01f80 g758806 ( .a(n_21869), .o(n_21870) );
in01f80 g778679 ( .a(n_2449), .o(n_2388) );
no02f80 g776048 ( .a(n_47004), .b(n_5178), .o(n_5325) );
no02f80 g773508 ( .a(n_7480), .b(n_6814), .o(n_7516) );
na02f80 g747726 ( .a(n_33702), .b(n_33516), .o(n_33745) );
na02f80 FE_RC_2928_0 ( .a(FE_OCPN964_n_27287), .b(FE_RN_1275_0), .o(FE_RN_1276_0) );
na02f80 g767426 ( .a(n_13503), .b(n_13209), .o(n_13587) );
no02f80 g754221 ( .a(n_25916), .b(n_25824), .o(n_26003) );
no02f80 g757343 ( .a(n_44068), .b(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .o(n_23462) );
na02f80 g738728 ( .a(n_41382), .b(n_41438), .o(n_41502) );
in01f80 g740950 ( .a(n_40177), .o(n_39426) );
no02f80 g748402 ( .a(n_31730), .b(FE_OCP_RBN1198_n_30619), .o(n_31763) );
na02f80 g767087 ( .a(n_13578), .b(n_13518), .o(n_13613) );
no02f80 FE_RC_2831_0 ( .a(FE_RN_1216_0), .b(n_23946), .o(FE_RN_1217_0) );
ao22s80 FE_RC_780_0 ( .a(FE_OCP_RBN2333_n_38446), .b(n_38160), .c(n_38161), .d(n_38446), .o(n_38534) );
in01f80 g752135 ( .a(n_28117), .o(n_28118) );
in01f80 g745610 ( .a(n_34532), .o(n_34993) );
na02f80 g755451 ( .a(FE_OCP_RBN1162_n_24701), .b(n_24574), .o(n_24697) );
in01f80 g776885 ( .a(n_4168), .o(n_4169) );
in01f80 newInst_1798 ( .a(newNet_1797), .o(newNet_1798) );
no02f80 g770047 ( .a(n_10906), .b(FE_OCP_RBN2749_n_9629), .o(n_10993) );
in01f80 newInst_901 ( .a(newNet_900), .o(newNet_901) );
in01f80 g753136 ( .a(n_27494), .o(n_27495) );
in01f80 g742260 ( .a(n_38120), .o(n_38026) );
na02f80 g773589 ( .a(n_7372), .b(delay_add_ln22_unr5_stage3_stallmux_q_20_), .o(n_7423) );
na02f80 g744460 ( .a(n_35442), .b(n_30633), .o(n_35471) );
in01f80 FE_OCP_RBC1201_n_25763 ( .a(FE_OCP_RBN1200_n_25763), .o(FE_OCP_RBN1201_n_25763) );
no02f80 g771574 ( .a(n_8973), .b(n_9013), .o(n_9190) );
na02f80 g771764 ( .a(n_9061), .b(FE_OCP_RBN3547_n_44575), .o(n_9232) );
na03f80 FE_RC_173_0 ( .a(n_18434), .b(n_18374), .c(n_18372), .o(n_18435) );
in01f80 newInst_3075 ( .a(newNet_826), .o(newNet_3075) );
ao12f80 g772896 ( .a(n_7698), .b(n_7902), .c(n_7751), .o(n_7976) );
ao22s80 g763094 ( .a(n_17816), .b(n_17602), .c(n_17817), .d(n_17603), .o(n_18488) );
in01f80 g766175 ( .a(n_47256), .o(n_14575) );
ao12f80 g739066 ( .a(n_41011), .b(n_41065), .c(n_40730), .o(n_41103) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_5_ ( .ck(newNet_3190), .d(n_35592), .o(delay_add_ln22_unr23_stage9_stallmux_q_5_) );
na02f80 g758070 ( .a(n_22650), .b(n_22728), .o(n_22786) );
no02f80 g766929 ( .a(n_13892), .b(n_13895), .o(n_14219) );
no02f80 g759743 ( .a(n_21667), .b(n_21374), .o(n_21718) );
no02f80 g737790 ( .a(n_42199), .b(n_42207), .o(n_42235) );
na02f80 g740939 ( .a(n_39215), .b(n_39027), .o(n_39258) );
no02f80 g743317 ( .a(n_36777), .b(n_36752), .o(n_36787) );
no02f80 g778117 ( .a(n_2855), .b(n_2806), .o(n_3626) );
na02f80 g773613 ( .a(n_7345), .b(n_7344), .o(n_7382) );
na02f80 g769717 ( .a(n_11198), .b(n_11200), .o(n_11229) );
na02f80 g760238 ( .a(FE_OCPN1261_n_20242), .b(FE_OCP_RBN3836_n_19241), .o(n_20459) );
no02f80 g766825 ( .a(n_14455), .b(n_14454), .o(n_15520) );
na02f80 g744692 ( .a(n_35285), .b(n_35264), .o(n_35307) );
in01f80 g780741 ( .a(n_601), .o(n_599) );
no02f80 g777931 ( .a(n_3142), .b(FE_OCP_RBN2344_FE_OCPN870_n_2737), .o(n_3183) );
no02f80 g756921 ( .a(n_23748), .b(n_23747), .o(n_23749) );
no02f80 g754709 ( .a(n_26231), .b(n_25683), .o(n_26345) );
in01f80 g771677 ( .a(n_9389), .o(n_9390) );
in01f80 newInst_2483 ( .a(newNet_2482), .o(newNet_2483) );
no02f80 g777253 ( .a(n_3640), .b(n_3672), .o(n_3828) );
in01f80 newInst_2404 ( .a(newNet_2403), .o(newNet_2404) );
no02f80 g761683 ( .a(n_18825), .b(n_18856), .o(n_18938) );
no02f80 g774942 ( .a(n_6144), .b(n_6114), .o(n_6145) );
in01f80 g737754 ( .a(n_42355), .o(n_42356) );
in01f80 newInst_2261 ( .a(newNet_2260), .o(newNet_2261) );
in01f80 g758116 ( .a(n_22129), .o(n_22128) );
ms00f80 delay_sub_ln23_unr17_stage6_stallmux_q_reg_1_ ( .ck(newNet_1056), .d(n_22549), .o(delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
no03m80 FE_RC_1667_0 ( .a(FE_OCPN1015_n_32820), .b(FE_OCP_RBN2154_n_32772), .c(n_32818), .o(n_32851) );
oa12f80 g744021 ( .a(n_36794), .b(n_36862), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36899) );
na02f80 g752911 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .o(n_27791) );
in01f80 newInst_2955 ( .a(newNet_1722), .o(newNet_2955) );
ao12f80 g771485 ( .a(n_9225), .b(n_9595), .c(n_9323), .o(n_9654) );
in01f80 g747328 ( .a(n_32754), .o(n_32715) );
no02f80 g747317 ( .a(FE_OCP_RBN2102_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .o(n_32554) );
in01f80 g768585 ( .a(n_12267), .o(n_12333) );
no02f80 g749422 ( .a(n_30561), .b(n_30539), .o(n_30622) );
in01f80 g738888 ( .a(n_41330), .o(n_41345) );
no02f80 g767036 ( .a(FE_OCP_RBN2458_n_13765), .b(n_13134), .o(n_13903) );
no02f80 g754034 ( .a(n_26086), .b(n_24433), .o(n_26212) );
in01f80 g752210 ( .a(n_28634), .o(n_28709) );
na02f80 g760101 ( .a(n_20456), .b(FE_OCP_RBN2392_n_19434), .o(n_20533) );
in01f80 g765401 ( .a(n_15296), .o(n_15412) );
in01f80 g782657 ( .a(n_44051), .o(n_44052) );
in01f80 g779116 ( .a(n_2034), .o(n_2035) );
no02f80 g761648 ( .a(n_18756), .b(n_18265), .o(n_18758) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_5_ ( .ck(newNet_2147), .d(n_1017), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_) );
na02f80 g745753 ( .a(n_34196), .b(FE_OCP_RBN3438_n_33750), .o(n_34218) );
na02f80 g775410 ( .a(n_5614), .b(n_4556), .o(n_5634) );
in01f80 g776605 ( .a(n_4430), .o(n_4431) );
no03m80 g752178 ( .a(n_27918), .b(n_27919), .c(n_27864), .o(n_28012) );
in01f80 g755122 ( .a(n_25349), .o(n_25445) );
na02f80 g753877 ( .a(n_26298), .b(n_26216), .o(n_26329) );
in01f80 g764192 ( .a(n_16594), .o(n_16595) );
in01f80 g764180 ( .a(n_16850), .o(n_16851) );
na02f80 g777191 ( .a(n_4873), .b(n_4745), .o(n_5774) );
in01f80 FE_RC_4076_0 ( .a(FE_RN_1776_0), .o(FE_RN_1774_0) );
oa22f80 FE_RC_1472_0 ( .a(FE_OFN767_n_15670), .b(n_17648), .c(n_17753), .d(n_17587), .o(n_17677) );
na02f80 g773417 ( .a(n_7544), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .o(n_7593) );
in01f80 newInst_1960 ( .a(newNet_1959), .o(newNet_1960) );
in01f80 newInst_2327 ( .a(newNet_2072), .o(newNet_2327) );
in01f80 g743966 ( .a(n_35952), .o(n_35953) );
in01f80 newInst_573 ( .a(newNet_572), .o(newNet_573) );
no02f80 g780505 ( .a(n_704), .b(n_730), .o(n_812) );
no02f80 g765312 ( .a(n_15208), .b(n_15207), .o(n_15339) );
no02f80 g739954 ( .a(n_40398), .b(n_40131), .o(n_40399) );
in01f80 FE_OCPUNCOC1806_n_19801 ( .a(FE_OCPUNCON1805_n_19801), .o(FE_OCPUNCON1806_n_19801) );
no02f80 g751405 ( .a(n_29226), .b(n_29225), .o(n_29227) );
in01f80 FE_OCP_RBC2225_n_12729 ( .a(n_12729), .o(FE_OCP_RBN2225_n_12729) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_9_ ( .ck(newNet_767), .d(n_1306), .o(delay_xor_ln21_unr3_stage2_stallmux_q_9_) );
in01f80 g759992 ( .a(n_20379), .o(n_20414) );
no02f80 g758931 ( .a(n_21233), .b(n_45024), .o(n_21365) );
na02f80 g739454 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .o(n_40873) );
in01f80 g743443 ( .a(n_36594), .o(n_36566) );
in01f80 g762155 ( .a(FE_OCP_RBN2205_n_18242), .o(n_18355) );
no03m80 g752239 ( .a(n_27937), .b(n_27970), .c(n_27936), .o(n_28037) );
in01f80 g749067 ( .a(n_31075), .o(n_31022) );
na02f80 g750553 ( .a(n_29583), .b(n_29633), .o(n_29584) );
in01f80 g743550 ( .a(n_36579), .o(n_36604) );
na02f80 g755167 ( .a(n_25042), .b(n_24694), .o(n_25048) );
in01f80 FE_OCP_RBC2973_n_5531 ( .a(n_5531), .o(FE_OCP_RBN2973_n_5531) );
no02f80 FE_RC_2643_0 ( .a(FE_RN_1102_0), .b(FE_RN_1101_0), .o(n_3545) );
no02f80 g761199 ( .a(n_19038), .b(n_19081), .o(n_19143) );
in01f80 g753733 ( .a(n_26614), .o(n_26615) );
na02f80 g777117 ( .a(n_3547), .b(n_3457), .o(n_3634) );
na02f80 g748377 ( .a(n_31449), .b(n_30322), .o(n_31477) );
in01f80 g753677 ( .a(n_26589), .o(n_26691) );
no02f80 g747321 ( .a(FE_OCP_RBN3331_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .o(n_32706) );
in01f80 FE_OCPC1428_n_13510 ( .a(FE_OCPN1427_n_13510), .o(FE_OCPN1428_n_13510) );
in01f80 FE_OCP_RBC1164_n_13726 ( .a(FE_OCP_RBN1163_n_13726), .o(FE_OCP_RBN1164_n_13726) );
no02f80 g745936 ( .a(n_33984), .b(n_34039), .o(n_34040) );
no02f80 g739945 ( .a(n_40089), .b(n_39982), .o(n_40091) );
in01f80 g750162 ( .a(n_29816), .o(n_29780) );
in01f80 FE_OCP_RBC2283_n_33846 ( .a(n_33846), .o(FE_OCP_RBN2283_n_33846) );
in01f80 g740740 ( .a(n_39551), .o(n_39550) );
ao12f80 g738093 ( .a(n_41710), .b(n_42059), .c(n_41592), .o(n_42089) );
in01f80 g776651 ( .a(n_4382), .o(n_4383) );
in01f80 FE_OCP_RBC2663_n_20333 ( .a(FE_OCP_RBN2662_n_20333), .o(FE_OCP_RBN2663_n_20333) );
na02f80 g767906 ( .a(n_12686), .b(n_12685), .o(n_12743) );
in01f80 FE_OCP_RBC2406_n_8242 ( .a(n_8242), .o(FE_OCP_RBN2406_n_8242) );
in01f80 newInst_3192 ( .a(newNet_3191), .o(newNet_3192) );
in01f80 g766577 ( .a(n_13932), .o(n_13992) );
in01f80 g779192 ( .a(n_1908), .o(n_2606) );
in01f80 g778982 ( .a(n_2226), .o(n_2227) );
in01f80 g775495 ( .a(n_5719), .o(n_5720) );
in01f80 g743665 ( .a(n_36437), .o(n_36438) );
in01f80 FE_OCP_RBC2725_n_4219 ( .a(FE_OCP_RBN2722_n_4219), .o(FE_OCP_RBN2725_n_4219) );
na02f80 g770986 ( .a(n_9472), .b(n_9465), .o(n_9541) );
in01f80 g751584 ( .a(n_28486), .o(n_28487) );
in01f80 FE_OCP_RBC2677_n_9247 ( .a(n_9247), .o(FE_OCP_RBN2677_n_9247) );
na02f80 g748752 ( .a(n_31233), .b(n_31100), .o(n_31299) );
no02f80 g768686 ( .a(n_12137), .b(delay_add_ln22_unr8_stage4_stallmux_q_5_), .o(n_12186) );
in01f80 g757939 ( .a(n_22811), .o(n_22885) );
in01f80 g755034 ( .a(n_25431), .o(n_25148) );
in01f80 g737281 ( .a(n_42888), .o(n_42900) );
in01f80 g758657 ( .a(n_21913), .o(n_21914) );
no02f80 g770318 ( .a(n_10538), .b(n_44464), .o(n_10601) );
no02f80 g756042 ( .a(n_25032), .b(n_25028), .o(n_25053) );
no02f80 g753562 ( .a(n_26724), .b(n_26333), .o(n_26757) );
in01f80 g747788 ( .a(n_33970), .o(n_33971) );
in01f80 newInst_3381 ( .a(newNet_3380), .o(newNet_3381) );
in01f80 g767591 ( .a(n_13011), .o(n_13012) );
ao12f80 g746850 ( .a(n_33225), .b(FE_OCP_RBN2169_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n_33260) );
oa12f80 g768768 ( .a(n_11698), .b(n_11958), .c(n_11924), .o(n_11964) );
oa12f80 g740566 ( .a(n_39681), .b(n_39680), .c(n_39679), .o(n_39708) );
in01f80 g771107 ( .a(n_9742), .o(n_9798) );
no02f80 g751791 ( .a(n_28251), .b(n_28030), .o(n_28287) );
in01f80 g767418 ( .a(n_13361), .o(n_13406) );
na02f80 g772502 ( .a(n_8345), .b(n_8375), .o(n_8416) );
na02f80 g763839 ( .a(n_16607), .b(n_16585), .o(n_16628) );
na02f80 g766641 ( .a(n_14261), .b(n_14260), .o(n_14262) );
no02f80 g763187 ( .a(FE_OCP_RBN3210_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .o(n_17289) );
in01f80 g738033 ( .a(n_42150), .o(n_42149) );
in01f80 g777140 ( .a(n_3750), .o(n_3843) );
in01f80 newInst_1528 ( .a(newNet_1527), .o(newNet_1528) );
no02f80 g762611 ( .a(FE_OCP_RBN2142_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .o(n_17975) );
in01f80 g766526 ( .a(FE_OCP_RBN2450_n_14114), .o(n_14274) );
no02f80 g755625 ( .a(n_24547), .b(n_24438), .o(n_24596) );
no02f80 g750124 ( .a(FE_OCP_RBN3568_n_29857), .b(n_29160), .o(n_30108) );
in01f80 g775936 ( .a(n_4849), .o(n_4850) );
na02f80 g766126 ( .a(n_14519), .b(n_13272), .o(n_14587) );
ao22s80 FE_RC_3271_0 ( .a(n_11427), .b(n_11504), .c(FE_RN_1440_0), .d(n_11503), .o(n_11669) );
no02f80 g762130 ( .a(n_18189), .b(n_17050), .o(n_18264) );
no02f80 g741504 ( .a(n_38756), .b(n_38755), .o(n_38757) );
in01f80 newInst_2780 ( .a(newNet_2779), .o(newNet_2780) );
ao22s80 FE_RC_12_0 ( .a(n_1473), .b(n_1421), .c(n_1467), .d(n_1472), .o(n_1588) );
in01f80 FE_OCPC3778_n_36126 ( .a(n_36126), .o(FE_OCPN3778_n_36126) );
oa22f80 g765259 ( .a(n_15156), .b(FE_OCP_RBN3496_n_13818), .c(FE_OCP_RBN2681_n_15048), .d(FE_OCPN1257_n_13831), .o(n_15266) );
in01f80 g779584 ( .a(n_2026), .o(n_2027) );
na02f80 g761766 ( .a(n_18789), .b(n_18744), .o(n_18745) );
in01f80 FE_OCP_RBC3666_n_10106 ( .a(FE_OCP_RBN2793_n_10106), .o(FE_OCP_RBN3666_n_10106) );
in01f80 g747124 ( .a(n_32889), .o(n_32928) );
in01f80 g736873 ( .a(n_43536), .o(n_43537) );
no02f80 g744682 ( .a(n_35213), .b(n_35207), .o(n_35214) );
in01f80 FE_OCP_RBC2334_n_24359 ( .a(n_24359), .o(FE_OCP_RBN2334_n_24359) );
no02f80 g745213 ( .a(n_34358), .b(n_34480), .o(n_34597) );
ao12f80 g755909 ( .a(n_25056), .b(n_25160), .c(n_25001), .o(n_25572) );
no02f80 FE_RC_4216_0 ( .a(FE_OCP_RBN2505_n_13896), .b(FE_RN_1845_0), .o(FE_RN_1846_0) );
in01f80 newInst_1194 ( .a(newNet_269), .o(newNet_1194) );
ao12f80 g746777 ( .a(n_34108), .b(n_34107), .c(n_34106), .o(n_34739) );
in01f80 g761528 ( .a(n_19648), .o(n_19952) );
in01f80 g755894 ( .a(n_24393), .o(n_24394) );
no02f80 g766930 ( .a(n_13970), .b(FE_RN_994_0), .o(n_14565) );
in01f80 g775890 ( .a(n_4968), .o(n_4969) );
no02f80 g771933 ( .a(n_8747), .b(n_8742), .o(n_8743) );
no02f80 g765565 ( .a(FE_OCP_RBN2716_n_14982), .b(n_14317), .o(n_15215) );
no02f80 g772751 ( .a(n_8216), .b(n_8183), .o(n_8358) );
oa22f80 g749010 ( .a(n_32233), .b(n_31633), .c(n_32232), .d(n_31634), .o(n_32274) );
oa22f80 g779026 ( .a(n_2110), .b(n_1917), .c(n_2118), .d(n_1918), .o(n_2187) );
no02f80 g749522 ( .a(n_30496), .b(n_30141), .o(n_30509) );
in01f80 fopt782736 ( .a(n_20843), .o(n_44144) );
na02f80 g776188 ( .a(n_4929), .b(n_4951), .o(n_4930) );
ao22s80 g739152 ( .a(n_40897), .b(n_40784), .c(n_40833), .d(n_40783), .o(n_41385) );
na02f80 g776950 ( .a(n_3558), .b(n_3488), .o(n_3630) );
na02f80 FE_RC_3762_0 ( .a(FE_RN_1651_0), .b(FE_RN_1652_0), .o(FE_RN_1653_0) );
in01f80 g762651 ( .a(n_18067), .o(n_18068) );
in01f80 FE_RC_2842_0 ( .a(FE_RN_1223_0), .o(n_13747) );
in01f80 newInst_2410 ( .a(newNet_1131), .o(newNet_2410) );
in01f80 g743711 ( .a(n_36390), .o(n_36391) );
in01f80 g753339 ( .a(n_27070), .o(n_27086) );
in01f80 FE_OCPC1002_n_45660 ( .a(FE_OCPN1000_n_45660), .o(FE_OCPN1002_n_45660) );
in01f80 newInst_2594 ( .a(newNet_1187), .o(newNet_2594) );
no02f80 g761881 ( .a(n_19020), .b(n_19019), .o(n_19021) );
in01f80 FE_OCP_RBC3702_n_31064 ( .a(FE_OCP_RBN3701_n_31064), .o(FE_OCP_RBN3702_n_31064) );
in01f80 newInst_2101 ( .a(newNet_394), .o(newNet_2101) );
no02f80 g759184 ( .a(n_21305), .b(n_45073), .o(n_21462) );
na02f80 g744157 ( .a(n_35545), .b(n_35517), .o(n_35573) );
oa22f80 FE_RC_289_0 ( .a(n_45091), .b(n_20941), .c(n_45013), .d(FE_OCP_RBN1335_n_20941), .o(n_21072) );
oa12f80 g764552 ( .a(n_16507), .b(n_16506), .c(n_16505), .o(n_16550) );
na02f80 g739308 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40933) );
in01f80 newInst_550 ( .a(newNet_549), .o(newNet_550) );
na02f80 g769051 ( .a(n_11592), .b(n_45224), .o(n_11779) );
in01f80 g742819 ( .a(n_37310), .o(n_37344) );
na02f80 g769781 ( .a(n_11113), .b(n_11064), .o(n_11197) );
na02f80 g750106 ( .a(FE_OCP_RBN2573_n_29922), .b(n_30191), .o(n_30213) );
na02f80 g756628 ( .a(n_24078), .b(n_23749), .o(n_24077) );
no02f80 g766726 ( .a(n_13778), .b(n_13260), .o(n_13776) );
no02f80 g772929 ( .a(n_7864), .b(FE_OCPN1392_n_7925), .o(n_7926) );
na02f80 g758650 ( .a(n_21815), .b(n_21899), .o(n_21916) );
ao12f80 g774384 ( .a(n_6826), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n_7408) );
in01f80 newInst_3505 ( .a(newNet_3504), .o(newNet_3505) );
in01f80 g775249 ( .a(n_46427), .o(n_5961) );
in01f80 g748400 ( .a(n_31763), .o(n_31788) );
no02f80 g742191 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38209), .o(n_38229) );
oa12f80 g768706 ( .a(n_12123), .b(n_12122), .c(n_12121), .o(n_13054) );
na02f80 g748952 ( .a(n_31128), .b(FE_OCPN1452_n_27518), .o(n_31236) );
ao12f80 g739399 ( .a(n_40838), .b(FE_OCPN898_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .o(n_41137) );
in01f80 g743628 ( .a(n_36501), .o(n_36532) );
na02f80 g766592 ( .a(n_13866), .b(n_47250), .o(n_13867) );
ms00f80 delay_sub_ln23_unr21_stage7_stallmux_q_reg_1_ ( .ck(newNet_1051), .d(n_27677), .o(delay_sub_ln23_unr21_stage7_stallmux_q_1_) );
na02f80 g754861 ( .a(n_25398), .b(n_25397), .o(n_25427) );
na04m80 FE_RC_1075_0 ( .a(n_46413), .b(n_32712), .c(n_32709), .d(FE_OCPN1236_n_32791), .o(n_32714) );
na02f80 g767708 ( .a(n_13129), .b(n_13126), .o(n_13212) );
no02f80 FE_RC_3494_0 ( .a(FE_RN_1506_0), .b(FE_OCP_RBN3422_n_12879), .o(n_13011) );
in01f80 g757973 ( .a(n_22108), .o(n_22109) );
na02f80 g779350 ( .a(n_1635), .b(n_1626), .o(n_1627) );
na02f80 g767554 ( .a(n_13011), .b(n_12987), .o(n_13063) );
no02f80 FE_RC_2405_0 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_3_), .b(n_6780), .o(FE_RN_947_0) );
na02f80 g747251 ( .a(n_32784), .b(delay_add_ln22_unr20_stage8_stallmux_q_3_), .o(n_32813) );
no02f80 g773467 ( .a(n_7560), .b(n_7157), .o(n_7563) );
na02f80 g743819 ( .a(n_36335), .b(n_36334), .o(n_36336) );
ao12f80 g764163 ( .a(n_16461), .b(n_16439), .c(n_16437), .o(n_16565) );
oa12f80 g778146 ( .a(n_2180), .b(n_2801), .c(n_2141), .o(n_2884) );
in01f80 g770402 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_8_), .o(n_10611) );
in01f80 newInst_3582 ( .a(newNet_3297), .o(newNet_3582) );
na02f80 g777667 ( .a(n_3447), .b(n_3408), .o(n_3519) );
in01f80 g737471 ( .a(n_46944), .o(n_42668) );
no02f80 g749927 ( .a(n_29918), .b(n_29986), .o(n_29963) );
in01f80 g745130 ( .a(n_36179), .o(n_36180) );
in01f80 g765864 ( .a(n_15711), .o(n_15360) );
in01f80 g739593 ( .a(n_40616), .o(n_40633) );
in01f80 FE_OCP_RBC2638_n_38806 ( .a(FE_OCP_RBN2636_n_38806), .o(FE_OCP_RBN2638_n_38806) );
na02f80 g745315 ( .a(n_35799), .b(n_35884), .o(n_35852) );
oa12f80 g752642 ( .a(n_27506), .b(n_27533), .c(n_27422), .o(n_27578) );
no02f80 g771236 ( .a(n_9639), .b(n_9616), .o(n_9879) );
no02f80 g780387 ( .a(n_937), .b(n_872), .o(n_873) );
no02f80 g773864 ( .a(n_7071), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .o(n_7095) );
no02f80 g768105 ( .a(n_12662), .b(n_12079), .o(n_12670) );
in01f80 g757529 ( .a(n_23897), .o(n_23341) );
oa22f80 FE_RC_403_0 ( .a(FE_OCP_RBN3497_n_13818), .b(n_14052), .c(FE_OCP_RBN3496_n_13818), .d(n_14088), .o(n_14278) );
na02f80 FE_RC_2892_0 ( .a(n_33881), .b(FE_RN_1252_0), .o(n_34017) );
ao22s80 g756512 ( .a(n_23606), .b(n_22717), .c(n_23599), .d(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n_23759) );
in01f80 g765973 ( .a(n_14811), .o(n_14812) );
in01f80 g761510 ( .a(n_19876), .o(n_19789) );
na02f80 g740369 ( .a(n_39787), .b(n_39085), .o(n_40045) );
oa12f80 g743911 ( .a(n_46249), .b(n_36861), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36978) );
no02f80 g750147 ( .a(n_29869), .b(n_29112), .o(n_29915) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_22_ ( .ck(newNet_1402), .d(n_36680), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_) );
na02f80 g753507 ( .a(n_26805), .b(n_26826), .o(n_26957) );
no02f80 g748681 ( .a(n_31329), .b(n_31075), .o(n_31400) );
in01f80 g767161 ( .a(n_14452), .o(n_14650) );
in01f80 FE_RC_2027_0 ( .a(FE_RN_675_0), .o(n_25939) );
na02f80 FE_RC_2114_0 ( .a(FE_RN_731_0), .b(n_21084), .o(FE_RN_732_0) );
in01f80 newInst_601 ( .a(newNet_600), .o(newNet_601) );
na02f80 g759774 ( .a(n_21248), .b(n_21826), .o(n_21375) );
in01f80 g754091 ( .a(n_26178), .o(n_26122) );
in01f80 g780821 ( .a(n_491), .o(n_492) );
na02f80 g778464 ( .a(n_2344), .b(n_2343), .o(n_2345) );
na02f80 g751026 ( .a(n_28894), .b(n_28893), .o(n_28934) );
in01f80 newInst_2878 ( .a(newNet_2877), .o(newNet_2878) );
ao12f80 g774194 ( .a(n_6772), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .o(n_6979) );
in01f80 g769992 ( .a(n_11003), .o(n_11022) );
oa12f80 g757792 ( .a(n_22173), .b(n_22356), .c(n_22042), .o(n_22450) );
in01f80 newInst_438 ( .a(newNet_437), .o(newNet_438) );
in01f80 g744879 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .o(n_36785) );
in01f80 g774686 ( .a(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6806) );
no02f80 g771699 ( .a(n_8841), .b(n_7582), .o(n_8910) );
no02f80 g774310 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .o(n_7006) );
in01f80 newInst_2186 ( .a(newNet_2185), .o(newNet_2186) );
in01f80 g774256 ( .a(n_6590), .o(n_6674) );
in01f80 g768446 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_20_), .o(n_12381) );
no02f80 g742802 ( .a(n_37281), .b(n_37121), .o(n_37282) );
in01f80 g772522 ( .a(n_8535), .o(n_8488) );
no02f80 g754912 ( .a(n_25327), .b(n_25390), .o(n_25393) );
in01f80 newInst_3689 ( .a(newNet_1816), .o(newNet_3689) );
na02f80 g742381 ( .a(n_37769), .b(n_37746), .o(n_37822) );
ao12f80 g780756 ( .a(n_544), .b(n_547), .c(n_543), .o(n_701) );
in01f80 g755207 ( .a(n_25374), .o(n_25373) );
in01f80 g754264 ( .a(n_25919), .o(n_25935) );
na02f80 g748604 ( .a(n_31333), .b(n_31382), .o(n_31401) );
na02f80 g768693 ( .a(n_12181), .b(n_12273), .o(n_12331) );
in01f80 newInst_1455 ( .a(newNet_1454), .o(newNet_1455) );
in01f80 FE_OCP_RBC3437_n_33750 ( .a(n_33750), .o(FE_OCP_RBN3437_n_33750) );
ao22s80 g740707 ( .a(n_39515), .b(n_39173), .c(n_39514), .d(n_39174), .o(n_39584) );
in01f80 FE_RC_3558_0 ( .a(FE_RN_1545_0), .o(n_29684) );
in01f80 newInst_866 ( .a(newNet_86), .o(newNet_866) );
na02f80 g761923 ( .a(n_18508), .b(n_18424), .o(n_18786) );
na02f80 g779203 ( .a(n_1847), .b(n_1846), .o(n_1848) );
na02f80 g776169 ( .a(n_4554), .b(n_4219), .o(n_4716) );
in01f80 g775099 ( .a(n_6096), .o(n_6097) );
na02f80 g780903 ( .a(n_420), .b(n_443), .o(n_461) );
na02f80 g773093 ( .a(n_7712), .b(n_7957), .o(n_7720) );
na02f80 g746591 ( .a(n_34666), .b(n_34774), .o(n_34839) );
oa12f80 g773111 ( .a(n_7854), .b(n_8362), .c(n_7888), .o(n_8716) );
no02f80 g759711 ( .a(n_20545), .b(n_45008), .o(n_20591) );
na02f80 g737085 ( .a(n_43097), .b(n_42957), .o(n_43273) );
na02f80 g749585 ( .a(n_31672), .b(n_31221), .o(n_31692) );
in01f80 FE_RC_2112_0 ( .a(n_45023), .o(FE_RN_731_0) );
in01f80 FE_OCP_RBC1196_n_30926 ( .a(n_30926), .o(FE_OCP_RBN1196_n_30926) );
in01f80 g781275 ( .a(n_104), .o(n_74) );
in01f80 g749530 ( .a(n_31885), .o(n_31886) );
in01f80 g769166 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .o(n_11558) );
na02f80 g764877 ( .a(n_15687), .b(n_15686), .o(n_15793) );
na02f80 g760649 ( .a(FE_OCP_RBN3520_n_19663), .b(FE_OCPN1426_n_18099), .o(n_19729) );
oa22f80 g748856 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .c(n_32271), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_33045) );
in01f80 newInst_2814 ( .a(newNet_2813), .o(newNet_2814) );
in01f80 g773520 ( .a(n_7494), .o(n_7495) );
oa12f80 g782664 ( .a(n_8493), .b(n_8443), .c(n_8316), .o(n_44058) );
ao12f80 g755196 ( .a(n_25642), .b(n_25660), .c(n_25641), .o(n_25712) );
in01f80 FE_RC_3294_0 ( .a(n_23015), .o(FE_RN_1449_0) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_15_ ( .ck(newNet_740), .d(n_46157), .o(delay_xor_ln21_unr6_stage3_stallmux_q_15_) );
ao12f80 g745249 ( .a(n_34131), .b(n_34275), .c(n_34150), .o(n_34570) );
in01f80 g737703 ( .a(n_42332), .o(n_42333) );
in01f80 g761758 ( .a(n_18439), .o(n_18519) );
na02f80 g763420 ( .a(n_16902), .b(n_16944), .o(n_17031) );
in01f80 FE_OCP_RBC2228_n_7598 ( .a(n_7598), .o(FE_OCP_RBN2228_n_7598) );
in01f80 newInst_2510 ( .a(newNet_706), .o(newNet_2510) );
in01f80 g779469 ( .a(n_1804), .o(n_1805) );
no02f80 g744949 ( .a(n_34862), .b(n_34882), .o(n_34955) );
na02f80 g774516 ( .a(n_6524), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .o(n_6540) );
na02f80 g771823 ( .a(n_9811), .b(n_9733), .o(n_9776) );
na02f80 g771078 ( .a(n_9840), .b(n_9706), .o(n_9887) );
in01f80 g744595 ( .a(n_35377), .o(n_35437) );
in01f80 FE_OCP_RBC3309_n_44722 ( .a(FE_OCP_RBN3310_n_44722), .o(FE_OCP_RBN3309_n_44722) );
na02f80 g763353 ( .a(FE_OCP_RBN3214_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .o(n_16915) );
in01f80 g772670 ( .a(n_8283), .o(n_8305) );
no02f80 g765053 ( .a(n_15530), .b(n_13742), .o(n_15531) );
in01f80 g751347 ( .a(n_29908), .o(n_29509) );
no02f80 g747466 ( .a(n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .o(n_32568) );
in01f80 g766818 ( .a(n_14352), .o(n_14353) );
no02f80 g769053 ( .a(FE_OCP_RBN3265_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .o(n_11882) );
in01f80 g763255 ( .a(n_17287), .o(n_17275) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_19_ ( .ck(newNet_2293), .d(n_40477), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_3_ ( .ck(newNet_3487), .d(n_21302), .o(delay_add_ln22_unr14_stage6_stallmux_q_3_) );
in01f80 g778657 ( .a(n_3319), .o(n_2416) );
na02f80 g764313 ( .a(n_16398), .b(n_14805), .o(n_16399) );
in01f80 g756026 ( .a(n_25031), .o(n_25086) );
na02f80 g764700 ( .a(n_16031), .b(n_16030), .o(n_16032) );
oa22f80 g736910 ( .a(n_43230), .b(n_43494), .c(FE_OCP_RBN3067_n_43230), .d(n_43121), .o(n_43632) );
na02f80 g758883 ( .a(n_22331), .b(n_45081), .o(n_21441) );
no02f80 g752949 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .o(n_28280) );
in01f80 g748032 ( .a(n_33003), .o(n_32982) );
na02f80 g745604 ( .a(n_34369), .b(FE_OCP_RBN1681_n_33491), .o(n_34458) );
no02f80 g738296 ( .a(n_41916), .b(n_41915), .o(n_41917) );
oa22f80 g779849 ( .a(n_44652), .b(n_1022), .c(n_44623), .d(n_957), .o(n_1355) );
oa12f80 g769848 ( .a(n_10161), .b(n_11180), .c(n_10160), .o(n_11267) );
in01f80 newInst_3189 ( .a(newNet_3188), .o(newNet_3189) );
in01f80 newInst_1606 ( .a(newNet_1605), .o(newNet_1606) );
na02f80 g752199 ( .a(n_28559), .b(n_28558), .o(n_28560) );
na02f80 g754907 ( .a(FE_OCP_RBN2596_n_25181), .b(n_24486), .o(n_25973) );
in01f80 g776204 ( .a(n_4946), .o(n_4995) );
in01f80 newInst_2723 ( .a(newNet_2722), .o(newNet_2723) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_4_ ( .ck(newNet_3195), .d(n_35518), .o(delay_add_ln22_unr23_stage9_stallmux_q_4_) );
in01f80 newInst_2764 ( .a(newNet_2763), .o(newNet_2764) );
in01f80 g762909 ( .a(n_18064), .o(n_18065) );
in01f80 g762317 ( .a(n_18091), .o(n_18092) );
in01f80 g747363 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_6_), .o(n_32440) );
ao22s80 g766360 ( .a(n_14176), .b(n_13514), .c(n_14225), .d(n_13515), .o(n_14362) );
in01f80 g770780 ( .a(n_10072), .o(n_10109) );
in01f80 g737220 ( .a(n_42948), .o(n_42949) );
na02f80 g765932 ( .a(n_14798), .b(FE_OCP_RBN3528_n_13765), .o(n_14796) );
in01f80 g747751 ( .a(n_32300), .o(n_32296) );
na02f80 g741467 ( .a(n_38808), .b(n_38807), .o(n_38809) );
oa12f80 g738306 ( .a(n_41454), .b(n_41648), .c(n_41477), .o(n_41842) );
na02f80 g748074 ( .a(n_32843), .b(n_32422), .o(n_32844) );
in01f80 g778529 ( .a(n_2556), .o(n_2629) );
in01f80 g773382 ( .a(n_7574), .o(n_7575) );
in01f80 g740324 ( .a(n_40396), .o(n_40397) );
ao12f80 g775680 ( .a(n_5160), .b(n_5539), .c(n_5204), .o(n_5571) );
in01f80 g760891 ( .a(FE_OCP_RBN2392_n_19434), .o(n_20528) );
in01f80 newInst_2801 ( .a(newNet_2139), .o(newNet_2801) );
in01f80 g738839 ( .a(n_41325), .o(n_41340) );
oa12f80 g779137 ( .a(n_1942), .b(n_2606), .c(FE_OFN810_n_1941), .o(n_4117) );
na02f80 g739330 ( .a(n_40873), .b(n_40761), .o(n_40762) );
in01f80 newInst_460 ( .a(newNet_459), .o(newNet_460) );
no02f80 g772415 ( .a(n_8530), .b(n_8541), .o(n_8584) );
in01f80 g742679 ( .a(n_37414), .o(n_37415) );
in01f80 newInst_675 ( .a(newNet_674), .o(newNet_675) );
na02f80 g737671 ( .a(FE_OCPN887_n_42367), .b(n_42710), .o(n_42766) );
no02f80 g775296 ( .a(n_5809), .b(n_5808), .o(n_5832) );
in01f80 g746708 ( .a(n_33112), .o(n_33163) );
na02f80 g742594 ( .a(n_37505), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37557) );
no02f80 g752631 ( .a(n_28242), .b(n_28241), .o(n_28243) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_24_ ( .ck(newNet_1982), .d(n_12150), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_) );
in01f80 newInst_3557 ( .a(newNet_3556), .o(newNet_3557) );
na02f80 FE_RC_2768_0 ( .a(n_2627), .b(n_2688), .o(FE_RN_1179_0) );
in01f80 g752742 ( .a(n_44046), .o(n_27960) );
in01f80 newInst_1749 ( .a(newNet_1748), .o(newNet_1749) );
no02f80 FE_RC_2716_0 ( .a(FE_RN_1144_0), .b(FE_RN_1145_0), .o(n_44219) );
ao12f80 g780352 ( .a(n_873), .b(n_937), .c(n_872), .o(n_972) );
na02f80 g752388 ( .a(FE_OCP_RBN3313_delay_xor_ln22_unr18_stage7_stallmux_q_2_), .b(n_44722), .o(n_27777) );
in01f80 g739697 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n_40508) );
in01f80 g767010 ( .a(n_14137), .o(n_14138) );
in01f80 g751775 ( .a(n_29047), .o(n_29029) );
na02f80 g768923 ( .a(n_11842), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n_11843) );
in01f80 g767597 ( .a(n_13050), .o(n_13051) );
in01f80 FE_OCPC1403_n_21007 ( .a(n_21007), .o(FE_OCPN1403_n_21007) );
na02f80 g776798 ( .a(n_47010), .b(n_4231), .o(n_4404) );
in01f80 g764240 ( .a(n_16515), .o(n_16524) );
no02f80 g748141 ( .a(n_31929), .b(n_31868), .o(n_31930) );
na02f80 g739085 ( .a(n_41072), .b(n_40866), .o(n_41096) );
na02f80 g775706 ( .a(n_5335), .b(n_4017), .o(n_5411) );
in01f80 g771415 ( .a(n_9655), .o(n_9833) );
oa22f80 FE_RC_234_0 ( .a(n_14148), .b(FE_OCP_RBN2253_n_13017), .c(n_14149), .d(n_13418), .o(n_14321) );
ao12f80 g754446 ( .a(n_25239), .b(n_25568), .c(n_25398), .o(n_25634) );
oa22f80 g784419 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .c(n_36358), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46231) );
no02f80 g764747 ( .a(n_15938), .b(n_15937), .o(n_16031) );
no02f80 g744726 ( .a(n_35101), .b(n_30587), .o(n_35156) );
oa12f80 g737358 ( .a(n_42747), .b(n_42838), .c(n_42727), .o(n_42850) );
na03f80 g756845 ( .a(n_23335), .b(n_23313), .c(n_23031), .o(n_23336) );
in01f80 g756137 ( .a(n_24998), .o(n_25032) );
no03m80 FE_RC_583_0 ( .a(FE_RN_179_0), .b(n_23388), .c(n_23389), .o(n_47245) );
in01f80 g753686 ( .a(n_26584), .o(n_26617) );
in01f80 g749642 ( .a(n_31433), .o(n_31434) );
no02f80 g776622 ( .a(n_3963), .b(n_3082), .o(n_4111) );
in01f80 g752707 ( .a(n_28993), .o(n_28134) );
in01f80 newInst_2109 ( .a(newNet_2108), .o(newNet_2109) );
in01f80 FE_OCPC1051_n_31674 ( .a(FE_OCP_RBN3713_n_31466), .o(FE_OCPN1051_n_31674) );
no02f80 g748248 ( .a(FE_OCP_RBN3083_n_31819), .b(n_44437), .o(n_31931) );
na02f80 g743219 ( .a(n_36872), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_), .o(n_36917) );
no02f80 g738673 ( .a(n_41478), .b(n_41296), .o(n_41688) );
no02f80 FE_RC_2200_0 ( .a(n_26359), .b(FE_RN_790_0), .o(n_26390) );
no02f80 g743088 ( .a(n_36591), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37111) );
oa12f80 g750935 ( .a(n_28972), .b(n_28971), .c(n_28970), .o(n_29059) );
in01f80 FE_OCP_RBC2480_n_8595 ( .a(n_8595), .o(FE_OCP_RBN2480_n_8595) );
in01f80 g743213 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_5_), .o(n_36918) );
ao22s80 FE_RC_3881_0 ( .a(FE_OCP_DRV_N3158_n_27062), .b(FE_OCP_RBN1197_n_30619), .c(FE_OCPN1410_n_27014), .d(n_30619), .o(n_30727) );
in01f80 fopt782851 ( .a(n_44275), .o(n_44277) );
na02f80 g751444 ( .a(n_28491), .b(n_28489), .o(n_28507) );
na02f80 g761816 ( .a(n_18435), .b(n_18373), .o(n_18554) );
na02f80 g759665 ( .a(n_21878), .b(n_21877), .o(n_21879) );
no03m80 FE_RC_3576_0 ( .a(n_35752), .b(n_35696), .c(FE_RN_1554_0), .o(FE_RN_1555_0) );
na02f80 g774004 ( .a(n_6907), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .o(n_6987) );
no02f80 g765506 ( .a(FE_OFN765_n_15670), .b(n_15087), .o(n_15826) );
ao12f80 g739397 ( .a(n_40777), .b(FE_OCPN898_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n_41177) );
na02f80 g751303 ( .a(n_29675), .b(n_29132), .o(n_29712) );
in01f80 newInst_3276 ( .a(newNet_3275), .o(newNet_3276) );
in01f80 g758376 ( .a(n_22014), .o(n_22015) );
na02f80 g778422 ( .a(n_2602), .b(n_2666), .o(n_2695) );
no02f80 g741547 ( .a(n_38680), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38707) );
no02f80 g742734 ( .a(n_37350), .b(n_37052), .o(n_37351) );
in01f80 newInst_775 ( .a(newNet_774), .o(newNet_775) );
in01f80 g759260 ( .a(n_21011), .o(n_21080) );
ao12f80 g755310 ( .a(n_24884), .b(n_24883), .c(n_24897), .o(n_26587) );
in01f80 fopt783156 ( .a(n_40578), .o(n_44687) );
in01f80 newInst_1207 ( .a(newNet_1158), .o(newNet_1207) );
ao22s80 g779333 ( .a(n_1602), .b(n_1454), .c(FE_OCP_RBN2155_n_1602), .d(n_1453), .o(n_1658) );
na02f80 g774809 ( .a(n_6290), .b(FE_OCP_RBN2979_n_5656), .o(n_6352) );
na02f80 g754370 ( .a(n_25761), .b(n_25389), .o(n_25818) );
oa12f80 g740802 ( .a(n_38980), .b(n_39468), .c(n_39395), .o(n_39489) );
in01f80 newInst_658 ( .a(newNet_657), .o(newNet_658) );
ao12f80 g746772 ( .a(n_32899), .b(n_32924), .c(n_32898), .o(n_34137) );
in01f80 g745144 ( .a(n_35667), .o(n_34724) );
in01f80 g755340 ( .a(n_24861), .o(n_24877) );
ao22s80 FE_RC_3942_0 ( .a(FE_RN_1704_0), .b(n_16972), .c(FE_RN_1705_0), .d(n_16970), .o(n_17230) );
in01f80 g758467 ( .a(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .o(n_23254) );
na02f80 g776729 ( .a(n_4275), .b(n_3977), .o(n_4301) );
in01f80 g775569 ( .a(FE_OFN76_n_5397), .o(n_6263) );
na02f80 g750370 ( .a(n_29661), .b(n_29698), .o(n_29733) );
in01f80 newInst_161 ( .a(newNet_1), .o(newNet_161) );
na02f80 g763073 ( .a(n_17200), .b(n_17044), .o(n_17252) );
na02f80 g738056 ( .a(n_42100), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42121) );
na02f80 g777156 ( .a(n_5298), .b(n_5297), .o(n_5299) );
oa22f80 g746743 ( .a(n_33016), .b(n_32984), .c(n_33066), .d(n_32983), .o(n_33945) );
ao12f80 g737527 ( .a(n_42453), .b(n_42472), .c(n_42461), .o(n_42512) );
in01f80 FE_OCP_RBC2534_n_47018 ( .a(FE_OCP_RBN2533_n_47018), .o(FE_OCP_RBN2534_n_47018) );
na02f80 g762129 ( .a(n_18217), .b(n_18216), .o(n_18244) );
in01f80 g772312 ( .a(n_8727), .o(n_8728) );
in01f80 g742623 ( .a(n_37974), .o(n_37566) );
no02f80 g742444 ( .a(n_37732), .b(n_37529), .o(n_37752) );
na02f80 g757452 ( .a(FE_OCP_RBN3822_n_44061), .b(n_22939), .o(n_23015) );
ao12f80 g750413 ( .a(n_29608), .b(n_29607), .c(n_29606), .o(n_31197) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_12_ ( .ck(newNet_2317), .d(n_40403), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_) );
na02f80 g736570 ( .a(n_43450), .b(n_43518), .o(n_43571) );
no02f80 g738682 ( .a(n_41525), .b(n_41654), .o(n_41685) );
no02f80 g741568 ( .a(n_38651), .b(n_38648), .o(n_38671) );
in01f80 g749440 ( .a(n_30723), .o(n_30724) );
na02f80 g777106 ( .a(n_4675), .b(n_3606), .o(n_5384) );
na02f80 g751599 ( .a(FE_OCP_RBN3404_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .o(n_28698) );
ao12f80 g760341 ( .a(n_20159), .b(n_20212), .c(n_20211), .o(n_20226) );
na02f80 g756364 ( .a(n_24498), .b(n_23927), .o(n_24645) );
no02f80 g761954 ( .a(n_18966), .b(n_18736), .o(n_19020) );
no02f80 g765378 ( .a(n_16135), .b(n_15566), .o(n_15633) );
in01f80 g763958 ( .a(n_16686), .o(n_16658) );
no02f80 g776145 ( .a(n_4944), .b(n_4490), .o(n_5077) );
na02f80 g770161 ( .a(n_10847), .b(n_10820), .o(n_10950) );
na02f80 g741608 ( .a(n_38613), .b(n_38625), .o(n_38658) );
in01f80 newInst_491 ( .a(newNet_490), .o(newNet_491) );
ao12f80 g773909 ( .a(n_6981), .b(n_6980), .c(n_6979), .o(n_7044) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_1_ ( .ck(newNet_382), .d(n_40589), .o(delay_xor_ln22_unr28_stage10_stallmux_q_1_) );
no02f80 g737566 ( .a(n_42266), .b(n_42210), .o(n_42265) );
na02f80 g778179 ( .a(n_2906), .b(n_2831), .o(n_3068) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_24_ ( .ck(newNet_229), .d(n_46191), .o(delay_xor_ln22_unr6_stage3_stallmux_q_24_) );
na02f80 g738336 ( .a(n_41795), .b(FE_OCP_RBN2316_n_41420), .o(n_41831) );
na02f80 g767983 ( .a(n_13115), .b(n_12988), .o(n_13671) );
oa12f80 g773804 ( .a(n_7210), .b(n_7209), .c(n_7208), .o(n_8114) );
oa12f80 g780255 ( .a(n_911), .b(n_910), .c(n_1159), .o(n_1025) );
ao12f80 g744109 ( .a(n_35490), .b(n_35556), .c(n_35515), .o(n_35574) );
in01f80 g739967 ( .a(n_40122), .o(n_40159) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_20_ ( .ck(newNet_1116), .d(n_10913), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_) );
in01f80 g747582 ( .a(n_33397), .o(n_33375) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_16_ ( .ck(newNet_2111), .d(n_6105), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_) );
na02f80 g778347 ( .a(n_2627), .b(n_2626), .o(n_2689) );
in01f80 FE_RC_2633_0 ( .a(n_11693), .o(FE_RN_1097_0) );
oa12f80 g771159 ( .a(n_9816), .b(n_9884), .c(n_9815), .o(n_9917) );
no03m80 FE_RC_1066_0 ( .a(n_37040), .b(FE_RN_314_0), .c(n_37395), .o(n_37467) );
in01f80 g757551 ( .a(n_22823), .o(n_22824) );
in01f80 FE_OCP_RBC3399_n_12751 ( .a(n_12751), .o(FE_OCP_RBN3399_n_12751) );
in01f80 FE_OCP_RBC2833_n_26081 ( .a(n_26081), .o(FE_OCP_RBN2833_n_26081) );
na02f80 g741878 ( .a(n_38407), .b(n_38406), .o(n_38408) );
no02f80 g753763 ( .a(n_26424), .b(n_23564), .o(n_26521) );
in01f80 newInst_835 ( .a(newNet_144), .o(newNet_835) );
no02f80 g749362 ( .a(n_30601), .b(n_30370), .o(n_30627) );
in01f80 g768235 ( .a(n_12753), .o(n_12677) );
in01f80 g759089 ( .a(n_21226), .o(n_21278) );
in01f80 newInst_1301 ( .a(newNet_1300), .o(newNet_1301) );
in01f80 FE_OFC773_n_46137 ( .a(n_46137), .o(FE_OFN773_n_46137) );
ao22s80 g743065 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .c(n_36991), .d(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37524) );
no02f80 g763672 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .o(n_17663) );
in01f80 newInst_1127 ( .a(newNet_887), .o(newNet_1127) );
in01f80 newInst_2207 ( .a(newNet_2206), .o(newNet_2207) );
in01f80 g769870 ( .a(n_11083), .o(n_11084) );
in01f80 g746095 ( .a(n_33957), .o(n_33941) );
in01f80 g751691 ( .a(n_28447), .o(n_28458) );
no02f80 g772862 ( .a(n_8051), .b(n_8050), .o(n_8102) );
in01f80 g767672 ( .a(n_13260), .o(n_13261) );
in01f80 FE_OCPC945_n_1780 ( .a(n_1780), .o(FE_OCPN945_n_1780) );
in01f80 FE_OCP_RBC3506_n_13860 ( .a(FE_OCP_RBN2388_n_13860), .o(FE_OCP_RBN3506_n_13860) );
na02f80 g753976 ( .a(FE_OCP_RBN3682_n_26171), .b(FE_OCP_RBN2833_n_26081), .o(n_26250) );
no02f80 g748798 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n_32425) );
in01f80 g746795 ( .a(n_32974), .o(n_32975) );
in01f80 g756668 ( .a(n_23606), .o(n_23599) );
na02f80 g775778 ( .a(n_5547), .b(n_5502), .o(n_5563) );
no02f80 g741067 ( .a(n_38891), .b(FE_OCP_RBN2549_n_44944), .o(n_38962) );
na02f80 g767958 ( .a(n_12994), .b(n_12916), .o(n_12995) );
in01f80 g745058 ( .a(n_36386), .o(n_36356) );
in01f80 newInst_736 ( .a(newNet_735), .o(newNet_736) );
ao12f80 g755376 ( .a(n_24833), .b(n_24832), .c(n_24834), .o(n_26530) );
no02f80 FE_RC_2203_0 ( .a(n_26412), .b(n_26337), .o(FE_RN_792_0) );
no02f80 g738079 ( .a(n_42051), .b(n_42196), .o(n_42075) );
no02f80 g772679 ( .a(n_8264), .b(n_8313), .o(n_8344) );
in01f80 g777638 ( .a(n_3470), .o(n_3471) );
oa12f80 g766513 ( .a(n_13948), .b(n_14027), .c(FE_OCP_RBN2246_n_13017), .o(n_14104) );
no02f80 g771252 ( .a(n_9314), .b(n_9298), .o(n_9509) );
in01f80 g769856 ( .a(FE_OCP_RBN3006_n_11087), .o(n_11112) );
in01f80 g764954 ( .a(n_15584), .o(n_15585) );
in01f80 g777916 ( .a(n_3133), .o(n_3120) );
na02f80 g769282 ( .a(FE_OCP_RBN3093_n_11475), .b(n_10797), .o(n_11580) );
in01f80 FE_OCP_RBC2732_n_4219 ( .a(FE_OCP_RBN2728_n_4219), .o(FE_OCP_RBN2732_n_4219) );
in01f80 g757252 ( .a(n_23170), .o(n_23171) );
in01f80 g738006 ( .a(n_42202), .o(n_42201) );
in01f80 g753927 ( .a(n_26320), .o(n_26321) );
na02f80 g769886 ( .a(n_10967), .b(n_10939), .o(n_11089) );
in01f80 g759499 ( .a(n_20932), .o(n_20933) );
no02f80 FE_RC_1786_0 ( .a(n_28018), .b(n_28050), .o(FE_RN_524_0) );
no02f80 g736559 ( .a(n_43532), .b(n_43152), .o(n_43573) );
no02f80 g769431 ( .a(n_11355), .b(n_11336), .o(n_11439) );
ao12f80 g741453 ( .a(n_38684), .b(n_38788), .c(n_38778), .o(n_38796) );
oa22f80 g780118 ( .a(n_1175), .b(FE_OFN761_n_45813), .c(n_1176), .d(n_1203), .o(n_1205) );
no02f80 g753719 ( .a(n_26531), .b(n_26530), .o(n_26658) );
in01f80 g738618 ( .a(n_41405), .o(n_41507) );
na02f80 g775178 ( .a(n_5818), .b(n_4556), .o(n_5815) );
in01f80 g768615 ( .a(n_12289), .o(n_12290) );
in01f80 FE_OCP_RBC3535_n_13765 ( .a(FE_OCP_RBN3531_n_13765), .o(FE_OCP_RBN3535_n_13765) );
no02f80 g741043 ( .a(n_38885), .b(n_38930), .o(n_38931) );
in01f80 newInst_374 ( .a(newNet_302), .o(newNet_374) );
na02f80 g748430 ( .a(n_31730), .b(n_30933), .o(n_31722) );
oa22f80 FE_RC_3518_0 ( .a(n_23017), .b(FE_OCPN1022_n_23195), .c(FE_RN_1519_0), .d(n_23212), .o(n_23266) );
no02f80 FE_RC_1802_0 ( .a(n_24217), .b(n_25239), .o(FE_RN_533_0) );
in01f80 g764531 ( .a(n_16086), .o(n_16117) );
na02f80 g781017 ( .a(sin_out_21), .b(FE_OFN3_n_43918), .o(n_290) );
in01f80 FE_OCP_RBC3397_n_37624 ( .a(n_37624), .o(FE_OCP_RBN3397_n_37624) );
in01f80 g768388 ( .a(n_12479), .o(n_12480) );
no02f80 g753626 ( .a(n_26583), .b(n_23590), .o(n_26666) );
no02f80 g750924 ( .a(n_30068), .b(n_30289), .o(n_30333) );
oa22f80 FE_RC_659_0 ( .a(n_6690), .b(n_6960), .c(n_6961), .d(n_6689), .o(n_7050) );
in01f80 g751862 ( .a(n_28210), .o(n_28211) );
oa12f80 g743856 ( .a(n_35672), .b(n_35671), .c(n_35670), .o(n_35757) );
in01f80 FE_OCPC975_n_46956 ( .a(FE_OCPN974_n_46956), .o(FE_OCPN975_n_46956) );
no02f80 g768328 ( .a(n_12469), .b(n_12468), .o(n_12502) );
oa22f80 g776000 ( .a(n_4784), .b(n_4182), .c(FE_OCP_RBN2841_n_4784), .d(FE_OCPN846_n_4046), .o(n_4959) );
na02f80 g772323 ( .a(n_8491), .b(FE_OCP_RBN3463_n_7886), .o(n_8528) );
na02f80 g775109 ( .a(n_6016), .b(n_5934), .o(n_6077) );
no02f80 g757946 ( .a(n_22133), .b(n_44277), .o(n_22235) );
no02f80 g749481 ( .a(n_30530), .b(n_30171), .o(n_30531) );
na02f80 g743020 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_30_), .o(n_37068) );
na02f80 g751634 ( .a(n_28421), .b(n_28388), .o(n_28658) );
no02f80 g777847 ( .a(n_3261), .b(n_3155), .o(n_3276) );
na02f80 g753175 ( .a(n_27103), .b(n_25596), .o(n_27157) );
na02f80 g738949 ( .a(n_41244), .b(n_41243), .o(n_41245) );
na02f80 g752827 ( .a(n_27272), .b(n_27206), .o(n_27402) );
in01f80 FE_RC_2122_0 ( .a(n_20836), .o(FE_RN_738_0) );
no02f80 g764737 ( .a(n_15847), .b(n_14524), .o(n_15849) );
na02f80 g761910 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .o(n_18914) );
oa22f80 g756152 ( .a(n_24145), .b(n_23790), .c(n_24147), .d(n_23791), .o(n_24178) );
oa12f80 g768860 ( .a(n_11657), .b(n_44356), .c(n_11647), .o(n_11913) );
in01f80 newInst_1279 ( .a(newNet_1278), .o(newNet_1279) );
no02f80 g781292 ( .a(beta_31), .b(beta_25), .o(n_52) );
na02f80 g765895 ( .a(n_15032), .b(n_14966), .o(n_14967) );
in01f80 newInst_65 ( .a(newNet_8), .o(newNet_65) );
na02f80 g776324 ( .a(n_4786), .b(n_4756), .o(n_4757) );
in01f80 FE_RC_2906_0 ( .a(n_9402), .o(FE_RN_1262_0) );
in01f80 g748420 ( .a(n_31704), .o(n_31727) );
na02f80 g764432 ( .a(n_16088), .b(n_14618), .o(n_16127) );
ao22s80 g780860 ( .a(n_420), .b(n_476), .c(n_403), .d(n_260), .o(n_477) );
in01f80 FE_OCPC956_n_39096 ( .a(FE_OCP_RBN2685_n_38870), .o(FE_OCPN956_n_39096) );
in01f80 newInst_1987 ( .a(newNet_1671), .o(newNet_1987) );
in01f80 g772640 ( .a(n_8321), .o(n_8348) );
na02f80 FE_RC_3973_0 ( .a(n_24592), .b(FE_RN_1720_0), .o(n_24779) );
oa12f80 g736353 ( .a(n_340), .b(n_43774), .c(FE_OFN3_n_43918), .o(n_43813) );
in01f80 newInst_1632 ( .a(newNet_1631), .o(newNet_1632) );
in01f80 g740136 ( .a(n_39802), .o(n_39820) );
no02f80 g762093 ( .a(n_18196), .b(n_18179), .o(n_18180) );
no02f80 g749079 ( .a(n_30978), .b(n_29555), .o(n_31093) );
no02f80 g771993 ( .a(n_44575), .b(n_7862), .o(n_9218) );
oa12f80 g745725 ( .a(n_34054), .b(n_34053), .c(n_34069), .o(n_35500) );
oa12f80 g743881 ( .a(n_36979), .b(n_36774), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37814) );
no02f80 g751002 ( .a(n_30438), .b(n_30164), .o(n_31041) );
oa22f80 FE_RC_536_0 ( .a(n_28732), .b(n_29117), .c(n_28733), .d(n_29116), .o(n_29217) );
in01f80 g764518 ( .a(n_16053), .o(n_16089) );
in01f80 FE_OCP_RBC2394_n_8288 ( .a(FE_OCP_RBN2393_n_8288), .o(FE_OCP_RBN2394_n_8288) );
ao12f80 g773658 ( .a(n_7266), .b(n_7267), .c(n_7265), .o(n_7345) );
no02f80 g775966 ( .a(n_5243), .b(n_5242), .o(n_5353) );
na02f80 g756919 ( .a(n_24025), .b(n_24024), .o(n_24026) );
na02f80 g740577 ( .a(n_39616), .b(n_39615), .o(n_39643) );
in01f80 FE_OCP_RBC2996_n_11004 ( .a(n_11004), .o(FE_OCP_RBN2996_n_11004) );
in01f80 newInst_2098 ( .a(newNet_2097), .o(newNet_2098) );
na02f80 g775286 ( .a(n_5718), .b(n_4556), .o(n_5772) );
na02f80 FE_RC_4163_0 ( .a(FE_RN_1813_0), .b(n_33501), .o(n_33518) );
na02f80 g773915 ( .a(n_6934), .b(n_5362), .o(n_7036) );
no02f80 g743454 ( .a(n_36538), .b(n_36554), .o(n_36612) );
na02f80 g777958 ( .a(n_3081), .b(n_3064), .o(n_3149) );
na02f80 g745453 ( .a(n_34512), .b(n_34566), .o(n_34626) );
no02f80 g764382 ( .a(n_16316), .b(n_16266), .o(n_16418) );
in01f80 g767509 ( .a(n_14733), .o(n_14896) );
na02f80 g744649 ( .a(n_36558), .b(n_36018), .o(n_36603) );
in01f80 g779940 ( .a(FE_OCP_RBN3242_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1800) );
in01f80 g780894 ( .a(n_389), .o(n_390) );
oa12f80 g779286 ( .a(n_1700), .b(n_1699), .c(n_1698), .o(n_2463) );
na02f80 g747103 ( .a(n_32927), .b(delay_add_ln22_unr20_stage8_stallmux_q_8_), .o(n_32988) );
na02f80 g763157 ( .a(n_17049), .b(n_16908), .o(n_17145) );
no02f80 g746691 ( .a(n_33328), .b(n_33253), .o(n_33329) );
in01f80 newInst_3434 ( .a(newNet_3433), .o(newNet_3434) );
na02f80 g773462 ( .a(n_7465), .b(n_7501), .o(n_7513) );
no02f80 g737322 ( .a(n_42879), .b(n_42487), .o(n_42891) );
in01f80 g739915 ( .a(n_40164), .o(n_40165) );
na02f80 g775523 ( .a(n_5522), .b(n_5488), .o(n_5651) );
na02f80 g736806 ( .a(n_43297), .b(n_46936), .o(n_43314) );
in01f80 g742538 ( .a(n_37597), .o(n_37596) );
in01f80 newInst_1736 ( .a(newNet_1613), .o(newNet_1736) );
na02f80 g750670 ( .a(n_29415), .b(n_29393), .o(n_29491) );
in01f80 g781348 ( .a(beta_1), .o(n_353) );
no02f80 g750435 ( .a(n_29590), .b(n_28476), .o(n_29611) );
no02f80 g772803 ( .a(n_8073), .b(n_47241), .o(n_8133) );
na02f80 g751055 ( .a(n_29932), .b(n_30033), .o(n_30062) );
in01f80 FE_OCPC1862_n_30319 ( .a(FE_OCPN1861_n_30319), .o(FE_OCPN1862_n_30319) );
in01f80 g754255 ( .a(n_25983), .o(n_25984) );
ao12f80 g738173 ( .a(n_41858), .b(n_41995), .c(n_41810), .o(n_41996) );
in01f80 g739933 ( .a(n_40374), .o(n_40371) );
na02f80 g759316 ( .a(n_21754), .b(n_21299), .o(n_21801) );
na02f80 g760936 ( .a(n_19383), .b(n_19422), .o(n_19506) );
in01f80 g769424 ( .a(n_11455), .o(n_11585) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_30_ ( .ck(newNet_2721), .d(n_17725), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_) );
na02f80 g778592 ( .a(n_2384), .b(n_2423), .o(n_2691) );
no02f80 g768050 ( .a(n_12790), .b(n_12850), .o(n_12882) );
na02f80 g736698 ( .a(n_43432), .b(n_43358), .o(n_43468) );
no02f80 g743704 ( .a(n_36279), .b(n_35641), .o(n_36327) );
na02f80 g742217 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37967), .o(n_38271) );
na02f80 g770268 ( .a(n_10776), .b(n_10775), .o(n_10777) );
in01f80 newInst_3628 ( .a(newNet_585), .o(newNet_3628) );
na02f80 g754547 ( .a(n_26606), .b(n_26605), .o(n_26607) );
na02f80 g740018 ( .a(n_39981), .b(FE_OCP_RBN3052_n_39913), .o(n_40044) );
no03m80 FE_RC_775_0 ( .a(n_11283), .b(n_11158), .c(n_11215), .o(n_11285) );
no02f80 FE_RC_3502_0 ( .a(FE_RN_1510_0), .b(FE_RN_1511_0), .o(n_27661) );
no02f80 g757018 ( .a(n_23803), .b(n_23746), .o(n_24169) );
no02f80 g750953 ( .a(n_30811), .b(n_30089), .o(n_30167) );
in01f80 g773279 ( .a(n_7712), .o(n_7730) );
in01f80 FE_OCP_RBC2601_n_34388 ( .a(FE_OCP_RBN2599_n_34388), .o(FE_OCP_RBN2601_n_34388) );
na02f80 g756817 ( .a(n_24006), .b(n_23950), .o(n_24032) );
in01f80 newInst_157 ( .a(newNet_156), .o(newNet_157) );
no02f80 g770594 ( .a(n_10356), .b(n_10407), .o(n_10529) );
in01f80 g747213 ( .a(n_32851), .o(n_32830) );
in01f80 g750723 ( .a(n_29271), .o(n_29272) );
na02f80 g749269 ( .a(n_30765), .b(n_30272), .o(n_30800) );
ao12f80 g777899 ( .a(n_2907), .b(n_3114), .c(n_2963), .o(n_3176) );
oa22f80 g745791 ( .a(n_44112), .b(n_34004), .c(n_44102), .d(n_33976), .o(n_34423) );
na02f80 g749072 ( .a(n_30991), .b(n_27366), .o(n_30992) );
in01f80 FE_OCP_RBC2493_n_8508 ( .a(n_8508), .o(FE_OCP_RBN2493_n_8508) );
in01f80 g760283 ( .a(n_20299), .o(n_20300) );
no02f80 g744640 ( .a(n_35256), .b(n_35213), .o(n_35257) );
na02f80 g766667 ( .a(n_13730), .b(n_12864), .o(n_13815) );
in01f80 g753316 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_7_), .o(n_28227) );
in01f80 newInst_336 ( .a(newNet_335), .o(newNet_336) );
no02f80 g757414 ( .a(n_22869), .b(n_22870), .o(n_22965) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_17_ ( .ck(newNet_734), .d(n_46147), .o(delay_xor_ln21_unr6_stage3_stallmux_q_17_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_10_ ( .ck(newNet_1433), .d(n_36453), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_) );
in01f80 FE_OCP_DRV_C1601_n_21639 ( .a(n_21639), .o(FE_OCP_DRV_N1601_n_21639) );
na02f80 g744828 ( .a(n_35065), .b(n_35037), .o(n_35207) );
na02f80 g767612 ( .a(n_12949), .b(n_12942), .o(n_12943) );
no02f80 g750690 ( .a(n_29161), .b(n_29266), .o(n_29325) );
in01f80 g760831 ( .a(n_19615), .o(n_19653) );
in01f80 g780789 ( .a(n_553), .o(n_554) );
in01f80 g752453 ( .a(n_27729), .o(n_27755) );
no03m80 g778497 ( .a(n_2721), .b(n_2729), .c(n_2803), .o(n_2804) );
na02f80 g737915 ( .a(n_42270), .b(n_41886), .o(n_42496) );
na02f80 g774984 ( .a(n_6129), .b(n_6143), .o(n_6243) );
in01f80 g770953 ( .a(n_10162), .o(n_10163) );
na02f80 g773995 ( .a(n_6913), .b(n_6890), .o(n_6990) );
na02f80 g753122 ( .a(n_27216), .b(n_27217), .o(n_27263) );
oa12f80 g746404 ( .a(n_33057), .b(n_33484), .c(n_33449), .o(n_33520) );
oa22f80 g752441 ( .a(n_27693), .b(n_24059), .c(n_27666), .d(n_27845), .o(n_27731) );
no02f80 g736642 ( .a(n_43413), .b(n_43215), .o(n_43414) );
na02f80 g753550 ( .a(n_26670), .b(n_26620), .o(n_26704) );
in01f80 g740782 ( .a(n_39891), .o(n_39513) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_20_ ( .ck(newNet_237), .d(n_46185), .o(delay_xor_ln22_unr6_stage3_stallmux_q_20_) );
na02f80 g778621 ( .a(n_2438), .b(n_2473), .o(n_2474) );
in01f80 g768899 ( .a(n_11850), .o(n_11870) );
in01f80 FE_OCP_RBC1992_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_ ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(FE_OCP_RBN1992_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
in01f80 FE_OCP_RBC1911_n_20545 ( .a(FE_OCP_RBN1909_n_20545), .o(FE_OCP_RBN1911_n_20545) );
in01f80 g780681 ( .a(n_662), .o(n_663) );
in01f80 g767532 ( .a(n_13154), .o(n_13185) );
in01f80 newInst_2143 ( .a(newNet_2142), .o(newNet_2143) );
in01f80 g761857 ( .a(n_20135), .o(n_20136) );
oa12f80 g776871 ( .a(n_4119), .b(n_4118), .c(FE_OFN78_n_4117), .o(n_4180) );
ao12f80 g757908 ( .a(n_22926), .b(n_22784), .c(n_22725), .o(n_22979) );
na02f80 g754464 ( .a(n_25601), .b(n_25321), .o(n_25654) );
na02f80 g774802 ( .a(n_45475), .b(n_5636), .o(n_6367) );
in01f80 g749413 ( .a(n_31977), .o(n_31978) );
oa12f80 g764807 ( .a(n_15219), .b(n_15589), .c(n_15144), .o(n_15698) );
in01f80 g749255 ( .a(n_30766), .o(n_30767) );
in01f80 g748169 ( .a(n_32210), .o(n_32211) );
na02f80 g741646 ( .a(n_38556), .b(n_38575), .o(n_38601) );
no02f80 g750608 ( .a(n_29421), .b(FE_OCPN1746_n_29420), .o(n_29498) );
in01f80 FE_OCP_RBC3423_n_37794 ( .a(n_37794), .o(FE_OCP_RBN3423_n_37794) );
no02f80 g771445 ( .a(n_9399), .b(n_9522), .o(n_9608) );
oa12f80 g768851 ( .a(n_12089), .b(n_12088), .c(n_12087), .o(n_12221) );
ao12f80 g776386 ( .a(n_3841), .b(n_4054), .c(n_3928), .o(n_4197) );
in01f80 FE_OCP_RBC2600_n_34388 ( .a(FE_OCP_RBN2599_n_34388), .o(FE_OCP_RBN2600_n_34388) );
ao22s80 g736266 ( .a(n_43894), .b(n_43539), .c(n_43895), .d(n_43540), .o(n_43912) );
in01f80 FE_OCP_RBC2698_n_4238 ( .a(n_4238), .o(FE_OCP_RBN2698_n_4238) );
no02f80 g770280 ( .a(n_10573), .b(n_8865), .o(n_10574) );
na02f80 FE_RC_4241_0 ( .a(FE_RN_1862_0), .b(FE_RN_1863_0), .o(FE_RN_1864_0) );
no02f80 FE_RC_1758_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .b(n_11973), .o(FE_RN_500_0) );
in01f80 g769145 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n_11696) );
na02f80 g749681 ( .a(n_31482), .b(n_31540), .o(n_31541) );
ao12f80 g743745 ( .a(n_37294), .b(n_36557), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37342) );
in01f80 newInst_1140 ( .a(newNet_1139), .o(newNet_1140) );
no02f80 g739467 ( .a(FE_OCPN898_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n_41107) );
in01f80 g773568 ( .a(n_7683), .o(n_8389) );
no02f80 g753663 ( .a(n_26562), .b(FE_OCP_RBN2981_n_26591), .o(n_26590) );
na02f80 FE_RC_2129_0 ( .a(n_15035), .b(n_15124), .o(FE_RN_743_0) );
in01f80 newInst_1436 ( .a(newNet_1435), .o(newNet_1436) );
oa12f80 g771789 ( .a(n_8682), .b(n_8751), .c(n_8661), .o(n_8848) );
na02f80 g779129 ( .a(n_1950), .b(n_1814), .o(n_1943) );
in01f80 g778614 ( .a(n_2814), .o(n_2781) );
na02f80 g750081 ( .a(n_29896), .b(n_29501), .o(n_30272) );
in01f80 newInst_1760 ( .a(newNet_200), .o(newNet_1760) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_21_ ( .ck(newNet_1115), .d(n_10981), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_) );
in01f80 g763752 ( .a(n_16801), .o(n_16802) );
na02f80 FE_RC_1727_0 ( .a(FE_RN_477_0), .b(n_23393), .o(FE_RN_478_0) );
in01f80 newInst_254 ( .a(newNet_253), .o(newNet_254) );
in01f80 g754347 ( .a(n_25849), .o(n_25850) );
in01f80 g738428 ( .a(n_41812), .o(n_41813) );
no02f80 g755103 ( .a(n_25201), .b(n_24093), .o(n_25292) );
in01f80 FE_RC_345_0 ( .a(n_11643), .o(FE_RN_99_0) );
in01f80 newInst_1806 ( .a(newNet_1805), .o(newNet_1806) );
oa12f80 g770771 ( .a(n_10219), .b(n_10218), .c(n_10217), .o(n_10295) );
in01f80 newInst_1249 ( .a(newNet_1248), .o(newNet_1249) );
no02f80 g773074 ( .a(n_7961), .b(n_8038), .o(n_8048) );
no02f80 g755392 ( .a(n_24726), .b(n_24788), .o(n_24729) );
in01f80 g749845 ( .a(n_31066), .o(n_31067) );
na02f80 g740559 ( .a(n_39630), .b(n_45841), .o(n_39654) );
ao12f80 g766233 ( .a(n_14171), .b(n_14780), .c(n_14213), .o(n_14839) );
na02f80 g759708 ( .a(n_20612), .b(n_20500), .o(n_20638) );
na02f80 g737315 ( .a(n_42850), .b(n_42756), .o(n_42875) );
na02f80 g737074 ( .a(FE_OCPN912_n_43022), .b(n_42794), .o(n_43164) );
in01f80 g749042 ( .a(n_31001), .o(n_31002) );
in01f80 g780636 ( .a(n_768), .o(n_769) );
na02f80 g740544 ( .a(n_39706), .b(n_39693), .o(n_39714) );
no02f80 FE_RC_2223_0 ( .a(n_32857), .b(FE_RN_805_0), .o(FE_RN_806_0) );
na02f80 g759950 ( .a(n_21691), .b(n_21720), .o(n_21824) );
oa22f80 g780016 ( .a(n_1263), .b(n_1072), .c(n_1262), .d(n_1073), .o(n_1273) );
in01f80 newInst_533 ( .a(newNet_532), .o(newNet_533) );
na02f80 g767640 ( .a(n_12746), .b(n_12520), .o(n_12804) );
in01f80 g738530 ( .a(n_41640), .o(n_41579) );
no02f80 g773451 ( .a(n_7583), .b(n_7563), .o(n_7881) );
in01f80 g757531 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .o(n_22754) );
na02f80 g771530 ( .a(n_9268), .b(n_9330), .o(n_9339) );
no02f80 g744274 ( .a(n_44180), .b(n_34966), .o(n_35736) );
na02f80 g755429 ( .a(n_25526), .b(n_25525), .o(n_25527) );
no02f80 FE_RC_1112_0 ( .a(FE_RN_334_0), .b(FE_RN_333_0), .o(FE_RN_335_0) );
in01f80 FE_OCP_RBC2574_n_34822 ( .a(n_34822), .o(FE_OCP_RBN2574_n_34822) );
oa22f80 g779851 ( .a(n_44652), .b(n_1124), .c(n_44637), .d(n_1100), .o(n_1303) );
no02f80 g747388 ( .a(n_32704), .b(n_32475), .o(n_32572) );
no02f80 g766707 ( .a(n_13759), .b(n_13776), .o(n_13860) );
na02f80 g757388 ( .a(n_22945), .b(n_22944), .o(n_22970) );
in01f80 newInst_1047 ( .a(newNet_564), .o(newNet_1047) );
na02f80 g766227 ( .a(n_14254), .b(FE_OCP_RBN2231_n_13141), .o(n_14378) );
in01f80 g779051 ( .a(n_2097), .o(n_2098) );
in01f80 g769287 ( .a(n_11478), .o(n_11598) );
no02f80 g778441 ( .a(n_2337), .b(n_1963), .o(n_2430) );
na02f80 g760703 ( .a(n_19688), .b(FE_OCPUNCON1804_n_18111), .o(n_19739) );
no02f80 g767757 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .o(n_13278) );
in01f80 g769376 ( .a(n_12007), .o(n_12008) );
in01f80 g760294 ( .a(n_20518), .o(n_20519) );
in01f80 newInst_3296 ( .a(newNet_3245), .o(newNet_3296) );
na02f80 g754567 ( .a(n_26709), .b(n_26708), .o(n_26736) );
in01f80 g743242 ( .a(n_36867), .o(n_36894) );
na02f80 g740275 ( .a(n_40169), .b(n_40170), .o(n_40210) );
na02f80 g763746 ( .a(n_16669), .b(n_16662), .o(n_16709) );
in01f80 g743735 ( .a(n_36208), .o(n_36248) );
no02f80 g776788 ( .a(n_4113), .b(n_3938), .o(n_4256) );
oa12f80 g745133 ( .a(n_34348), .b(n_34820), .c(n_34764), .o(n_34848) );
in01f80 g770115 ( .a(n_10906), .o(n_10907) );
no02f80 g750335 ( .a(n_29716), .b(FE_OCPN1768_n_29715), .o(n_29728) );
in01f80 FE_OCP_RBC2751_n_15239 ( .a(n_15239), .o(FE_OCP_RBN2751_n_15239) );
na02f80 g769335 ( .a(FE_OCP_RBN2001_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .o(n_11525) );
in01f80 FE_OCP_RBC2503_n_13896 ( .a(FE_OCP_RBN3528_n_13765), .o(FE_OCP_RBN2503_n_13896) );
in01f80 FE_OCP_RBC2335_n_24359 ( .a(n_24359), .o(FE_OCP_RBN2335_n_24359) );
in01f80 g779253 ( .a(n_1812), .o(n_1807) );
in01f80 g773897 ( .a(n_7045), .o(n_7046) );
no02f80 g771460 ( .a(n_9245), .b(n_9074), .o(n_9274) );
in01f80 g743498 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_26_), .o(n_36610) );
in01f80 g742693 ( .a(n_37889), .o(n_38251) );
no02f80 g764250 ( .a(n_46426), .b(n_16293), .o(n_16716) );
oa12f80 g749808 ( .a(n_31284), .b(FE_OCP_RBN3011_n_31117), .c(n_31216), .o(n_31623) );
no02f80 g755237 ( .a(n_25660), .b(n_25641), .o(n_25642) );
no02f80 g749850 ( .a(n_31064), .b(n_30103), .o(n_31114) );
na02f80 g764195 ( .a(n_16401), .b(n_16490), .o(n_16530) );
oa12f80 g749895 ( .a(FE_OCP_RBN3019_n_31117), .b(n_31251), .c(n_31253), .o(n_31276) );
na02f80 g768007 ( .a(n_12613), .b(n_11492), .o(n_12664) );
na02f80 g746637 ( .a(n_33205), .b(n_33065), .o(n_33206) );
in01f80 g761940 ( .a(n_18398), .o(n_18472) );
in01f80 g750529 ( .a(n_29530), .o(n_29501) );
no02f80 g748593 ( .a(n_31364), .b(n_31337), .o(n_31446) );
in01f80 fopt783921 ( .a(n_36508), .o(n_45625) );
na02f80 g764493 ( .a(FE_OCP_RBN1133_n_16041), .b(n_14650), .o(n_16119) );
in01f80 g746823 ( .a(n_33080), .o(n_33081) );
na02f80 g748324 ( .a(n_31521), .b(n_31500), .o(n_31556) );
in01f80 g770898 ( .a(n_9978), .o(n_10010) );
no02f80 g738745 ( .a(n_41355), .b(n_41372), .o(n_41361) );
no02f80 g775404 ( .a(n_5543), .b(n_4182), .o(n_5586) );
na03f80 FE_RC_503_0 ( .a(n_27802), .b(n_27868), .c(n_27777), .o(n_27919) );
in01f80 FE_RC_995_0 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .o(FE_RN_285_0) );
na02f80 g737712 ( .a(n_42394), .b(n_42391), .o(n_42446) );
in01f80 g743403 ( .a(n_36655), .o(n_36656) );
oa12f80 g749731 ( .a(n_29828), .b(n_29875), .c(n_29784), .o(n_29970) );
in01f80 g756448 ( .a(n_25002), .o(n_24258) );
oa22f80 FE_RC_721_0 ( .a(n_45511), .b(n_40631), .c(n_40601), .d(n_40632), .o(n_40663) );
in01f80 g775070 ( .a(n_6112), .o(n_6113) );
no02f80 g763739 ( .a(n_17574), .b(n_17573), .o(n_18350) );
na02f80 g760747 ( .a(n_19603), .b(n_19322), .o(n_19673) );
ao12f80 g755280 ( .a(n_24940), .b(n_24939), .c(n_24938), .o(n_25013) );
in01f80 g751534 ( .a(n_28673), .o(n_28721) );
in01f80 FE_OCP_RBC3704_n_26231 ( .a(FE_OCP_RBN3703_n_26231), .o(FE_OCP_RBN3704_n_26231) );
oa12f80 g745435 ( .a(n_34198), .b(n_34298), .c(n_34247), .o(n_34326) );
in01f80 g758028 ( .a(n_22381), .o(n_22382) );
no02f80 g774619 ( .a(n_6247), .b(n_6486), .o(n_6499) );
in01f80 g739876 ( .a(n_40432), .o(n_40412) );
in01f80 g767945 ( .a(n_13255), .o(n_13167) );
no02f80 g739326 ( .a(n_45147), .b(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n_40750) );
in01f80 FE_OFC744_n_23604 ( .a(n_23604), .o(FE_OFN744_n_23604) );
in01f80 newInst_1565 ( .a(newNet_765), .o(newNet_1565) );
na02f80 g774115 ( .a(n_6867), .b(n_6782), .o(n_6936) );
ao12f80 g768267 ( .a(n_11974), .b(n_12573), .c(n_11894), .o(n_12602) );
na02f80 g766420 ( .a(n_14127), .b(n_13437), .o(n_14128) );
no02f80 g764616 ( .a(n_16080), .b(n_15856), .o(n_15998) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_0_ ( .ck(newNet_1045), .d(n_16633), .o(n_44847) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_3_ ( .ck(newNet_2913), .d(n_4679), .o(delay_add_ln22_unr5_stage3_stallmux_q_3_) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_0_ ( .ck(newNet_2981), .d(n_4180), .o(delay_add_ln22_unr5_stage3_stallmux_q_0_) );
na02f80 g737048 ( .a(n_43103), .b(n_43102), .o(n_43127) );
ao12f80 g753691 ( .a(n_26815), .b(n_27135), .c(n_26710), .o(n_27201) );
oa12f80 g776410 ( .a(n_4709), .b(n_4708), .c(n_4710), .o(n_4793) );
na02f80 g736868 ( .a(n_43400), .b(n_43454), .o(n_43539) );
no02f80 g736711 ( .a(n_43392), .b(FE_OCPN1247_n_43120), .o(n_43467) );
na02f80 g780718 ( .a(n_618), .b(n_496), .o(n_628) );
no02f80 g755570 ( .a(n_24561), .b(n_23941), .o(n_24617) );
in01f80 FE_OCP_RBC1151_n_13460 ( .a(n_13460), .o(FE_OCP_RBN1151_n_13460) );
in01f80 newInst_3542 ( .a(newNet_447), .o(newNet_3542) );
in01f80 FE_OCP_RBC1177_n_18981 ( .a(FE_OCP_RBN1176_n_18981), .o(FE_OCP_RBN1177_n_18981) );
in01f80 newInst_1062 ( .a(newNet_1061), .o(newNet_1062) );
in01f80 g765019 ( .a(n_15498), .o(n_15674) );
na02f80 g742007 ( .a(n_44031), .b(n_47252), .o(n_38164) );
in01f80 newInst_3671 ( .a(newNet_3670), .o(newNet_3671) );
na02f80 g780101 ( .a(n_1119), .b(n_1096), .o(n_1097) );
in01f80 g745179 ( .a(n_34540), .o(n_34541) );
in01f80 newInst_2706 ( .a(newNet_540), .o(newNet_2706) );
na02f80 g760745 ( .a(n_19622), .b(n_19617), .o(n_19690) );
in01f80 g750257 ( .a(n_30895), .o(n_30896) );
no02f80 g748564 ( .a(n_31588), .b(n_31547), .o(n_31720) );
in01f80 FE_OCP_DRV_C3159_n_31303 ( .a(n_31303), .o(FE_OCP_DRV_N3159_n_31303) );
in01f80 newInst_1188 ( .a(newNet_1187), .o(newNet_1188) );
in01f80 newInst_284 ( .a(newNet_14), .o(newNet_284) );
in01f80 g739097 ( .a(n_41444), .o(n_41050) );
in01f80 g744202 ( .a(n_36291), .o(n_36292) );
in01f80 g747826 ( .a(n_33461), .o(n_33513) );
na02f80 g738562 ( .a(n_41567), .b(n_41568), .o(n_41665) );
na02f80 g737591 ( .a(n_42766), .b(n_42725), .o(n_42788) );
na02f80 g774043 ( .a(n_6804), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .o(n_6842) );
no02f80 g777762 ( .a(n_3318), .b(n_2485), .o(n_3298) );
no02f80 g765579 ( .a(n_15396), .b(n_14045), .o(n_15447) );
na02f80 g761824 ( .a(n_19125), .b(n_18731), .o(n_19197) );
in01f80 newInst_3212 ( .a(newNet_3211), .o(newNet_3212) );
na02f80 g769303 ( .a(n_11475), .b(n_10544), .o(n_11510) );
no02f80 g745096 ( .a(n_34714), .b(n_34687), .o(n_34688) );
in01f80 g770204 ( .a(n_10711), .o(n_10770) );
in01f80 newInst_2274 ( .a(newNet_2273), .o(newNet_2274) );
in01f80 g768258 ( .a(n_12599), .o(n_12600) );
no02f80 g748657 ( .a(n_31269), .b(n_31300), .o(n_31330) );
na02f80 g740684 ( .a(n_39567), .b(n_39453), .o(n_39601) );
in01f80 g771352 ( .a(n_9353), .o(n_9372) );
oa22f80 FE_RC_1398_0 ( .a(n_35971), .b(n_36447), .c(n_45617), .d(n_35972), .o(n_36520) );
no02f80 FE_RC_4015_0 ( .a(FE_RN_1314_0), .b(n_15316), .o(FE_RN_1743_0) );
na02f80 g771064 ( .a(FE_OCP_RBN2750_n_9629), .b(FE_OCP_RBN2619_n_44561), .o(n_9717) );
in01f80 g765149 ( .a(n_15380), .o(n_15381) );
no02f80 g767468 ( .a(n_13444), .b(n_13443), .o(n_13445) );
no02f80 g746813 ( .a(n_32961), .b(n_32897), .o(n_33485) );
in01f80 g774740 ( .a(n_6408), .o(n_6409) );
in01f80 g760644 ( .a(n_19754), .o(n_19778) );
in01f80 g770001 ( .a(n_10991), .o(n_11012) );
na02f80 g748572 ( .a(n_32658), .b(n_32447), .o(n_32676) );
no02f80 g776966 ( .a(n_5356), .b(n_6250), .o(n_5439) );
in01f80 g761891 ( .a(n_18481), .o(n_18432) );
na02f80 g769179 ( .a(n_11797), .b(n_11710), .o(n_12071) );
in01f80 FE_OCP_RBC3441_n_37945 ( .a(n_37945), .o(FE_OCP_RBN3441_n_37945) );
ao12f80 FE_RC_2955_0 ( .a(FE_RN_1289_0), .b(FE_RN_1290_0), .c(n_10944), .o(n_11118) );
in01f80 FE_OCP_RBC2427_n_19599 ( .a(n_19599), .o(FE_OCP_RBN2427_n_19599) );
in01f80 fopt784724 ( .a(n_22682), .o(n_47207) );
no02f80 g780929 ( .a(n_457), .b(n_479), .o(n_463) );
na02f80 g751978 ( .a(n_28793), .b(n_28937), .o(n_28988) );
in01f80 g749534 ( .a(n_31871), .o(n_30554) );
ao12f80 g784674 ( .a(n_5012), .b(n_4933), .c(n_4348), .o(n_47004) );
in01f80 g775829 ( .a(n_5198), .o(n_5199) );
in01f80 FE_OCP_RBC2788_n_4294 ( .a(n_4294), .o(FE_OCP_RBN2788_n_4294) );
no02f80 g778731 ( .a(FE_OCPN871_n_2737), .b(n_2738), .o(n_2838) );
na02f80 g738717 ( .a(n_41378), .b(n_41401), .o(n_41445) );
in01f80 g736416 ( .a(n_43759), .o(n_43772) );
na02f80 g777648 ( .a(n_3469), .b(FE_OCP_RBN2486_n_3498), .o(n_3538) );
in01f80 g780447 ( .a(n_935), .o(n_782) );
no02f80 g755877 ( .a(n_25771), .b(n_25735), .o(n_26134) );
na02f80 g761965 ( .a(n_18225), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .o(n_18434) );
na02f80 g749456 ( .a(n_30575), .b(FE_OCPN1410_n_27014), .o(n_30621) );
na02f80 g751948 ( .a(n_28757), .b(n_28756), .o(n_28758) );
in01f80 newInst_1815 ( .a(newNet_1814), .o(newNet_1815) );
in01f80 g780842 ( .a(n_571), .o(n_572) );
in01f80 g765944 ( .a(n_14772), .o(n_14792) );
no02f80 g747798 ( .a(n_33315), .b(n_32900), .o(n_33393) );
oa12f80 g736318 ( .a(n_339), .b(n_43845), .c(n_43918), .o(n_43886) );
in01f80 newInst_3218 ( .a(newNet_2208), .o(newNet_3218) );
in01f80 newInst_718 ( .a(newNet_717), .o(newNet_718) );
ao12f80 g770350 ( .a(n_10638), .b(n_10659), .c(n_10637), .o(n_10716) );
in01f80 g770262 ( .a(n_10784), .o(n_10785) );
na02f80 g736774 ( .a(n_43043), .b(n_43024), .o(n_43055) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_15_ ( .ck(newNet_967), .d(n_22960), .o(delay_xor_ln21_unr15_stage6_stallmux_q_15_) );
oa12f80 g736603 ( .a(n_43159), .b(n_43157), .c(n_43038), .o(n_43335) );
in01f80 g749383 ( .a(n_30608), .o(n_30626) );
na02f80 g774899 ( .a(n_6168), .b(n_6190), .o(n_6297) );
oa12f80 g755824 ( .a(n_25368), .b(n_25160), .c(n_25304), .o(n_26237) );
no02f80 g748574 ( .a(FE_OCP_RBN1211_n_31515), .b(n_27536), .o(n_31589) );
no02f80 g742149 ( .a(FE_OCP_RBN2256_n_37844), .b(n_37617), .o(n_38036) );
in01f80 g754853 ( .a(n_25650), .o(n_25651) );
in01f80 g776934 ( .a(n_3724), .o(n_3744) );
oa12f80 g775995 ( .a(n_4688), .b(n_4624), .c(n_4601), .o(n_4815) );
na02f80 g743420 ( .a(n_36646), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36717) );
no02f80 g770146 ( .a(n_10871), .b(n_10805), .o(n_10872) );
no02f80 g760402 ( .a(n_20095), .b(n_18605), .o(n_20170) );
no03m80 FE_RC_1128_0 ( .a(n_40688), .b(n_40781), .c(n_40734), .o(n_40798) );
na02f80 g761669 ( .a(n_18649), .b(n_18681), .o(n_18754) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_28_ ( .ck(newNet_3126), .d(n_40585), .o(delay_add_ln22_unr27_stage10_stallmux_q_28_) );
no02f80 g762267 ( .a(FE_OFN750_n_45003), .b(n_18660), .o(n_18818) );
no02f80 g748976 ( .a(n_31023), .b(FE_OCPN1486_n_27315), .o(n_31108) );
in01f80 newInst_3449 ( .a(newNet_3448), .o(newNet_3449) );
oa22f80 FE_RC_37_0 ( .a(FE_OFN84_n_46137), .b(n_6725), .c(FE_OFN806_n_46196), .d(n_6774), .o(n_46193) );
oa12f80 g780218 ( .a(n_749), .b(n_1056), .c(n_845), .o(n_1093) );
in01f80 newInst_2671 ( .a(newNet_2670), .o(newNet_2671) );
oa12f80 g746153 ( .a(n_34701), .b(n_35045), .c(n_34639), .o(n_35109) );
in01f80 g748667 ( .a(n_31437), .o(n_31438) );
in01f80 FE_OCP_RBC3565_n_29857 ( .a(FE_OCP_RBN3561_n_29857), .o(FE_OCP_RBN3565_n_29857) );
na02f80 g736531 ( .a(n_43686), .b(n_43217), .o(n_43687) );
in01f80 FE_RC_580_0 ( .a(n_23390), .o(FE_RN_177_0) );
na02f80 g778393 ( .a(n_2446), .b(n_2445), .o(n_2447) );
in01f80 FE_OCP_RBC3481_n_13667 ( .a(n_13667), .o(FE_OCP_RBN3481_n_13667) );
in01f80 g765517 ( .a(n_15667), .o(n_15668) );
in01f80 g738394 ( .a(n_41705), .o(n_41706) );
no02f80 g779629 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .o(n_2030) );
in01f80 g763455 ( .a(n_17313), .o(n_17314) );
na02f80 g757832 ( .a(n_22447), .b(n_22472), .o(n_22553) );
in01f80 newInst_848 ( .a(newNet_510), .o(newNet_848) );
na02f80 g780405 ( .a(n_881), .b(n_778), .o(n_800) );
no02f80 FE_RC_1306_0 ( .a(FE_RN_383_0), .b(n_20404), .o(n_20654) );
in01f80 FE_OCPC914_n_7832 ( .a(n_7832), .o(FE_OCPN914_n_7832) );
in01f80 FE_OCP_RBC3630_n_25656 ( .a(n_25656), .o(FE_OCP_RBN3630_n_25656) );
na02f80 g779094 ( .a(n_2004), .b(delay_add_ln22_unr2_stage2_stallmux_q_13_), .o(n_2049) );
no02f80 g768125 ( .a(n_12716), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .o(n_12731) );
no02f80 g741472 ( .a(n_38781), .b(n_38780), .o(n_38782) );
in01f80 FE_OCP_RBC2951_n_21489 ( .a(n_21489), .o(FE_OCP_RBN2951_n_21489) );
in01f80 newInst_2370 ( .a(newNet_2369), .o(newNet_2370) );
no02f80 g752548 ( .a(n_28281), .b(n_27953), .o(n_28339) );
na02f80 g772837 ( .a(n_8023), .b(n_8011), .o(n_8342) );
na02f80 g765261 ( .a(n_15230), .b(n_15263), .o(n_15376) );
in01f80 g776496 ( .a(n_4538), .o(n_4525) );
in01f80 newInst_2057 ( .a(newNet_2056), .o(newNet_2057) );
no02f80 g777775 ( .a(n_3498), .b(n_2759), .o(n_3312) );
no02f80 g758066 ( .a(n_23295), .b(n_22730), .o(n_23296) );
na02f80 g737385 ( .a(n_42810), .b(n_42795), .o(n_43104) );
in01f80 newInst_1093 ( .a(newNet_1092), .o(newNet_1093) );
na02f80 g757201 ( .a(n_23225), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .o(n_23289) );
oa12f80 g769385 ( .a(FE_OCP_RBN2105_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_11542), .c(n_9777), .o(n_11543) );
in01f80 g737340 ( .a(n_42843), .o(n_42889) );
na02f80 g778733 ( .a(n_2235), .b(n_2234), .o(n_2261) );
in01f80 g777682 ( .a(n_47019), .o(n_3439) );
in01f80 g744976 ( .a(n_46953), .o(n_36402) );
in01f80 g765841 ( .a(n_14908), .o(n_14925) );
na02f80 g737308 ( .a(n_42873), .b(n_42859), .o(n_42910) );
ao12f80 g761366 ( .a(n_19828), .b(n_20086), .c(n_19760), .o(n_20328) );
in01f80 FE_OCP_DRV_C1551_n_19010 ( .a(n_19010), .o(FE_OCP_DRV_N1551_n_19010) );
oa22f80 g758202 ( .a(n_22657), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(FE_OCP_RBN2046_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .d(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n_23157) );
in01f80 g778166 ( .a(n_2872), .o(n_2873) );
no02f80 g749911 ( .a(n_29899), .b(n_29898), .o(n_29900) );
no03m80 FE_RC_3186_0 ( .a(FE_RN_1414_0), .b(FE_OCP_RBN3372_n_6745), .c(n_6523), .o(n_6802) );
in01f80 FE_OCP_RBC3549_n_44575 ( .a(FE_OCP_RBN3543_n_44575), .o(FE_OCP_RBN3549_n_44575) );
no02f80 g771441 ( .a(n_9521), .b(n_9398), .o(n_9562) );
no02f80 g784100 ( .a(n_7156), .b(delay_add_ln22_unr5_stage3_stallmux_q_14_), .o(n_45843) );
na02f80 g757290 ( .a(n_23187), .b(n_23125), .o(n_23204) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_21_ ( .ck(newNet_2472), .d(n_32384), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_) );
na02f80 g737661 ( .a(n_42502), .b(n_42519), .o(n_42585) );
na02f80 g773942 ( .a(n_7217), .b(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .o(n_7255) );
no02f80 g751906 ( .a(n_28897), .b(n_29041), .o(n_29069) );
in01f80 newInst_3638 ( .a(newNet_1712), .o(newNet_3638) );
in01f80 FE_OCP_RBC1356_n_44259 ( .a(n_44259), .o(FE_OCP_RBN1356_n_44259) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_4_ ( .ck(newNet_3483), .d(n_21341), .o(delay_add_ln22_unr14_stage6_stallmux_q_4_) );
ao22s80 g778905 ( .a(FE_OCP_RBN2287_n_2268), .b(n_2001), .c(n_2268), .d(n_2002), .o(n_2380) );
in01f80 g759241 ( .a(n_21266), .o(n_21306) );
no02f80 g769630 ( .a(n_11183), .b(FE_OCP_RBN3038_n_47269), .o(n_11251) );
in01f80 g762415 ( .a(n_18443), .o(n_18534) );
na02f80 g738981 ( .a(n_41207), .b(n_40934), .o(n_41246) );
no02f80 g775640 ( .a(n_5570), .b(n_5591), .o(n_5746) );
na02f80 g775759 ( .a(n_5452), .b(n_4908), .o(n_5468) );
oa12f80 g736274 ( .a(n_296), .b(n_43887), .c(FE_OFN4_n_43918), .o(n_43910) );
no02f80 g753596 ( .a(n_26654), .b(n_26584), .o(n_26696) );
in01f80 g775318 ( .a(n_5974), .o(n_5975) );
ao12f80 g779432 ( .a(n_2108), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .o(n_2116) );
in01f80 g769808 ( .a(n_11194), .o(n_11218) );
in01f80 g775408 ( .a(n_5751), .o(n_5752) );
in01f80 newInst_936 ( .a(newNet_935), .o(newNet_936) );
in01f80 g775039 ( .a(FE_OCP_RBN3048_n_6013), .o(n_6028) );
na02f80 g736788 ( .a(n_43389), .b(n_43520), .o(n_43558) );
oa12f80 g775642 ( .a(n_5482), .b(n_5510), .c(n_5481), .o(n_5618) );
ao22s80 FE_RC_1296_0 ( .a(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_24366), .c(n_22089), .d(n_24395), .o(n_24465) );
in01f80 newInst_2928 ( .a(newNet_1360), .o(newNet_2928) );
in01f80 FE_OCP_RBC2379_n_3502 ( .a(n_3502), .o(FE_OCP_RBN2379_n_3502) );
na02f80 g771271 ( .a(n_9342), .b(n_8309), .o(n_9424) );
in01f80 newInst_2387 ( .a(newNet_298), .o(newNet_2387) );
in01f80 g747095 ( .a(n_32800), .o(n_32801) );
in01f80 newInst_289 ( .a(newNet_192), .o(newNet_289) );
in01f80 g775699 ( .a(n_5499), .o(n_5500) );
no02f80 g756167 ( .a(n_24864), .b(n_24845), .o(n_24846) );
no02f80 g759419 ( .a(n_20886), .b(n_20885), .o(n_20956) );
na02f80 g756850 ( .a(n_23363), .b(delay_add_ln22_unr14_stage6_stallmux_q_10_), .o(n_23369) );
in01f80 g774862 ( .a(n_6222), .o(n_6223) );
no02f80 g767252 ( .a(n_13606), .b(n_13551), .o(n_13607) );
no02f80 g767764 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .o(n_13356) );
no02f80 g745855 ( .a(n_35391), .b(n_35335), .o(n_35392) );
in01f80 newInst_2038 ( .a(newNet_2037), .o(newNet_2038) );
na02f80 g751610 ( .a(n_29252), .b(n_29105), .o(n_29177) );
in01f80 FE_OCP_RBC3083_n_31819 ( .a(n_31819), .o(FE_OCP_RBN3083_n_31819) );
in01f80 newInst_52 ( .a(newNet_51), .o(newNet_52) );
in01f80 newInst_1417 ( .a(newNet_119), .o(newNet_1417) );
in01f80 g753932 ( .a(n_26263), .o(n_26264) );
no02f80 g740824 ( .a(n_39440), .b(n_38981), .o(n_39406) );
na02f80 g740191 ( .a(FE_OCP_RBN3718_n_39913), .b(n_39586), .o(n_40188) );
na02f80 g777005 ( .a(n_4063), .b(n_4036), .o(n_4140) );
oa12f80 g754942 ( .a(FE_OCP_RBN3586_n_25295), .b(n_25201), .c(n_25294), .o(n_25453) );
no02f80 g756866 ( .a(n_23811), .b(n_23704), .o(n_23705) );
no02f80 g763487 ( .a(FE_OCP_RBN3081_n_16977), .b(n_15549), .o(n_17118) );
in01f80 g765242 ( .a(n_15453), .o(n_15454) );
in01f80 g765735 ( .a(n_15514), .o(n_15599) );
no02f80 g756381 ( .a(n_24016), .b(n_23857), .o(n_24498) );
na02f80 g753813 ( .a(n_26373), .b(FE_OCPN1508_n_23414), .o(n_26409) );
in01f80 g763316 ( .a(n_16917), .o(n_16918) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_20_ ( .ck(newNet_3144), .d(n_40487), .o(delay_add_ln22_unr27_stage10_stallmux_q_20_) );
in01f80 FE_RC_1241_0 ( .a(FE_RN_374_0), .o(n_8981) );
oa12f80 g741484 ( .a(n_38740), .b(n_38774), .c(n_38754), .o(n_38807) );
in01f80 g779510 ( .a(n_1983), .o(n_1984) );
in01f80 g755931 ( .a(n_24429), .o(n_24457) );
in01f80 newInst_1873 ( .a(newNet_829), .o(newNet_1873) );
no03m80 g751290 ( .a(n_29078), .b(n_29721), .c(n_29306), .o(n_29758) );
in01f80 g778619 ( .a(n_2295), .o(n_2296) );
oa22f80 FE_RC_2594_0 ( .a(n_1401), .b(n_1491), .c(n_1494), .d(n_1492), .o(n_1585) );
no02f80 g767525 ( .a(n_13183), .b(n_13290), .o(n_13184) );
in01f80 g764771 ( .a(n_15765), .o(n_15797) );
na02f80 g754924 ( .a(n_25542), .b(n_24546), .o(n_25543) );
no02f80 g777660 ( .a(n_3495), .b(n_3494), .o(n_3539) );
ao12f80 g765582 ( .a(n_14426), .b(n_15481), .c(n_14388), .o(n_15573) );
no02f80 g740861 ( .a(n_39342), .b(n_39046), .o(n_39379) );
no02f80 g763470 ( .a(n_16987), .b(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n_17125) );
no02f80 g761689 ( .a(n_18602), .b(FE_OCPN1776_n_18263), .o(n_18601) );
no02f80 g762829 ( .a(FE_OCP_RBN2140_FE_OCPN861_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .o(n_17845) );
no02f80 g767959 ( .a(n_13104), .b(n_13200), .o(n_13201) );
ao12f80 g757075 ( .a(n_23567), .b(n_23566), .c(n_23565), .o(n_23806) );
oa12f80 g763961 ( .a(n_16564), .b(n_16565), .c(n_16535), .o(n_16607) );
in01f80 g776672 ( .a(n_4050), .o(n_4051) );
na02f80 g740980 ( .a(n_39059), .b(n_38984), .o(n_39313) );
oa22f80 g784540 ( .a(n_11778), .b(FE_OFN802_n_46285), .c(n_11725), .d(FE_OCP_RBN3043_n_46337), .o(n_46361) );
no02f80 g745064 ( .a(n_34858), .b(n_34857), .o(n_34859) );
in01f80 newInst_2837 ( .a(newNet_1627), .o(newNet_2837) );
no02f80 g746766 ( .a(n_33062), .b(n_33015), .o(n_33143) );
oa22f80 g779885 ( .a(n_44652), .b(n_1164), .c(n_44637), .d(n_1157), .o(n_1298) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_5_ ( .ck(newNet_2810), .d(n_10222), .o(delay_add_ln22_unr8_stage4_stallmux_q_5_) );
oa22f80 g757785 ( .a(n_22425), .b(n_22801), .c(n_22390), .d(n_22580), .o(n_22480) );
na02f80 g753522 ( .a(n_27449), .b(n_26770), .o(n_27540) );
ao12f80 g751423 ( .a(n_28460), .b(n_28533), .c(n_28523), .o(n_28534) );
in01f80 g761508 ( .a(n_19820), .o(n_19821) );
in01f80 FE_OCP_DRV_C3151_n_13264 ( .a(n_13264), .o(FE_OCP_DRV_N3151_n_13264) );
no02f80 g763815 ( .a(n_17498), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .o(n_17574) );
ao12f80 g747164 ( .a(n_32759), .b(n_32758), .c(FE_OCP_RBN1339_n_32653), .o(n_33958) );
in01f80 FE_OCP_RBC2431_n_14018 ( .a(FE_OCP_RBN2430_n_14018), .o(FE_OCP_RBN2431_n_14018) );
na02f80 g739881 ( .a(n_40478), .b(n_40480), .o(n_40737) );
in01f80 newInst_978 ( .a(newNet_651), .o(newNet_978) );
na02f80 g748508 ( .a(n_31518), .b(n_30989), .o(n_31702) );
na02f80 g753579 ( .a(n_26662), .b(n_26316), .o(n_26726) );
in01f80 FE_OCP_RBC3440_n_33803 ( .a(n_33803), .o(FE_OCP_RBN3440_n_33803) );
ao12f80 g765634 ( .a(n_15399), .b(n_15446), .c(n_15398), .o(n_15870) );
in01f80 g736361 ( .a(n_43811), .o(n_43812) );
in01f80 g759514 ( .a(n_20883), .o(n_20884) );
no02f80 g759424 ( .a(n_21059), .b(FE_OCPUNCON3146_n_21058), .o(n_21174) );
ao22s80 FE_RC_2660_0 ( .a(n_27970), .b(n_27935), .c(n_27934), .d(FE_OCP_RBN3371_n_27970), .o(n_28085) );
ao12f80 g756504 ( .a(n_23735), .b(n_23678), .c(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n_23786) );
in01f80 FE_OFC771_n_46337 ( .a(FE_OCP_RBN3040_n_46337), .o(FE_OFN771_n_46337) );
in01f80 g745460 ( .a(n_34433), .o(n_34434) );
oa22f80 g746642 ( .a(n_33204), .b(n_33011), .c(n_33162), .d(n_33010), .o(n_34051) );
no02f80 g758133 ( .a(n_22411), .b(n_22554), .o(n_22502) );
no02f80 g751965 ( .a(n_28836), .b(n_28837), .o(n_28864) );
no02f80 g736700 ( .a(n_43225), .b(n_43188), .o(n_43329) );
in01f80 FE_OCP_RBC2296_n_2438 ( .a(FE_OCP_RBN2292_n_2438), .o(FE_OCP_RBN2296_n_2438) );
na02f80 g753909 ( .a(n_26189), .b(FE_RN_1643_0), .o(n_26292) );
no02f80 g743519 ( .a(n_36608), .b(n_36750), .o(n_36609) );
na02f80 g762915 ( .a(n_17683), .b(n_17592), .o(n_17624) );
ao22s80 FE_RC_3883_0 ( .a(n_20749), .b(n_21093), .c(n_20751), .d(n_21143), .o(n_21194) );
no02f80 g738676 ( .a(n_41525), .b(n_41339), .o(n_41724) );
oa12f80 g772453 ( .a(n_45213), .b(n_8387), .c(n_7464), .o(n_8476) );
no02f80 g765839 ( .a(n_14877), .b(n_14878), .o(n_14953) );
in01f80 g777136 ( .a(n_3780), .o(n_3781) );
na02f80 g754889 ( .a(n_25385), .b(n_25421), .o(n_25507) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_14_ ( .ck(newNet_3553), .d(n_22275), .o(delay_add_ln22_unr14_stage6_stallmux_q_14_) );
oa12f80 g751933 ( .a(n_28755), .b(n_28754), .c(n_28753), .o(n_29077) );
oa12f80 g736378 ( .a(n_315), .b(n_43793), .c(n_43918), .o(n_43851) );
na02f80 g771278 ( .a(n_9292), .b(FE_OCPN901_n_44593), .o(n_9302) );
na02f80 g759555 ( .a(n_20872), .b(n_19098), .o(n_20930) );
in01f80 newInst_639 ( .a(newNet_615), .o(newNet_639) );
no02f80 g759063 ( .a(n_21230), .b(n_21229), .o(n_21280) );
na02f80 g775346 ( .a(n_5860), .b(n_5859), .o(n_5861) );
in01f80 g746300 ( .a(n_35678), .o(n_34988) );
in01f80 FE_OCP_RBC3480_n_13664 ( .a(n_13664), .o(FE_OCP_RBN3480_n_13664) );
no02f80 g757698 ( .a(n_22705), .b(n_22667), .o(n_22668) );
no02f80 g739344 ( .a(n_45147), .b(delay_add_ln22_unr27_stage10_stallmux_q_15_), .o(n_40705) );
in01f80 g768646 ( .a(n_12319), .o(n_12320) );
ao12f80 g768992 ( .a(n_11885), .b(FE_OCP_RBN2119_n_45224), .c(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .o(n_12295) );
no02f80 g750021 ( .a(n_30279), .b(n_30258), .o(n_30316) );
in01f80 newInst_1669 ( .a(newNet_1668), .o(newNet_1669) );
na02f80 g778663 ( .a(FE_OCPN1234_n_2414), .b(n_2515), .o(n_2544) );
na02f80 g767775 ( .a(n_13015), .b(n_12986), .o(n_13016) );
no02f80 g742683 ( .a(n_37545), .b(n_37452), .o(n_37546) );
in01f80 g737452 ( .a(n_42671), .o(n_42672) );
na02f80 g774089 ( .a(n_6798), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .o(n_6824) );
na02f80 g762742 ( .a(n_17875), .b(FE_OCP_RBN2144_FE_OCPN861_n_45450), .o(n_17917) );
oa12f80 g770476 ( .a(n_9942), .b(n_10277), .c(n_9978), .o(n_10404) );
in01f80 g736765 ( .a(n_43353), .o(n_43354) );
no02f80 g777339 ( .a(n_4556), .b(FE_OFN824_n_3500), .o(n_4818) );
no02f80 g760723 ( .a(n_19567), .b(n_19641), .o(n_19642) );
no02f80 FE_RC_2377_0 ( .a(FE_RN_924_0), .b(n_12279), .o(FE_RN_925_0) );
na02f80 g776091 ( .a(n_4946), .b(n_4546), .o(n_5055) );
oa12f80 g780198 ( .a(n_1115), .b(n_1114), .c(n_1113), .o(n_1167) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_20_ ( .ck(newNet_340), .d(n_1295), .o(delay_xor_ln22_unr3_stage2_stallmux_q_20_) );
na02f80 g779255 ( .a(n_1755), .b(n_1558), .o(n_1818) );
na02f80 g778607 ( .a(n_2259), .b(n_2261), .o(n_2396) );
oa12f80 g751624 ( .a(n_28250), .b(n_28373), .c(n_28210), .o(n_28428) );
no02f80 g749150 ( .a(n_30772), .b(FE_OCPN1486_n_27315), .o(n_30890) );
no02f80 g747227 ( .a(n_33913), .b(n_33912), .o(n_33914) );
in01f80 fopt782905 ( .a(n_44352), .o(n_44351) );
na02f80 FE_RC_2268_0 ( .a(FE_RN_843_0), .b(FE_RN_841_0), .o(n_25640) );
in01f80 g766332 ( .a(n_14279), .o(n_14280) );
oa22f80 FE_RC_942_0 ( .a(n_20231), .b(n_22774), .c(n_22580), .d(n_22751), .o(n_22826) );
oa22f80 FE_RC_1679_0 ( .a(delay_sub_ln23_0_unr30_stage10_stallmux_q), .b(n_43009), .c(n_43012), .d(n_42998), .o(n_43013) );
na02f80 g747990 ( .a(n_33070), .b(n_33069), .o(n_33071) );
no02f80 g752142 ( .a(n_28060), .b(n_28114), .o(n_28164) );
na02f80 g751892 ( .a(n_28812), .b(n_28811), .o(n_28838) );
in01f80 g746370 ( .a(n_33613), .o(n_33580) );
no02f80 g763403 ( .a(n_16975), .b(n_16146), .o(n_17216) );
no02f80 g756466 ( .a(n_23758), .b(n_23823), .o(n_23848) );
na02f80 g738477 ( .a(n_41387), .b(n_41412), .o(n_41475) );
in01f80 newInst_319 ( .a(newNet_318), .o(newNet_319) );
in01f80 g774405 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .o(n_6496) );
na02f80 g741747 ( .a(n_38462), .b(n_38461), .o(n_38463) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_23_ ( .ck(newNet_1106), .d(n_11153), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_) );
oa12f80 g769739 ( .a(n_11266), .b(n_11267), .c(n_10124), .o(n_11287) );
no02f80 g742775 ( .a(n_37514), .b(n_36997), .o(n_37290) );
no02f80 g777849 ( .a(n_3135), .b(n_3026), .o(n_3193) );
in01f80 g746181 ( .a(n_33868), .o(n_33918) );
no02f80 g773061 ( .a(n_7636), .b(n_7628), .o(n_7629) );
in01f80 FE_RC_2793_0 ( .a(FE_RN_1194_0), .o(n_14203) );
oa12f80 FE_RC_2971_0 ( .a(FE_RN_1298_0), .b(FE_RN_1297_0), .c(n_26153), .o(n_26291) );
in01f80 g740697 ( .a(n_39475), .o(n_39476) );
no02f80 g744217 ( .a(n_36030), .b(n_36059), .o(n_36186) );
na02f80 g780708 ( .a(n_634), .b(n_582), .o(n_638) );
in01f80 g750443 ( .a(n_29663), .o(n_29640) );
in01f80 g736963 ( .a(n_43316), .o(n_43305) );
no02f80 g740723 ( .a(n_39408), .b(n_39455), .o(n_39494) );
na02f80 g779490 ( .a(n_1376), .b(n_1455), .o(n_1472) );
in01f80 fopt783437 ( .a(n_45032), .o(n_45024) );
na02f80 FE_RC_3860_0 ( .a(n_31246), .b(FE_RN_1685_0), .o(FE_RN_1686_0) );
ao22s80 FE_RC_1271_0 ( .a(n_9764), .b(n_44819), .c(n_9676), .d(n_9712), .o(n_9904) );
in01f80 newInst_2136 ( .a(newNet_2135), .o(newNet_2136) );
no02f80 g766590 ( .a(n_13884), .b(n_13364), .o(n_13926) );
no02f80 g745509 ( .a(n_34357), .b(n_34318), .o(n_34412) );
in01f80 FE_OCP_RBC1217_n_20595 ( .a(n_20595), .o(FE_OCP_RBN1217_n_20595) );
in01f80 FE_OCP_RBC2342_FE_OCPN870_n_2737 ( .a(FE_OCPN870_n_2737), .o(FE_OCP_RBN2342_FE_OCPN870_n_2737) );
no02f80 g757291 ( .a(n_23072), .b(n_23071), .o(n_23073) );
no02f80 g751197 ( .a(n_29909), .b(n_29851), .o(n_29937) );
na02f80 g762200 ( .a(n_18148), .b(n_17948), .o(n_18166) );
no02f80 g756324 ( .a(n_24514), .b(n_24513), .o(n_24515) );
in01f80 FE_OCPC3796_n_26115 ( .a(n_26115), .o(FE_OCPN3796_n_26115) );
in01f80 FE_OCP_RBC2676_n_4061 ( .a(n_4061), .o(FE_OCP_RBN2676_n_4061) );
in01f80 g745815 ( .a(n_34162), .o(n_34163) );
no02f80 g747845 ( .a(n_32188), .b(n_31970), .o(n_32238) );
in01f80 newInst_2364 ( .a(newNet_2363), .o(newNet_2364) );
in01f80 g767811 ( .a(n_13378), .o(n_13314) );
na02f80 g756060 ( .a(n_25188), .b(n_24793), .o(n_25290) );
in01f80 g739822 ( .a(n_40453), .o(n_40470) );
na02f80 g740362 ( .a(n_39761), .b(n_39760), .o(n_39762) );
na02f80 FE_RC_3296_0 ( .a(n_23040), .b(FE_RN_1450_0), .o(n_23064) );
na02f80 g747811 ( .a(n_33315), .b(n_33314), .o(n_33357) );
no02f80 g769118 ( .a(n_11583), .b(n_11405), .o(n_11702) );
na02f80 g754948 ( .a(n_25327), .b(n_24392), .o(n_25455) );
in01f80 g747197 ( .a(n_33888), .o(n_33952) );
no02f80 g744074 ( .a(n_44223), .b(n_35980), .o(n_36068) );
in01f80 g746827 ( .a(n_33182), .o(n_33183) );
na02f80 g750296 ( .a(n_29762), .b(FE_OCP_RBN2376_n_29480), .o(n_29786) );
no02f80 g778042 ( .a(n_2862), .b(n_2980), .o(n_3051) );
in01f80 g746167 ( .a(n_33731), .o(n_33732) );
oa22f80 FE_RC_960_0 ( .a(n_28336), .b(n_32394), .c(n_32566), .d(n_32463), .o(n_32511) );
na02f80 g755535 ( .a(n_24748), .b(n_24747), .o(n_24822) );
no02f80 g743980 ( .a(n_35947), .b(n_35974), .o(n_36008) );
na02f80 g774882 ( .a(n_6270), .b(n_6186), .o(n_6324) );
no02f80 FE_RC_2464_0 ( .a(FE_RN_989_0), .b(n_14217), .o(FE_RN_990_0) );
in01f80 g773287 ( .a(n_7612), .o(n_7576) );
in01f80 g755408 ( .a(n_24911), .o(n_24912) );
no02f80 g770578 ( .a(n_10465), .b(FE_OCP_RBN3560_n_8809), .o(n_10463) );
in01f80 g771615 ( .a(n_9439), .o(n_9440) );
ao12f80 g760523 ( .a(n_19837), .b(n_19817), .c(n_19775), .o(n_19950) );
na02f80 g742060 ( .a(FE_OCP_RBN2256_n_37844), .b(n_37912), .o(n_37914) );
in01f80 g754162 ( .a(n_26083), .o(n_26084) );
in01f80 g738098 ( .a(n_42103), .o(n_42104) );
in01f80 g747865 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .o(n_32275) );
in01f80 FE_OCP_RBC2313_n_41420 ( .a(n_41420), .o(FE_OCP_RBN2313_n_41420) );
oa22f80 g739729 ( .a(n_40434), .b(n_40285), .c(n_40435), .d(n_40286), .o(n_40477) );
in01f80 g756908 ( .a(n_23365), .o(n_23420) );
na02f80 g736790 ( .a(n_43519), .b(n_43087), .o(n_43556) );
na02f80 g773231 ( .a(n_7556), .b(n_7549), .o(n_7592) );
in01f80 g771288 ( .a(n_9836), .o(n_9837) );
na02f80 g772582 ( .a(n_8483), .b(n_8555), .o(n_8566) );
no02f80 g768915 ( .a(n_11845), .b(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n_11846) );
in01f80 newInst_445 ( .a(newNet_152), .o(newNet_445) );
oa12f80 g778157 ( .a(n_2755), .b(n_2754), .c(n_2753), .o(n_4433) );
in01f80 g775117 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .o(n_6061) );
in01f80 newInst_885 ( .a(newNet_203), .o(newNet_885) );
in01f80 g747660 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .o(n_32329) );
no02f80 g741922 ( .a(n_38074), .b(n_38071), .o(n_38072) );
no02f80 g740941 ( .a(n_39212), .b(n_39157), .o(n_39236) );
in01f80 FE_RC_3163_0 ( .a(FE_OCP_RBN1134_n_16041), .o(FE_RN_1402_0) );
no02f80 g745757 ( .a(n_34278), .b(n_34003), .o(n_34306) );
na02f80 g745560 ( .a(n_47255), .b(n_34454), .o(n_34558) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_3_ ( .ck(newNet_1576), .d(n_26998), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_) );
in01f80 g780147 ( .a(n_1189), .o(n_1179) );
in01f80 g768333 ( .a(n_12618), .o(n_12975) );
na02f80 g743433 ( .a(n_36588), .b(n_36750), .o(n_36589) );
oa12f80 g738996 ( .a(n_41145), .b(n_41144), .c(n_41143), .o(n_41492) );
in01f80 g755150 ( .a(n_25743), .o(n_25744) );
na02f80 g760057 ( .a(n_20375), .b(n_20436), .o(n_20499) );
no02f80 FE_RC_4211_0 ( .a(n_14554), .b(FE_RN_1843_0), .o(FE_RN_1844_0) );
no02f80 g765532 ( .a(n_15664), .b(n_15665), .o(n_15839) );
no02f80 g775510 ( .a(n_5739), .b(n_5681), .o(n_5763) );
na02f80 g756547 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .o(n_23767) );
oa22f80 g754891 ( .a(n_25542), .b(FE_OCPN1048_n_24819), .c(n_25481), .d(n_24865), .o(n_25721) );
in01f80 newInst_593 ( .a(newNet_592), .o(newNet_593) );
no02f80 g751809 ( .a(n_29151), .b(n_29127), .o(n_29202) );
in01f80 g756207 ( .a(n_24102), .o(n_24101) );
oa12f80 g778901 ( .a(n_2178), .b(n_2177), .c(n_2176), .o(n_2644) );
in01f80 g779655 ( .a(n_1778), .o(n_1779) );
no02f80 g737510 ( .a(n_42454), .b(n_42632), .o(n_42664) );
no02f80 g748581 ( .a(n_31404), .b(FE_OCPN1520_n_31403), .o(n_31424) );
in01f80 g776100 ( .a(n_5116), .o(n_5117) );
in01f80 g748519 ( .a(n_31468), .o(n_31469) );
no02f80 g739958 ( .a(n_40024), .b(n_40047), .o(n_40048) );
in01f80 newInst_2818 ( .a(newNet_2817), .o(newNet_2818) );
no02f80 g736782 ( .a(n_43359), .b(n_43349), .o(n_43394) );
no03m80 FE_RC_3547_0 ( .a(FE_RN_1536_0), .b(n_32741), .c(n_32740), .o(FE_RN_1537_0) );
no02f80 g759680 ( .a(n_21781), .b(n_21718), .o(n_21796) );
na02f80 FE_RC_16_0 ( .a(n_2365), .b(FE_RN_5_0), .o(n_2431) );
na02f80 g752175 ( .a(n_28592), .b(n_28054), .o(n_28638) );
no02f80 g746817 ( .a(n_33211), .b(n_33252), .o(n_33265) );
in01f80 newInst_3169 ( .a(newNet_374), .o(newNet_3169) );
no02f80 g745842 ( .a(n_44104), .b(FE_OCP_RBN3458_n_33872), .o(n_34278) );
na02f80 g778765 ( .a(n_2222), .b(n_2007), .o(n_2207) );
no02f80 g774856 ( .a(n_6266), .b(n_6250), .o(n_6251) );
in01f80 FE_OCPC875_n_44672 ( .a(FE_OCPN873_n_44672), .o(FE_OCPN875_n_44672) );
in01f80 g756410 ( .a(n_24014), .o(n_24052) );
no02f80 g739054 ( .a(n_41092), .b(n_40704), .o(n_41093) );
in01f80 newInst_2320 ( .a(newNet_2319), .o(newNet_2320) );
ao12f80 g779394 ( .a(n_1538), .b(n_1537), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n_1909) );
no02f80 g753966 ( .a(n_26198), .b(n_23466), .o(n_26389) );
no02f80 g748802 ( .a(n_32390), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n_32424) );
oa22f80 g776680 ( .a(n_4190), .b(n_4097), .c(n_4191), .d(n_4096), .o(n_4438) );
no02f80 g766490 ( .a(n_13997), .b(FE_OCPN1468_n_12968), .o(n_14100) );
na02f80 g740960 ( .a(n_39135), .b(n_39272), .o(n_39305) );
no02f80 g754081 ( .a(n_26029), .b(n_25650), .o(n_26105) );
na02f80 g742095 ( .a(FE_OCP_RBN3451_n_37945), .b(n_37556), .o(n_38136) );
in01f80 FE_RC_1119_0 ( .a(n_3217), .o(FE_RN_337_0) );
in01f80 FE_OCP_RBC3617_n_20249 ( .a(FE_OCP_RBN2670_n_20249), .o(FE_OCP_RBN3617_n_20249) );
na02f80 g780390 ( .a(n_739), .b(n_717), .o(n_718) );
na02f80 g784767 ( .a(n_13489), .b(FE_OCPN860_n_12880), .o(n_47253) );
na02f80 g776732 ( .a(n_3956), .b(n_4083), .o(n_4165) );
oa12f80 g766778 ( .a(n_13743), .b(n_13827), .c(n_13800), .o(n_13828) );
in01f80 newInst_3001 ( .a(newNet_3000), .o(newNet_3001) );
no02f80 FE_RC_2695_0 ( .a(n_8021), .b(n_8776), .o(FE_RN_1129_0) );
no02f80 g751286 ( .a(n_29712), .b(n_29711), .o(n_29713) );
in01f80 g739409 ( .a(n_41022), .o(n_41023) );
in01f80 FE_OCPC1240_n_7721 ( .a(n_7721), .o(FE_OCPN1240_n_7721) );
no02f80 FE_RC_2380_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .b(FE_RN_927_0), .o(FE_RN_928_0) );
na02f80 g758682 ( .a(n_21911), .b(n_21947), .o(n_21962) );
no02f80 g755355 ( .a(n_24839), .b(n_24838), .o(n_24887) );
na02f80 g753235 ( .a(n_27377), .b(n_26201), .o(n_27381) );
ao12f80 g748695 ( .a(n_32559), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n_33130) );
ao12f80 g779500 ( .a(n_1930), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .o(n_2164) );
in01f80 g768424 ( .a(n_12447), .o(n_12448) );
in01f80 newInst_21 ( .a(newNet_20), .o(newNet_21) );
no02f80 g773214 ( .a(n_7886), .b(n_7885), .o(n_8038) );
in01f80 newInst_2564 ( .a(newNet_2563), .o(newNet_2564) );
in01f80 g760582 ( .a(n_19919), .o(n_19936) );
na02f80 g737534 ( .a(n_42291), .b(n_42318), .o(n_43021) );
no02f80 g763298 ( .a(n_17042), .b(n_16957), .o(n_17140) );
in01f80 newInst_3158 ( .a(newNet_3157), .o(newNet_3158) );
na02f80 g762071 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_26_), .o(n_18390) );
no02f80 g772429 ( .a(n_8639), .b(n_8638), .o(n_8640) );
no02f80 g743989 ( .a(n_36297), .b(n_35755), .o(n_36367) );
ao12f80 g784149 ( .a(n_38372), .b(n_38371), .c(n_45894), .o(n_45899) );
na02f80 g770803 ( .a(n_10255), .b(n_10237), .o(n_10238) );
no02f80 g741274 ( .a(n_38529), .b(FE_OCP_RBN2547_n_44944), .o(n_38981) );
ao12f80 g768603 ( .a(n_12319), .b(n_45659), .c(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .o(n_12363) );
no02f80 g759075 ( .a(n_21978), .b(n_21407), .o(n_22053) );
na02f80 FE_RC_2085_0 ( .a(FE_RN_713_0), .b(n_30727), .o(FE_RN_714_0) );
in01f80 newInst_385 ( .a(newNet_384), .o(newNet_385) );
in01f80 newInst_1625 ( .a(newNet_1624), .o(newNet_1625) );
no02f80 g775822 ( .a(n_5395), .b(n_5142), .o(n_5407) );
no02f80 g765940 ( .a(n_14774), .b(FE_OCP_RBN2272_n_13489), .o(n_14794) );
in01f80 g759004 ( .a(n_21604), .o(n_21634) );
oa12f80 g739078 ( .a(n_41022), .b(n_41083), .c(n_41052), .o(n_41112) );
in01f80 newInst_1393 ( .a(newNet_210), .o(newNet_1393) );
no02f80 g771815 ( .a(n_8932), .b(n_8931), .o(n_8933) );
no02f80 g740170 ( .a(n_39812), .b(n_46948), .o(n_40118) );
na02f80 g772685 ( .a(n_8237), .b(n_8269), .o(n_8270) );
na02f80 g746016 ( .a(n_33980), .b(n_33960), .o(n_34059) );
na02f80 g761873 ( .a(n_47247), .b(n_18345), .o(n_18370) );
in01f80 g739871 ( .a(n_40381), .o(n_40382) );
in01f80 g781252 ( .a(n_147), .o(n_148) );
no02f80 g774850 ( .a(n_45474), .b(n_5637), .o(n_6319) );
no02f80 g750643 ( .a(n_29281), .b(n_28673), .o(n_29349) );
no02f80 g752797 ( .a(n_27901), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n_27954) );
na02f80 FE_RC_562_0 ( .a(n_31697), .b(n_31678), .o(FE_RN_171_0) );
in01f80 g775314 ( .a(n_6011), .o(n_6044) );
no02f80 FE_RC_4031_0 ( .a(n_25673), .b(n_25648), .o(FE_RN_1751_0) );
na02f80 g769832 ( .a(n_11086), .b(n_11024), .o(n_11138) );
in01f80 g750157 ( .a(n_29951), .o(n_30016) );
in01f80 g775927 ( .a(n_5412), .o(n_5475) );
in01f80 g773743 ( .a(n_7236), .o(n_7226) );
in01f80 FE_OCP_RBC2399_FE_RN_347_0 ( .a(FE_RN_347_0), .o(FE_OCP_RBN2399_FE_RN_347_0) );
no02f80 g778724 ( .a(n_2438), .b(n_1888), .o(n_2534) );
na02f80 g769256 ( .a(n_11585), .b(n_10962), .o(n_11586) );
in01f80 g740954 ( .a(n_39112), .o(n_39810) );
no02f80 g761704 ( .a(n_18855), .b(FE_OCP_DRV_N1544_n_18854), .o(n_18940) );
na02f80 FE_RC_3063_0 ( .a(FE_RN_1344_0), .b(n_20694), .o(FE_RN_1345_0) );
oa12f80 g780175 ( .a(n_1117), .b(n_1116), .c(n_1148), .o(n_1168) );
in01f80 g761267 ( .a(n_19932), .o(n_19933) );
oa12f80 g765250 ( .a(n_15333), .b(n_15332), .c(n_15331), .o(n_15406) );
na02f80 g780837 ( .a(n_392), .b(n_409), .o(n_522) );
no02f80 g753664 ( .a(n_26540), .b(n_26434), .o(n_26597) );
in01f80 g775729 ( .a(n_5659), .o(n_5660) );
ao12f80 g759954 ( .a(n_20989), .b(n_20988), .c(n_20987), .o(n_21599) );
na02f80 g754732 ( .a(n_26541), .b(n_26634), .o(n_26770) );
in01f80 g745514 ( .a(n_34511), .o(n_34512) );
in01f80 FE_OCP_RBC2761_n_15200 ( .a(n_15200), .o(FE_OCP_RBN2761_n_15200) );
no02f80 g765351 ( .a(n_15224), .b(n_15223), .o(n_15340) );
oa22f80 FE_RC_2406_0 ( .a(FE_OCP_RBN1057_n_18267), .b(n_18128), .c(FE_OCP_RBN1058_n_18267), .d(n_18129), .o(n_18405) );
no02f80 g750301 ( .a(n_29778), .b(FE_OCP_DRV_N1570_n_29777), .o(n_29784) );
oa12f80 g756335 ( .a(n_24481), .b(n_24480), .c(n_24479), .o(n_25027) );
in01f80 FE_OCP_RBC3092_n_11475 ( .a(n_11475), .o(FE_OCP_RBN3092_n_11475) );
ao12f80 g779236 ( .a(FE_OCPN3755_n_1451), .b(n_1806), .c(n_1591), .o(n_1863) );
in01f80 g758711 ( .a(n_21742), .o(n_21743) );
oa22f80 FE_RC_4188_0 ( .a(FE_RN_1832_0), .b(FE_RN_1830_0), .c(FE_RN_1833_0), .d(n_24306), .o(n_24336) );
in01f80 FE_OCP_RBC1684_n_33491 ( .a(FE_OCP_RBN1682_n_33491), .o(FE_OCP_RBN1684_n_33491) );
in01f80 newInst_3315 ( .a(newNet_3314), .o(newNet_3315) );
no02f80 g741193 ( .a(FE_OCP_RBN3625_n_38870), .b(n_39393), .o(n_39421) );
in01f80 g760913 ( .a(n_19428), .o(n_19429) );
in01f80 g750086 ( .a(n_29956), .o(n_29957) );
in01f80 newInst_1939 ( .a(newNet_1938), .o(newNet_1939) );
no02f80 g749956 ( .a(n_29986), .b(n_29893), .o(n_30014) );
no02f80 g757745 ( .a(n_23158), .b(n_23157), .o(n_23159) );
in01f80 g753869 ( .a(n_26332), .o(n_26333) );
in01f80 g742455 ( .a(n_37697), .o(n_37692) );
na02f80 g740009 ( .a(n_40136), .b(n_40063), .o(n_40255) );
na02f80 g761269 ( .a(n_19679), .b(n_19845), .o(n_19991) );
no02f80 g777804 ( .a(n_3222), .b(n_2503), .o(n_3223) );
in01f80 FE_OCP_RBC3678_n_21051 ( .a(FE_OCP_RBN3677_n_21051), .o(FE_OCP_RBN3678_n_21051) );
no02f80 g753115 ( .a(n_27152), .b(n_27151), .o(n_27153) );
in01f80 g740969 ( .a(n_39212), .o(n_39254) );
in01f80 g753298 ( .a(n_27168), .o(n_27208) );
na02f80 g779558 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .o(n_2113) );
na02f80 g744464 ( .a(n_35449), .b(n_35460), .o(n_35450) );
in01f80 newInst_353 ( .a(newNet_352), .o(newNet_353) );
oa22f80 g765411 ( .a(n_15874), .b(n_16244), .c(n_16245), .d(n_16138), .o(n_16358) );
no02f80 g752209 ( .a(n_28058), .b(n_28004), .o(n_28083) );
ao12f80 g738255 ( .a(n_41892), .b(n_41891), .c(n_41890), .o(n_42312) );
ao22s80 g777713 ( .a(n_3405), .b(n_3301), .c(n_3373), .d(n_4022), .o(n_3495) );
in01f80 g738662 ( .a(n_41425), .o(n_41420) );
in01f80 newInst_1087 ( .a(newNet_211), .o(newNet_1087) );
no02f80 g765131 ( .a(n_15204), .b(n_14215), .o(n_15239) );
no02f80 g756731 ( .a(n_23464), .b(n_23478), .o(n_23555) );
in01f80 FE_RC_2210_0 ( .a(n_20914), .o(FE_RN_796_0) );
in01f80 g753305 ( .a(n_27206), .o(n_27250) );
in01f80 FE_RC_3425_0 ( .a(FE_RN_1481_0), .o(FE_RN_1482_0) );
na02f80 g769048 ( .a(n_11561), .b(n_45224), .o(n_11762) );
in01f80 newInst_2988 ( .a(newNet_2987), .o(newNet_2988) );
na02f80 g752585 ( .a(n_27593), .b(n_27353), .o(n_27608) );
oa22f80 FE_RC_3357_0 ( .a(n_27521), .b(n_27670), .c(n_27522), .d(n_27690), .o(n_27782) );
na02f80 g772886 ( .a(n_8004), .b(n_8003), .o(n_8005) );
in01f80 FE_RC_2827_0 ( .a(n_29603), .o(FE_RN_1214_0) );
na02f80 g744835 ( .a(n_35003), .b(n_30633), .o(n_35037) );
in01f80 g758194 ( .a(n_22496), .o(n_22497) );
in01f80 FE_RC_563_0 ( .a(n_31648), .o(FE_RN_172_0) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_16_ ( .ck(newNet_1021), .d(n_17808), .o(delay_xor_ln21_unr12_stage5_stallmux_q_16_) );
na02f80 g752574 ( .a(n_27585), .b(n_27597), .o(n_27653) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_28_ ( .ck(newNet_1206), .d(n_6323), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_) );
in01f80 g774529 ( .a(n_6528), .o(n_6582) );
na02f80 g766089 ( .a(n_14580), .b(n_14602), .o(n_14684) );
no02f80 FE_RC_2860_0 ( .a(n_10377), .b(FE_RN_1232_0), .o(n_10624) );
na02f80 FE_RC_2395_0 ( .a(FE_RN_940_0), .b(n_42522), .o(FE_RN_941_0) );
na02f80 g781226 ( .a(n_80), .b(beta_31), .o(n_130) );
ao12f80 g747313 ( .a(n_33864), .b(n_33863), .c(n_33862), .o(n_34474) );
no02f80 g758939 ( .a(n_21605), .b(n_21634), .o(n_21726) );
oa12f80 g736424 ( .a(n_303), .b(n_43749), .c(FE_OFN2_n_43918), .o(n_43797) );
no03m80 FE_RC_256_0 ( .a(n_20077), .b(n_20093), .c(n_20048), .o(n_20097) );
in01f80 g751879 ( .a(n_28926), .o(n_28927) );
in01f80 g775599 ( .a(n_5695), .o(n_5696) );
na02f80 g741958 ( .a(n_38138), .b(n_37996), .o(n_38185) );
oa22f80 FE_RC_3023_0 ( .a(n_40279), .b(n_40519), .c(n_40280), .d(n_40520), .o(n_40554) );
no02f80 FE_RC_1923_0 ( .a(FE_RN_607_0), .b(n_29192), .o(n_29233) );
in01f80 FE_RC_1323_0 ( .a(n_10071), .o(FE_RN_391_0) );
na02f80 g742420 ( .a(n_37738), .b(n_37737), .o(n_37765) );
in01f80 g771857 ( .a(n_10206), .o(n_10207) );
no02f80 g764656 ( .a(n_15813), .b(n_15770), .o(n_15948) );
ao22s80 g780539 ( .a(n_745), .b(n_893), .c(n_779), .d(n_748), .o(n_894) );
no02f80 g779569 ( .a(FE_OCP_RBN3249_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .o(n_1440) );
oa22f80 g740713 ( .a(n_39497), .b(n_39504), .c(n_39386), .d(n_39505), .o(n_39581) );
no02f80 g749725 ( .a(n_31409), .b(n_31408), .o(n_31431) );
no02f80 g751541 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_18_), .o(n_28494) );
ao12f80 g768614 ( .a(n_12141), .b(n_12140), .c(n_12139), .o(n_12256) );
in01f80 FE_OCPC1512_n_22280 ( .a(FE_OCPN1511_n_22280), .o(FE_OCPN1512_n_22280) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_24_ ( .ck(newNet_2549), .d(FE_OCP_RBN3133_n_27736), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_) );
in01f80 g767994 ( .a(n_12852), .o(n_12853) );
oa12f80 g751493 ( .a(n_28734), .b(n_28460), .c(n_28630), .o(n_28766) );
in01f80 g751658 ( .a(n_28419), .o(n_28438) );
in01f80 g740673 ( .a(n_39543), .o(n_39544) );
na02f80 g736710 ( .a(n_43268), .b(FE_OCPN913_n_43022), .o(n_43405) );
in01f80 g777757 ( .a(FE_OFN824_n_3500), .o(n_3501) );
na02f80 g753156 ( .a(n_27393), .b(n_27409), .o(n_27523) );
na02f80 g743243 ( .a(n_36831), .b(n_36786), .o(n_36867) );
no02f80 g754821 ( .a(n_25282), .b(n_25244), .o(n_25245) );
ao22s80 g739656 ( .a(n_40565), .b(n_40271), .c(n_40566), .d(n_40272), .o(n_40586) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_26_ ( .ck(newNet_1721), .d(n_22548), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_) );
in01f80 g758474 ( .a(n_23354), .o(n_23271) );
no02f80 g744665 ( .a(n_35212), .b(n_35185), .o(n_35293) );
in01f80 FE_RC_1797_0 ( .a(n_34037), .o(FE_RN_530_0) );
in01f80 g774221 ( .a(n_6926), .o(n_6927) );
oa22f80 FE_RC_1249_0 ( .a(n_6456), .b(n_6503), .c(n_6457), .d(n_6493), .o(n_6627) );
na02f80 g763451 ( .a(n_17119), .b(n_17169), .o(n_17317) );
in01f80 g740974 ( .a(n_39143), .o(n_39144) );
na02f80 g763225 ( .a(FE_OCP_RBN3082_n_16977), .b(n_17196), .o(n_17281) );
na02f80 g768245 ( .a(n_12675), .b(n_12674), .o(n_12676) );
na02f80 g741154 ( .a(n_38806), .b(n_38060), .o(n_38836) );
na02f80 g770063 ( .a(n_10952), .b(n_10929), .o(n_11061) );
in01f80 g755021 ( .a(n_25210), .o(n_25327) );
in01f80 FE_OCP_RBC2849_n_46982 ( .a(FE_OCP_RBN3669_n_46982), .o(FE_OCP_RBN2849_n_46982) );
ao22s80 g736396 ( .a(n_43778), .b(n_43606), .c(n_43777), .d(n_43605), .o(n_43838) );
in01f80 g758192 ( .a(n_22457), .o(n_22458) );
no02f80 g754239 ( .a(n_25940), .b(n_25565), .o(n_25966) );
in01f80 g757337 ( .a(n_23129), .o(n_23388) );
no03m80 g743658 ( .a(n_37473), .b(n_37472), .c(n_37307), .o(n_37475) );
no02f80 g758697 ( .a(n_21712), .b(n_21502), .o(n_21768) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_9_ ( .ck(newNet_2602), .d(n_21810), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_) );
in01f80 g775856 ( .a(n_5286), .o(n_5379) );
na02f80 g767929 ( .a(n_12652), .b(n_12454), .o(n_12685) );
oa12f80 g761949 ( .a(n_18109), .b(n_18267), .c(n_18071), .o(n_18318) );
in01f80 newInst_2284 ( .a(newNet_2283), .o(newNet_2284) );
no02f80 g776504 ( .a(n_4074), .b(n_2976), .o(n_4184) );
in01f80 g739678 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n_40575) );
in01f80 FE_RC_2932_0 ( .a(FE_RN_1278_0), .o(n_10810) );
in01f80 g736365 ( .a(n_43807), .o(n_43808) );
in01f80 g760393 ( .a(n_20203), .o(n_20204) );
no02f80 g766920 ( .a(n_13892), .b(n_13903), .o(n_13906) );
in01f80 g762145 ( .a(n_18774), .o(n_18775) );
na02f80 g738373 ( .a(n_41633), .b(FE_OCP_RBN2314_n_41420), .o(n_41792) );
no02f80 g770247 ( .a(n_10517), .b(n_10364), .o(n_10553) );
in01f80 g763128 ( .a(n_17863), .o(n_17862) );
in01f80 FE_RC_490_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(FE_RN_145_0) );
no02f80 g749259 ( .a(n_46958), .b(n_27130), .o(n_30821) );
in01f80 newInst_1658 ( .a(newNet_1657), .o(newNet_1658) );
in01f80 g736565 ( .a(n_43638), .o(n_43651) );
in01f80 g767268 ( .a(n_13559), .o(n_13558) );
in01f80 g752685 ( .a(n_27404), .o(n_27442) );
no02f80 g749051 ( .a(n_31019), .b(n_30990), .o(n_31126) );
in01f80 g736831 ( .a(n_43309), .o(n_43310) );
in01f80 newInst_1727 ( .a(newNet_26), .o(newNet_1727) );
na02f80 g751944 ( .a(n_28123), .b(n_28184), .o(n_28217) );
in01f80 g759731 ( .a(n_20420), .o(n_20419) );
ao12f80 g739266 ( .a(n_44797), .b(n_40882), .c(n_40558), .o(n_40941) );
no02f80 g765829 ( .a(n_14932), .b(FE_OCP_RBN2509_n_13896), .o(n_14933) );
in01f80 g771734 ( .a(n_8915), .o(n_8884) );
in01f80 g766745 ( .a(n_13849), .o(n_13850) );
in01f80 newInst_1494 ( .a(newNet_156), .o(newNet_1494) );
ms00f80 sin_out_reg_5_ ( .ck(newNet_21), .d(n_43703), .o(sin_out_5) );
na02f80 g767438 ( .a(n_13331), .b(n_13330), .o(n_13403) );
no02f80 g779013 ( .a(n_2195), .b(n_1913), .o(n_2224) );
no02f80 g754149 ( .a(n_26002), .b(FE_OCP_RBN2826_FE_RN_1573_0), .o(n_26057) );
no02f80 FE_RC_2913_0 ( .a(FE_RN_1267_0), .b(FE_RN_1265_0), .o(n_13295) );
in01f80 g770529 ( .a(n_10513), .o(n_10497) );
in01f80 newInst_2779 ( .a(newNet_2778), .o(newNet_2779) );
oa12f80 g775474 ( .a(n_5475), .b(n_5755), .c(n_5534), .o(n_5756) );
ao12f80 g747170 ( .a(n_32573), .b(n_46413), .c(n_32712), .o(n_32741) );
no02f80 g772741 ( .a(n_8179), .b(n_8165), .o(n_8235) );
in01f80 g777211 ( .a(n_3547), .o(n_3575) );
na02f80 g736489 ( .a(n_43675), .b(n_43183), .o(n_43691) );
in01f80 g736922 ( .a(n_43035), .o(n_43036) );
in01f80 FE_RC_3985_0 ( .a(FE_RN_1728_0), .o(n_14613) );
in01f80 g769150 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_19_), .o(n_11492) );
in01f80 FE_OCP_RBC3522_n_8242 ( .a(FE_OCP_RBN2407_n_8242), .o(FE_OCP_RBN3522_n_8242) );
in01f80 newInst_699 ( .a(newNet_698), .o(newNet_699) );
oa22f80 g737874 ( .a(n_42270), .b(n_41953), .c(FE_OCPN1231_n_42201), .d(n_42272), .o(n_42614) );
in01f80 newInst_3320 ( .a(newNet_3319), .o(newNet_3320) );
no02f80 g776909 ( .a(n_3762), .b(n_3029), .o(n_3919) );
in01f80 g744619 ( .a(n_35346), .o(n_35347) );
oa12f80 g780093 ( .a(n_1146), .b(n_1153), .c(n_1145), .o(n_1166) );
oa12f80 g764943 ( .a(n_15608), .b(n_15674), .c(n_15611), .o(n_15684) );
na02f80 g764958 ( .a(n_15472), .b(n_14210), .o(n_15440) );
in01f80 g754169 ( .a(n_26021), .o(n_26091) );
na02f80 g744213 ( .a(n_35857), .b(n_35814), .o(n_35971) );
oa22f80 FE_RC_1477_0 ( .a(n_17336), .b(n_17697), .c(n_16339), .d(n_17681), .o(n_17776) );
no02f80 g779100 ( .a(n_2004), .b(delay_add_ln22_unr2_stage2_stallmux_q_13_), .o(n_2017) );
no02f80 g761444 ( .a(n_20086), .b(n_19928), .o(n_20176) );
in01f80 g765174 ( .a(n_15124), .o(n_15160) );
na02f80 g740749 ( .a(n_39490), .b(n_39452), .o(n_39537) );
na02f80 g740558 ( .a(n_45531), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39668) );
no02f80 g749475 ( .a(n_30556), .b(n_30532), .o(n_30619) );
in01f80 g738102 ( .a(n_42116), .o(n_42101) );
na02f80 g747188 ( .a(n_32884), .b(n_32847), .o(n_32903) );
oa22f80 FE_RC_2951_0 ( .a(n_14722), .b(n_14665), .c(n_14693), .d(n_14723), .o(n_14823) );
na02f80 g766081 ( .a(n_14585), .b(n_13329), .o(n_14664) );
no02f80 g740059 ( .a(n_40119), .b(n_40118), .o(n_40145) );
ao12f80 g765626 ( .a(n_15443), .b(n_15481), .c(n_15442), .o(n_15961) );
oa12f80 g749626 ( .a(n_29963), .b(n_30180), .c(n_29988), .o(n_30483) );
na02f80 g776158 ( .a(n_4911), .b(n_4910), .o(n_4912) );
in01f80 FE_OCP_RBC2585_n_9009 ( .a(n_9009), .o(FE_OCP_RBN2585_n_9009) );
na02f80 g742108 ( .a(n_37970), .b(n_37968), .o(n_38082) );
no02f80 g742062 ( .a(FE_OCP_RBN2255_n_37844), .b(n_37384), .o(n_37980) );
na02f80 g759524 ( .a(n_21455), .b(n_21380), .o(n_21885) );
ao12f80 g755443 ( .a(n_25111), .b(n_25224), .c(n_25057), .o(n_25494) );
no02f80 g772014 ( .a(FE_OFN754_n_44461), .b(n_9367), .o(n_9433) );
na02f80 g737583 ( .a(n_42700), .b(n_42659), .o(n_42712) );
oa22f80 g739648 ( .a(n_40585), .b(n_40598), .c(n_40574), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40591) );
no02f80 g762835 ( .a(n_18084), .b(n_18083), .o(n_18085) );
na02f80 g764156 ( .a(n_16526), .b(n_16515), .o(n_16560) );
oa12f80 g762295 ( .a(n_18025), .b(n_18009), .c(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_18173) );
in01f80 g773154 ( .a(n_7767), .o(n_7830) );
in01f80 g748915 ( .a(n_32407), .o(n_32488) );
in01f80 g772945 ( .a(n_7843), .o(n_7894) );
in01f80 FE_OCP_RBC2884_n_26292 ( .a(n_26292), .o(FE_OCP_RBN2884_n_26292) );
na02f80 g774186 ( .a(n_6672), .b(n_6671), .o(n_6673) );
no02f80 g760146 ( .a(n_20488), .b(FE_OCP_RBN2739_n_20432), .o(n_20570) );
in01f80 FE_OCP_RBC2184_FE_RN_464_0 ( .a(FE_RN_464_0), .o(FE_OCP_RBN2184_FE_RN_464_0) );
oa12f80 g779088 ( .a(n_1982), .b(n_1987), .c(n_1981), .o(n_2766) );
na02f80 g760571 ( .a(FE_OCP_RBN2469_n_19806), .b(n_19862), .o(n_19865) );
in01f80 newInst_941 ( .a(newNet_940), .o(newNet_941) );
oa12f80 g784622 ( .a(n_38479), .b(n_38478), .c(n_38085), .o(n_46951) );
oa22f80 g767249 ( .a(n_13697), .b(n_13274), .c(n_13716), .d(n_13275), .o(n_14207) );
in01f80 fopt782893 ( .a(n_11403), .o(n_44336) );
no02f80 g751389 ( .a(n_29363), .b(n_28927), .o(n_29361) );
no02f80 g736701 ( .a(n_43285), .b(n_43185), .o(n_43286) );
in01f80 g745362 ( .a(n_35805), .o(n_35764) );
oa22f80 g784368 ( .a(FE_OFN775_n_46137), .b(n_5285), .c(FE_OFN805_n_46196), .d(n_5323), .o(n_46174) );
in01f80 newInst_1252 ( .a(newNet_156), .o(newNet_1252) );
no02f80 g756453 ( .a(n_23885), .b(n_23884), .o(n_23886) );
no02f80 g751609 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n_28867) );
oa22f80 g784359 ( .a(FE_OCP_RBN3075_FE_OFN807_n_46195), .b(n_5273), .c(FE_OFN775_n_46137), .d(n_5196), .o(n_46165) );
in01f80 g743320 ( .a(n_36737), .o(n_36738) );
no02f80 g759588 ( .a(n_20445), .b(n_20439), .o(n_20481) );
in01f80 g747575 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(n_36898) );
oa12f80 g743812 ( .a(n_37218), .b(n_37217), .c(n_46231), .o(n_37246) );
in01f80 g744968 ( .a(n_34934), .o(n_34933) );
in01f80 newInst_1012 ( .a(newNet_1011), .o(newNet_1012) );
na02f80 g761201 ( .a(n_18989), .b(n_18511), .o(n_19060) );
na02f80 g745820 ( .a(n_44101), .b(n_33604), .o(n_34184) );
in01f80 g753241 ( .a(n_27216), .o(n_27601) );
ao12f80 g779455 ( .a(n_1706), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .o(n_1992) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_27_ ( .ck(newNet_1716), .d(n_22588), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_) );
in01f80 FE_OCP_RBC2856_n_10176 ( .a(n_10176), .o(FE_OCP_RBN2856_n_10176) );
na02f80 g778032 ( .a(n_3085), .b(n_3084), .o(n_3102) );
na02f80 g760424 ( .a(n_20123), .b(n_20211), .o(n_20183) );
oa12f80 g751320 ( .a(n_29582), .b(n_29601), .c(n_29581), .o(n_30082) );
in01f80 g779475 ( .a(n_1824), .o(n_1825) );
in01f80 g773906 ( .a(n_6952), .o(n_6953) );
oa22f80 FE_RC_3916_0 ( .a(n_22492), .b(n_22573), .c(n_22593), .d(FE_OCP_RBN1730_n_22492), .o(n_22750) );
in01f80 g772707 ( .a(n_8185), .o(n_8203) );
na02f80 g767678 ( .a(n_13203), .b(n_12271), .o(n_13259) );
oa22f80 FE_RC_1466_0 ( .a(FE_OFN767_n_15670), .b(n_17685), .c(n_17753), .d(n_44147), .o(n_17754) );
in01f80 g762777 ( .a(n_18157), .o(n_18210) );
na02f80 g756477 ( .a(n_23683), .b(n_23605), .o(n_23686) );
ao12f80 g752843 ( .a(n_27990), .b(n_27762), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .o(n_28241) );
in01f80 g741638 ( .a(n_38622), .o(n_38633) );
no02f80 FE_RC_3693_0 ( .a(FE_RN_1624_0), .b(FE_RN_1246_0), .o(n_39575) );
na02f80 FE_RC_1993_0 ( .a(FE_OCP_DRV_N1556_n_19384), .b(n_19344), .o(FE_RN_651_0) );
oa12f80 g784649 ( .a(n_16559), .b(n_16527), .c(n_16486), .o(n_46979) );
ao22s80 g774238 ( .a(FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .c(n_6496), .d(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6594) );
oa12f80 g778506 ( .a(n_2352), .b(n_2369), .c(n_2351), .o(n_2558) );
in01f80 newInst_2831 ( .a(newNet_2830), .o(newNet_2831) );
in01f80 newInst_1750 ( .a(newNet_1157), .o(newNet_1750) );
in01f80 g758144 ( .a(n_22413), .o(n_22439) );
no02f80 g748004 ( .a(n_33004), .b(n_32489), .o(n_33005) );
oa12f80 g778939 ( .a(n_2130), .b(n_2129), .c(n_2128), .o(n_2472) );
in01f80 g737041 ( .a(n_43128), .o(n_43216) );
in01f80 newInst_3426 ( .a(newNet_3425), .o(newNet_3426) );
no02f80 g740503 ( .a(n_39711), .b(n_39655), .o(n_39727) );
no02f80 g739214 ( .a(n_40705), .b(n_40704), .o(n_40706) );
oa22f80 FE_RC_3204_0 ( .a(n_1118), .b(FE_OCPN875_n_44672), .c(n_1068), .d(n_44637), .o(n_1289) );
no02f80 g749877 ( .a(n_31311), .b(n_31371), .o(n_31409) );
in01f80 g756093 ( .a(n_24262), .o(n_24281) );
in01f80 newInst_2150 ( .a(newNet_2149), .o(newNet_2150) );
na02f80 g779746 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .o(n_1580) );
na02f80 g776560 ( .a(n_4286), .b(n_4345), .o(n_4424) );
no02f80 g765536 ( .a(n_14987), .b(n_15012), .o(n_15075) );
no02f80 g742913 ( .a(n_37073), .b(n_37072), .o(n_37322) );
in01f80 g761793 ( .a(n_18645), .o(n_18646) );
oa22f80 FE_RC_3208_0 ( .a(n_1001), .b(FE_OCPN875_n_44672), .c(FE_RN_1426_0), .d(n_44637), .o(n_1332) );
na02f80 g774499 ( .a(n_6524), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .o(n_6561) );
na02f80 g755866 ( .a(n_25548), .b(n_25054), .o(n_25110) );
na02f80 g774921 ( .a(n_6257), .b(n_6141), .o(n_6276) );
in01f80 newInst_2307 ( .a(newNet_2024), .o(newNet_2307) );
in01f80 g748347 ( .a(n_31796), .o(n_31797) );
oa12f80 g766041 ( .a(n_14686), .b(n_14689), .c(n_14685), .o(n_14740) );
in01f80 FE_RC_1557_0 ( .a(FE_OCP_RBN2290_n_2438), .o(FE_RN_441_0) );
in01f80 g765374 ( .a(n_16302), .o(n_16303) );
oa12f80 g754199 ( .a(n_25618), .b(n_26016), .c(n_25749), .o(n_26040) );
na02f80 g741008 ( .a(n_38969), .b(n_38968), .o(n_38970) );
na02f80 g738586 ( .a(n_41461), .b(n_41419), .o(n_41736) );
na02f80 g741260 ( .a(n_39148), .b(n_39118), .o(n_39226) );
no02f80 g739376 ( .a(n_41107), .b(n_41078), .o(n_41183) );
na02f80 g765305 ( .a(n_15710), .b(n_15969), .o(n_15962) );
na02f80 g750456 ( .a(n_29482), .b(n_25738), .o(n_29532) );
in01f80 newInst_2219 ( .a(newNet_2218), .o(newNet_2219) );
in01f80 g744788 ( .a(n_35148), .o(n_35175) );
na02f80 g755487 ( .a(n_24648), .b(n_24620), .o(n_24754) );
na02f80 g763924 ( .a(n_17018), .b(FE_OCP_RBN3359_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17257) );
na02f80 g768494 ( .a(n_12352), .b(n_11899), .o(n_12394) );
na02f80 g744550 ( .a(n_35397), .b(n_35396), .o(n_35398) );
na02f80 g746316 ( .a(n_33635), .b(n_33271), .o(n_33655) );
no02f80 g737937 ( .a(n_42201), .b(n_42108), .o(n_42298) );
ao12f80 g739219 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_21_), .b(n_45181), .c(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n_40681) );
no02f80 g766566 ( .a(n_14020), .b(n_13982), .o(n_14088) );
in01f80 g761983 ( .a(n_18284), .o(n_18704) );
no02f80 g748219 ( .a(n_32780), .b(n_32763), .o(n_32764) );
in01f80 newInst_1681 ( .a(newNet_192), .o(newNet_1681) );
in01f80 g753641 ( .a(n_26718), .o(n_26719) );
oa12f80 g737205 ( .a(n_42351), .b(n_42975), .c(n_42342), .o(n_42983) );
in01f80 FE_RC_2492_0 ( .a(delay_xor_ln23_unr3_stage2_stallmux_q), .o(FE_RN_1009_0) );
no02f80 g771592 ( .a(n_8923), .b(n_8309), .o(n_8973) );
no02f80 g764378 ( .a(n_16285), .b(n_14730), .o(n_16321) );
in01f80 FE_OCP_RBC1687_n_18986 ( .a(FE_OCP_RBN1685_n_18986), .o(FE_OCP_RBN1687_n_18986) );
no02f80 g784706 ( .a(n_11308), .b(FE_OCP_RBN2821_n_10023), .o(n_47182) );
no02f80 g769130 ( .a(n_11628), .b(n_11589), .o(n_11741) );
in01f80 newInst_2871 ( .a(newNet_2870), .o(newNet_2871) );
in01f80 g767728 ( .a(n_13440), .o(n_13441) );
no02f80 g754806 ( .a(n_26008), .b(n_25309), .o(n_26161) );
ao22s80 FE_RC_529_0 ( .a(n_28643), .b(n_28978), .c(n_28644), .d(n_28977), .o(n_29062) );
no02f80 g751038 ( .a(n_30092), .b(n_30091), .o(n_30093) );
na02f80 g745257 ( .a(n_34275), .b(n_34264), .o(n_34265) );
no02f80 g778015 ( .a(n_3021), .b(n_3051), .o(n_4719) );
in01f80 newInst_2442 ( .a(newNet_2441), .o(newNet_2442) );
no02f80 g747163 ( .a(n_32869), .b(n_32852), .o(n_32953) );
in01f80 FE_OCP_RBC3294_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3294_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
ao12f80 g736575 ( .a(n_43162), .b(n_43446), .c(n_43529), .o(n_43569) );
no02f80 g771783 ( .a(n_8863), .b(n_7592), .o(n_8885) );
no02f80 g739471 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n_40716) );
in01f80 g769317 ( .a(n_11972), .o(n_12050) );
in01f80 g750928 ( .a(n_30233), .o(n_30234) );
in01f80 FE_OCPC1507_n_23414 ( .a(n_23414), .o(FE_OCPN1507_n_23414) );
na02f80 g741403 ( .a(n_38811), .b(n_38067), .o(n_38841) );
na02f80 g765509 ( .a(n_15599), .b(n_15631), .o(n_15632) );
in01f80 g738511 ( .a(n_41696), .o(n_41668) );
na02f80 g736986 ( .a(n_43242), .b(n_43003), .o(n_43454) );
ao12f80 g738308 ( .a(n_41738), .b(n_41737), .c(n_41736), .o(n_41796) );
in01f80 newInst_3333 ( .a(newNet_1261), .o(newNet_3333) );
na02f80 g743697 ( .a(n_37382), .b(n_37381), .o(n_37383) );
no02f80 g784591 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n_46414) );
oa22f80 g744708 ( .a(n_36477), .b(n_36217), .c(n_36478), .d(n_36218), .o(n_36528) );
na02f80 g740231 ( .a(n_39764), .b(n_39763), .o(n_39795) );
in01f80 g772344 ( .a(n_8585), .o(n_8629) );
na02f80 g752180 ( .a(n_27921), .b(n_44735), .o(n_27976) );
in01f80 g749429 ( .a(n_30541), .o(n_30540) );
na02f80 g747005 ( .a(n_32833), .b(n_32801), .o(n_33025) );
no02f80 g760773 ( .a(n_19566), .b(n_19565), .o(n_19567) );
no02f80 g745095 ( .a(n_34897), .b(n_34896), .o(n_34898) );
in01f80 g779348 ( .a(n_1672), .o(n_1716) );
na02f80 g739440 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .o(n_40720) );
no02f80 g762287 ( .a(n_18444), .b(n_18452), .o(n_18626) );
in01f80 g772375 ( .a(n_8553), .o(n_8574) );
no02f80 g764865 ( .a(n_15554), .b(n_15547), .o(n_15621) );
in01f80 g760687 ( .a(n_19772), .o(n_19773) );
na02f80 g749265 ( .a(FE_OCP_RBN2829_n_30731), .b(FE_OCP_RBN2807_n_30643), .o(n_30803) );
ms00f80 delay_xor_ln23_unr3_stage2_stallmux_q_reg ( .ck(newNet_132), .d(n_44626), .o(delay_xor_ln23_unr3_stage2_stallmux_q) );
in01f80 g775785 ( .a(n_5490), .o(n_5491) );
no02f80 g771475 ( .a(n_9305), .b(n_9304), .o(n_9402) );
no02f80 g737027 ( .a(n_43032), .b(n_43031), .o(n_43066) );
in01f80 fopt782968 ( .a(n_41311), .o(n_44430) );
no02f80 g743091 ( .a(n_36951), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37097) );
oa12f80 g744533 ( .a(n_35439), .b(n_35438), .c(n_35437), .o(n_35464) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_16_ ( .ck(newNet_1865), .d(n_16767), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_) );
in01f80 FE_OCPC911_n_43022 ( .a(FE_OCPN910_n_43022), .o(FE_OCPN911_n_43022) );
ao22s80 g736371 ( .a(n_43820), .b(n_43516), .c(n_43821), .d(n_43517), .o(n_43853) );
ao12f80 g772279 ( .a(n_7531), .b(n_8409), .c(n_7559), .o(n_8471) );
oa12f80 g745696 ( .a(n_34109), .b(n_34191), .c(n_34134), .o(n_34250) );
in01f80 g772893 ( .a(n_7969), .o(n_7970) );
in01f80 g751184 ( .a(n_29881), .o(n_29850) );
in01f80 fopt782864 ( .a(n_21985), .o(n_44296) );
na02f80 g767805 ( .a(n_13065), .b(n_12996), .o(n_13066) );
no02f80 g745156 ( .a(n_34574), .b(n_34287), .o(n_34683) );
na02f80 g772810 ( .a(n_8100), .b(n_8099), .o(n_8224) );
no03m80 FE_RC_3807_0 ( .a(n_31947), .b(n_31992), .c(n_31993), .o(n_32021) );
in01f80 g754519 ( .a(n_26313), .o(n_26314) );
in01f80 g736722 ( .a(n_43281), .o(n_43372) );
na02f80 g765963 ( .a(n_14669), .b(n_14632), .o(n_14699) );
in01f80 FE_OCP_RBC3680_n_10338 ( .a(n_10338), .o(FE_OCP_RBN3680_n_10338) );
na02f80 g737735 ( .a(n_42392), .b(n_41994), .o(n_42434) );
no02f80 g765884 ( .a(FE_OCP_RBN2695_n_14814), .b(n_14758), .o(n_14879) );
no02f80 g740040 ( .a(n_40254), .b(n_40047), .o(n_40293) );
in01f80 g763418 ( .a(n_17132), .o(n_17121) );
na02f80 g773102 ( .a(FE_OCP_RBN3453_FE_OCPN1240_n_7721), .b(n_7950), .o(n_8110) );
in01f80 newInst_1794 ( .a(newNet_1793), .o(newNet_1794) );
no02f80 g778174 ( .a(n_2864), .b(n_2863), .o(n_2902) );
na02f80 g778197 ( .a(n_2692), .b(n_2691), .o(n_2693) );
in01f80 g770699 ( .a(n_10022), .o(n_10063) );
na02f80 g762923 ( .a(n_17679), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .o(n_17766) );
in01f80 g746284 ( .a(n_33640), .o(n_35268) );
na02f80 g763711 ( .a(n_16710), .b(n_16709), .o(n_16810) );
na02f80 g760990 ( .a(n_19250), .b(n_19215), .o(n_19353) );
oa12f80 g761953 ( .a(n_18735), .b(n_18911), .c(n_18533), .o(n_18994) );
no02f80 FE_RC_2828_0 ( .a(FE_RN_1213_0), .b(FE_RN_1214_0), .o(FE_RN_1215_0) );
in01f80 newInst_1579 ( .a(newNet_1578), .o(newNet_1579) );
na02f80 g766156 ( .a(n_14513), .b(n_14477), .o(n_14645) );
in01f80 g751964 ( .a(n_28864), .o(n_29042) );
in01f80 newInst_70 ( .a(newNet_69), .o(newNet_70) );
na02f80 g779295 ( .a(n_1658), .b(n_1039), .o(n_1744) );
na02f80 g759283 ( .a(n_20944), .b(n_20943), .o(n_20976) );
na02f80 g738064 ( .a(n_42145), .b(n_42141), .o(n_42142) );
in01f80 newInst_3331 ( .a(newNet_3330), .o(newNet_3331) );
no02f80 g761146 ( .a(n_19148), .b(n_17900), .o(n_19172) );
na02f80 g751401 ( .a(n_28652), .b(n_28533), .o(n_28653) );
in01f80 g770518 ( .a(n_10551), .o(n_10633) );
in01f80 g747784 ( .a(n_32260), .o(n_32261) );
ao12f80 g778257 ( .a(n_2576), .b(n_2575), .c(n_2574), .o(n_3911) );
oa12f80 g771482 ( .a(n_9189), .b(n_9077), .c(n_9074), .o(n_9208) );
oa12f80 g744560 ( .a(n_36121), .b(n_36623), .c(n_36050), .o(n_36683) );
no02f80 g759400 ( .a(n_20972), .b(n_20488), .o(n_21037) );
in01f80 g770321 ( .a(n_10690), .o(n_10691) );
oa12f80 g758600 ( .a(n_21842), .b(n_21898), .c(n_21783), .o(n_21950) );
na02f80 g739886 ( .a(n_40199), .b(n_39987), .o(n_40232) );
no02f80 g776951 ( .a(n_3758), .b(n_3529), .o(n_3789) );
no02f80 g766344 ( .a(n_14162), .b(n_14193), .o(n_14328) );
in01f80 g775807 ( .a(n_5461), .o(n_5462) );
in01f80 g747985 ( .a(n_31883), .o(n_31884) );
na02f80 g771137 ( .a(n_9509), .b(FE_OCPN1253_n_8348), .o(n_9670) );
na02f80 g754122 ( .a(FE_OCP_RBN2837_FE_RN_745_0), .b(n_25947), .o(n_26061) );
no02f80 g754980 ( .a(n_25414), .b(n_25482), .o(n_25504) );
no02f80 g752940 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .o(n_27878) );
no02f80 g746264 ( .a(n_33508), .b(n_33063), .o(n_33531) );
in01f80 g745120 ( .a(n_36232), .o(n_36233) );
no02f80 g764612 ( .a(n_16001), .b(n_15946), .o(n_16036) );
na02f80 g764289 ( .a(n_16333), .b(FE_OCPN3775_n_14730), .o(n_16442) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_24_ ( .ck(newNet_1503), .d(n_32256), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_) );
no02f80 g772750 ( .a(n_8234), .b(n_8209), .o(n_8351) );
na02f80 g759506 ( .a(n_20595), .b(n_20468), .o(n_20596) );
ao12f80 g759080 ( .a(n_21017), .b(n_21164), .c(n_21092), .o(n_21195) );
in01f80 g768438 ( .a(n_12450), .o(n_12481) );
in01f80 g743362 ( .a(n_36690), .o(n_36691) );
in01f80 g768486 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .o(n_12318) );
in01f80 g760268 ( .a(n_20456), .o(n_20537) );
no02f80 g751059 ( .a(n_30332), .b(n_29836), .o(n_30433) );
no02f80 g740847 ( .a(n_39379), .b(n_39400), .o(n_39841) );
na02f80 g745804 ( .a(n_44133), .b(n_34122), .o(n_34328) );
ao12f80 g752057 ( .a(n_28114), .b(n_28059), .c(n_27910), .o(n_28186) );
ao12f80 g746841 ( .a(n_33264), .b(FE_OCP_RBN3384_n_33108), .c(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n_33287) );
na02f80 g766899 ( .a(n_13685), .b(n_13684), .o(n_13686) );
na02f80 g778245 ( .a(n_2724), .b(n_2670), .o(n_2760) );
na03f80 g765168 ( .a(n_15407), .b(FE_OCP_RBN2737_n_15300), .c(n_15410), .o(n_15492) );
na02f80 g744523 ( .a(n_35421), .b(n_35420), .o(n_35440) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_14_ ( .ck(newNet_1339), .d(n_1207), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_) );
ao12f80 g741884 ( .a(n_38339), .b(n_38338), .c(n_38337), .o(n_38468) );
in01f80 fopt783245 ( .a(n_40736), .o(n_44800) );
in01f80 newInst_1786 ( .a(newNet_1785), .o(newNet_1786) );
na02f80 g753893 ( .a(n_26361), .b(FE_OCPN1498_n_26360), .o(n_26461) );
oa12f80 g760889 ( .a(n_20119), .b(n_20118), .c(n_20117), .o(n_20198) );
in01f80 newInst_932 ( .a(newNet_217), .o(newNet_932) );
in01f80 g737886 ( .a(n_42307), .o(n_42279) );
na02f80 g753954 ( .a(n_26194), .b(n_23447), .o(n_26363) );
in01f80 newInst_3187 ( .a(newNet_3186), .o(newNet_3187) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_26_ ( .ck(newNet_1212), .d(n_6229), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_) );
no02f80 g779787 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n_1445) );
in01f80 newInst_2258 ( .a(newNet_1918), .o(newNet_2258) );
in01f80 newInst_961 ( .a(newNet_358), .o(newNet_961) );
na02f80 g770614 ( .a(n_10313), .b(n_10264), .o(n_10338) );
na02f80 g760172 ( .a(n_20290), .b(n_20227), .o(n_20291) );
na02f80 g739290 ( .a(n_40713), .b(n_40766), .o(n_40768) );
no02f80 g784410 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .o(n_46222) );
no02f80 g764563 ( .a(n_45332), .b(n_16080), .o(n_16082) );
in01f80 FE_OCPC1793_n_30612 ( .a(n_30612), .o(FE_OCPN1793_n_30612) );
in01f80 g753720 ( .a(n_26532), .o(n_26533) );
in01f80 newInst_3647 ( .a(newNet_3646), .o(newNet_3647) );
in01f80 newInst_894 ( .a(newNet_866), .o(newNet_894) );
in01f80 g752637 ( .a(n_28239), .o(n_28240) );
na02f80 g771687 ( .a(n_9125), .b(FE_OCP_RBN2336_n_8269), .o(n_9237) );
no02f80 g749437 ( .a(n_30576), .b(n_30562), .o(n_30643) );
in01f80 newInst_2585 ( .a(newNet_2584), .o(newNet_2585) );
in01f80 g748743 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n_32462) );
in01f80 g775068 ( .a(n_6108), .o(n_6109) );
no02f80 g775124 ( .a(n_5839), .b(n_5769), .o(n_5878) );
na02f80 FE_RC_3630_0 ( .a(n_13642), .b(n_13683), .o(FE_RN_1591_0) );
in01f80 g738817 ( .a(n_41386), .o(n_41382) );
in01f80 g755857 ( .a(n_24958), .o(n_25059) );
in01f80 g750275 ( .a(n_29787), .o(n_29829) );
in01f80 g747499 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .o(n_32387) );
na02f80 g771582 ( .a(n_8881), .b(n_8880), .o(n_8985) );
no02f80 g750689 ( .a(n_29265), .b(n_29143), .o(n_29302) );
na02f80 g751390 ( .a(n_29363), .b(n_29336), .o(n_29337) );
in01f80 newInst_1291 ( .a(newNet_1290), .o(newNet_1291) );
in01f80 FE_OCP_RBC3019_n_31117 ( .a(FE_OCP_RBN3015_n_31117), .o(FE_OCP_RBN3019_n_31117) );
na02f80 g773192 ( .a(n_7802), .b(n_8062), .o(n_8036) );
in01f80 g770870 ( .a(n_10212), .o(n_10334) );
na02f80 g746034 ( .a(n_33780), .b(n_32985), .o(n_33880) );
in01f80 g744534 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .o(n_36745) );
in01f80 g746805 ( .a(n_33215), .o(n_33216) );
in01f80 newInst_3401 ( .a(newNet_3400), .o(newNet_3401) );
in01f80 newInst_1186 ( .a(newNet_225), .o(newNet_1186) );
na02f80 g761551 ( .a(n_18861), .b(FE_OCP_DRV_N1546_n_18860), .o(n_18863) );
na02f80 g741181 ( .a(FE_OCP_RBN2636_n_38806), .b(n_38964), .o(n_39013) );
in01f80 newInst_1349 ( .a(newNet_1091), .o(newNet_1349) );
ao22s80 g747087 ( .a(n_32904), .b(n_32931), .c(n_32903), .d(n_32888), .o(n_32985) );
in01f80 g743481 ( .a(n_36632), .o(n_36611) );
na02f80 g761432 ( .a(n_18897), .b(n_18335), .o(n_18923) );
ao12f80 g760167 ( .a(n_20902), .b(n_20929), .c(n_20901), .o(n_21514) );
oa12f80 g759539 ( .a(n_20798), .b(n_20820), .c(n_20797), .o(n_20915) );
na02f80 g776475 ( .a(n_4391), .b(n_4318), .o(n_4443) );
in01f80 g763042 ( .a(n_17460), .o(n_17456) );
no02f80 g769221 ( .a(n_11439), .b(n_45300), .o(n_11437) );
na02f80 g741997 ( .a(n_38352), .b(n_38312), .o(n_38376) );
ao22s80 FE_RC_927_0 ( .a(n_25534), .b(n_25903), .c(n_25902), .d(n_25533), .o(n_25999) );
in01f80 g752311 ( .a(n_29109), .o(n_27914) );
in01f80 g750964 ( .a(n_30229), .o(n_30230) );
in01f80 newInst_653 ( .a(newNet_652), .o(newNet_653) );
in01f80 newInst_310 ( .a(newNet_104), .o(newNet_310) );
no02f80 g747617 ( .a(n_45755), .b(n_47272), .o(n_32333) );
ao22s80 FE_RC_670_0 ( .a(n_45314), .b(n_6571), .c(n_6642), .d(n_6649), .o(n_6759) );
no02f80 g739343 ( .a(n_45146), .b(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n_40707) );
in01f80 newInst_2896 ( .a(newNet_523), .o(newNet_2896) );
in01f80 g780609 ( .a(n_746), .o(n_747) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_0_ ( .ck(newNet_1350), .d(n_419), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_) );
oa12f80 g780798 ( .a(n_383), .b(n_386), .c(n_382), .o(n_412) );
in01f80 g780730 ( .a(n_609), .o(n_619) );
oa12f80 g762463 ( .a(n_17966), .b(n_18070), .c(n_17912), .o(n_18130) );
na02f80 g758267 ( .a(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .o(n_22643) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_5_ ( .ck(newNet_1283), .d(n_1133), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_) );
in01f80 g742403 ( .a(n_37838), .o(n_37823) );
in01f80 g738049 ( .a(n_42154), .o(n_42155) );
no02f80 g776171 ( .a(n_4655), .b(FE_OCPN846_n_4046), .o(n_4843) );
in01f80 g743258 ( .a(n_36864), .o(n_36865) );
no03m80 g752052 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .b(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .c(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .o(n_27978) );
oa12f80 g761828 ( .a(n_19071), .b(n_19097), .c(n_19070), .o(n_19758) );
in01f80 FE_OCP_RBC2198_n_41256 ( .a(n_41256), .o(FE_OCP_RBN2198_n_41256) );
no02f80 g762376 ( .a(FE_OFN750_n_45003), .b(n_18572), .o(n_18765) );
na02f80 g775625 ( .a(n_5460), .b(n_5425), .o(n_5504) );
na02f80 g777076 ( .a(n_3825), .b(n_3794), .o(n_4208) );
oa12f80 g772627 ( .a(n_8251), .b(n_8275), .c(n_8159), .o(n_8276) );
in01f80 g757306 ( .a(n_23450), .o(n_23451) );
in01f80 g776424 ( .a(n_4397), .o(n_4468) );
na02f80 g753489 ( .a(n_26851), .b(n_26850), .o(n_26875) );
in01f80 newInst_3624 ( .a(newNet_3623), .o(newNet_3624) );
in01f80 g770058 ( .a(n_11008), .o(n_11019) );
ao12f80 g768475 ( .a(n_12355), .b(n_45659), .c(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .o(n_12581) );
in01f80 g761458 ( .a(n_19651), .o(n_19652) );
in01f80 g737716 ( .a(n_42389), .o(n_42448) );
in01f80 g780714 ( .a(n_748), .o(n_633) );
no02f80 g739975 ( .a(n_39929), .b(n_39818), .o(n_39959) );
in01f80 g778340 ( .a(n_2526), .o(n_2527) );
na02f80 g745027 ( .a(n_34792), .b(n_34538), .o(n_34878) );
in01f80 g738703 ( .a(n_41533), .o(n_41663) );
no02f80 g778264 ( .a(n_4073), .b(n_2976), .o(n_2997) );
na02f80 g765199 ( .a(n_15157), .b(n_15081), .o(n_15196) );
na02f80 g774781 ( .a(n_6352), .b(n_6325), .o(n_6453) );
in01f80 FE_OCP_RBC2842_n_4784 ( .a(n_4784), .o(FE_OCP_RBN2842_n_4784) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_2_ ( .ck(newNet_2629), .d(n_21066), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_) );
oa22f80 FE_RC_1417_0 ( .a(n_45066), .b(n_20462), .c(n_45012), .d(n_20461), .o(n_20636) );
in01f80 FE_OCP_DRV_C1543_n_18854 ( .a(n_18854), .o(FE_OCP_DRV_N1543_n_18854) );
in01f80 g750934 ( .a(n_29059), .o(n_29913) );
in01f80 newInst_2455 ( .a(newNet_727), .o(newNet_2455) );
no02f80 g761099 ( .a(n_19147), .b(n_19113), .o(n_19243) );
no02f80 g770815 ( .a(n_9944), .b(n_44464), .o(n_10025) );
in01f80 g760114 ( .a(n_20337), .o(n_20338) );
no02f80 g751459 ( .a(n_28521), .b(n_28571), .o(n_28603) );
ao12f80 g762459 ( .a(n_18137), .b(FE_OCP_RBN2147_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .o(n_17973) );
na02f80 g758120 ( .a(FE_OCPN1249_n_44267), .b(n_21339), .o(n_22305) );
na02f80 g737964 ( .a(n_42182), .b(n_42181), .o(n_42183) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_16_ ( .ck(newNet_1335), .d(n_1224), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_) );
na02f80 g760178 ( .a(n_20456), .b(n_19664), .o(n_20660) );
na02f80 g754753 ( .a(n_26161), .b(n_26134), .o(n_26135) );
in01f80 FE_RC_2968_0 ( .a(n_25670), .o(FE_RN_1297_0) );
na02f80 g765967 ( .a(n_45520), .b(FE_OCP_RBN3528_n_13765), .o(n_14859) );
in01f80 FE_OCPC845_n_4046 ( .a(n_4046), .o(FE_OCPN845_n_4046) );
oa12f80 g771550 ( .a(n_8880), .b(n_8871), .c(FE_OCP_RBN3472_n_7886), .o(n_8976) );
na02f80 g751823 ( .a(FE_OCP_RBN2164_n_28249), .b(n_28088), .o(n_28283) );
no02f80 g746080 ( .a(n_33755), .b(n_33691), .o(n_33809) );
ao22s80 g784430 ( .a(n_36773), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_46242) );
na02f80 g760604 ( .a(n_19774), .b(n_19704), .o(n_19841) );
in01f80 g779769 ( .a(n_1479), .o(n_1410) );
na02f80 g737296 ( .a(n_42875), .b(n_42885), .o(n_42941) );
in01f80 FE_OFC812_n_2405 ( .a(FE_OFN829_n_2405), .o(FE_OFN812_n_2405) );
ms00f80 cos_out_reg_4_ ( .ck(newNet_3684), .d(n_43694), .o(cos_out_4) );
in01f80 FE_RC_306_0 ( .a(n_21269), .o(FE_RN_90_0) );
na02f80 g744281 ( .a(n_44180), .b(n_34925), .o(n_35732) );
na02f80 g739221 ( .a(n_40742), .b(n_40694), .o(n_40783) );
in01f80 newInst_1530 ( .a(newNet_1529), .o(newNet_1530) );
na02f80 g745390 ( .a(n_34463), .b(n_34411), .o(n_34514) );
ao12f80 g752830 ( .a(n_28199), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n_28753) );
in01f80 newInst_503 ( .a(newNet_502), .o(newNet_503) );
oa12f80 g765803 ( .a(n_14390), .b(n_15290), .c(n_14345), .o(n_15324) );
no02f80 g745296 ( .a(n_35888), .b(n_35839), .o(n_35889) );
ao22s80 FE_RC_3344_0 ( .a(n_25623), .b(n_26000), .c(n_25622), .d(n_26022), .o(n_26152) );
in01f80 g774874 ( .a(n_6205), .o(n_6247) );
in01f80 g750713 ( .a(n_29322), .o(n_29495) );
na02f80 g742559 ( .a(n_37619), .b(n_37618), .o(n_37638) );
oa22f80 g743635 ( .a(n_36394), .b(n_35738), .c(n_36395), .d(n_35737), .o(n_36442) );
no02f80 g746936 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n_32948) );
na02f80 g738341 ( .a(n_41771), .b(n_41345), .o(n_41795) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_19_ ( .ck(newNet_3232), .d(n_36469), .o(delay_add_ln22_unr23_stage9_stallmux_q_19_) );
ao12f80 g778965 ( .a(n_2094), .b(n_2093), .c(n_2092), .o(n_2140) );
no02f80 g757185 ( .a(n_23193), .b(n_23192), .o(n_23215) );
na02f80 g777322 ( .a(n_4759), .b(n_5197), .o(n_5368) );
na02f80 g772647 ( .a(n_8289), .b(n_8281), .o(n_8282) );
ms00f80 cos_out_reg_17_ ( .ck(newNet_3737), .d(n_43852), .o(cos_out_17) );
na02f80 g759637 ( .a(n_20640), .b(n_45012), .o(n_20683) );
na02f80 g739797 ( .a(n_40406), .b(n_39976), .o(n_40425) );
in01f80 newInst_185 ( .a(newNet_184), .o(newNet_185) );
no02f80 g776328 ( .a(n_4363), .b(n_4416), .o(n_4453) );
in01f80 g742784 ( .a(n_37875), .o(n_37334) );
in01f80 newInst_994 ( .a(newNet_993), .o(newNet_994) );
oa12f80 g768970 ( .a(n_11976), .b(n_11866), .c(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12053) );
in01f80 FE_OCPC917_n_46991 ( .a(FE_OCPN916_n_46991), .o(FE_OCPN917_n_46991) );
na02f80 g781095 ( .a(n_252), .b(n_251), .o(n_253) );
in01f80 g751929 ( .a(n_28207), .o(n_28208) );
in01f80 g773176 ( .a(n_7963), .o(n_8012) );
na02f80 g778600 ( .a(n_2423), .b(n_2402), .o(n_2424) );
na02f80 g740343 ( .a(n_40169), .b(n_40205), .o(n_40306) );
no02f80 g752820 ( .a(n_27168), .b(n_27236), .o(n_27357) );
na02f80 g747834 ( .a(n_33571), .b(n_33511), .o(n_33667) );
oa12f80 g745959 ( .a(n_35280), .b(n_35299), .c(n_35279), .o(n_35335) );
na02f80 g739963 ( .a(n_40121), .b(n_40044), .o(n_40228) );
in01f80 newInst_1598 ( .a(newNet_1175), .o(newNet_1598) );
oa12f80 g753746 ( .a(n_26711), .b(n_27097), .c(n_26571), .o(n_27132) );
oa12f80 g740785 ( .a(n_39080), .b(n_39354), .c(n_39081), .o(n_39408) );
no02f80 g779533 ( .a(n_1643), .b(n_1801), .o(n_1741) );
oa12f80 g772825 ( .a(n_7371), .b(n_7798), .c(n_7341), .o(n_7905) );
ao22s80 g736517 ( .a(n_43640), .b(n_43607), .c(n_43639), .d(n_43608), .o(n_43672) );
in01f80 FE_RC_2423_0 ( .a(n_6737), .o(FE_RN_960_0) );
in01f80 g772755 ( .a(n_8043), .o(n_8044) );
no02f80 g761070 ( .a(n_19172), .b(n_19111), .o(n_19211) );
in01f80 g741893 ( .a(n_38190), .o(n_38191) );
in01f80 fopt782728 ( .a(n_44100), .o(n_44101) );
in01f80 g760807 ( .a(n_19538), .o(n_19560) );
in01f80 FE_OCP_RBC3012_n_31117 ( .a(FE_OCP_RBN3702_n_31064), .o(FE_OCP_RBN3012_n_31117) );
no02f80 g767326 ( .a(n_13454), .b(FE_OCPN860_n_12880), .o(n_13499) );
in01f80 g763897 ( .a(n_17302), .o(n_17422) );
no02f80 g748262 ( .a(FE_OCP_RBN3085_n_31819), .b(FE_OCP_RBN2804_n_30534), .o(n_32020) );
no02f80 FE_RC_1663_0 ( .a(FE_RN_462_0), .b(FE_OCP_RBN3391_n_37557), .o(FE_RN_464_0) );
na02f80 g743788 ( .a(n_37283), .b(n_46230), .o(n_37262) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_29_ ( .ck(newNet_2160), .d(n_1014), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_) );
ao12f80 g779166 ( .a(n_1875), .b(n_1874), .c(n_1873), .o(n_2218) );
oa12f80 g747639 ( .a(n_31821), .b(n_32150), .c(n_32149), .o(n_32172) );
in01f80 newInst_779 ( .a(newNet_778), .o(newNet_779) );
no02f80 g764201 ( .a(n_16484), .b(n_14784), .o(n_16583) );
no02f80 g747589 ( .a(n_32302), .b(n_47273), .o(n_32364) );
in01f80 newInst_3525 ( .a(newNet_512), .o(newNet_3525) );
no02f80 g754719 ( .a(FE_OCP_RBN2959_n_26231), .b(n_26544), .o(n_26571) );
na02f80 g764998 ( .a(n_15500), .b(n_15348), .o(n_15537) );
no02f80 g754144 ( .a(n_25972), .b(n_26002), .o(n_26027) );
na02f80 g758237 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .o(n_23052) );
in01f80 g770123 ( .a(n_10904), .o(n_10905) );
no02f80 g742984 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_14_), .o(n_37072) );
no02f80 g764976 ( .a(n_15933), .b(n_15563), .o(n_16066) );
no02f80 g741858 ( .a(n_38434), .b(n_38432), .o(n_38435) );
ao12f80 g777944 ( .a(n_3049), .b(n_3116), .c(n_2759), .o(n_3159) );
in01f80 g767077 ( .a(n_13642), .o(n_13643) );
no02f80 g763244 ( .a(n_17736), .b(n_17713), .o(n_17714) );
in01f80 g759468 ( .a(n_21055), .o(n_21056) );
oa12f80 g777741 ( .a(n_2909), .b(n_3291), .c(n_2838), .o(n_3354) );
oa22f80 g764231 ( .a(n_16575), .b(n_17584), .c(n_16551), .d(n_16338), .o(n_16619) );
in01f80 newInst_2917 ( .a(newNet_2916), .o(newNet_2917) );
no02f80 g780508 ( .a(n_667), .b(n_687), .o(n_708) );
no02f80 g737411 ( .a(n_42740), .b(n_42753), .o(n_43129) );
in01f80 g776783 ( .a(n_4115), .o(n_4116) );
na02f80 FE_RC_2328_0 ( .a(n_33034), .b(FE_RN_887_0), .o(FE_RN_888_0) );
in01f80 g781319 ( .a(n_65), .o(n_117) );
no02f80 g745867 ( .a(n_44102), .b(n_33939), .o(n_34266) );
oa12f80 g739782 ( .a(n_40256), .b(n_40470), .c(n_40060), .o(n_40496) );
no02f80 g749866 ( .a(FE_OCP_RBN3011_n_31117), .b(n_31214), .o(n_31324) );
oa22f80 FE_RC_783_0 ( .a(FE_OFN803_n_46285), .b(n_12143), .c(FE_OFN771_n_46337), .d(n_12067), .o(n_46358) );
in01f80 newInst_1222 ( .a(newNet_747), .o(newNet_1222) );
no02f80 g769027 ( .a(FE_OCP_RBN2119_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .o(n_11860) );
na02f80 g752394 ( .a(n_44759), .b(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .o(n_27821) );
in01f80 g763978 ( .a(FE_OFN779_n_17093), .o(n_19222) );
no02f80 g772776 ( .a(n_8157), .b(n_8176), .o(n_8266) );
na02f80 g780917 ( .a(n_521), .b(n_274), .o(n_582) );
no02f80 g778951 ( .a(n_2260), .b(n_1990), .o(n_2305) );
in01f80 g739463 ( .a(n_40672), .o(n_40673) );
in01f80 newInst_3145 ( .a(newNet_537), .o(newNet_3145) );
ao12f80 g748839 ( .a(n_32443), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n_32864) );
no02f80 g737019 ( .a(FE_OCP_RBN3729_n_43230), .b(n_43132), .o(n_43489) );
na02f80 g756490 ( .a(n_23676), .b(n_23733), .o(n_23763) );
in01f80 g749278 ( .a(n_30711), .o(n_30738) );
no02f80 g741571 ( .a(n_38658), .b(n_38778), .o(n_38715) );
oa12f80 g763049 ( .a(n_17554), .b(n_17588), .c(n_17553), .o(n_17643) );
in01f80 newInst_1611 ( .a(newNet_1610), .o(newNet_1611) );
oa12f80 g755758 ( .a(n_25221), .b(n_25259), .c(n_25160), .o(n_26234) );
na02f80 g741126 ( .a(n_39271), .b(n_38904), .o(n_39299) );
in01f80 g737050 ( .a(n_43204), .o(n_43245) );
na02f80 g759188 ( .a(n_21094), .b(n_19407), .o(n_21159) );
no02f80 g742633 ( .a(n_37424), .b(n_37423), .o(n_37425) );
in01f80 newInst_748 ( .a(newNet_747), .o(newNet_748) );
no02f80 g770892 ( .a(n_9868), .b(n_9909), .o(n_9965) );
ao12f80 g767535 ( .a(n_13307), .b(n_13306), .c(n_13305), .o(n_13875) );
na02f80 g775875 ( .a(n_47003), .b(n_47016), .o(n_5431) );
in01f80 newInst_2042 ( .a(newNet_2041), .o(newNet_2042) );
no02f80 g757953 ( .a(n_44267), .b(n_22201), .o(n_22313) );
oa22f80 FE_RC_424_0 ( .a(n_15071), .b(n_15161), .c(n_15160), .d(n_15072), .o(n_15314) );
na02f80 g770322 ( .a(n_10663), .b(n_44490), .o(n_10664) );
in01f80 g758763 ( .a(n_21893), .o(n_21894) );
in01f80 g744771 ( .a(n_35281), .o(n_35282) );
no02f80 g764573 ( .a(n_15993), .b(n_14650), .o(n_16046) );
in01f80 g778643 ( .a(n_3084), .o(n_2294) );
no02f80 g755624 ( .a(n_24548), .b(n_24458), .o(n_24615) );
na02f80 g755582 ( .a(n_24506), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24532) );
in01f80 g752774 ( .a(n_27158), .o(n_27159) );
oa12f80 g764470 ( .a(n_16270), .b(n_16269), .c(n_16268), .o(n_16362) );
in01f80 FE_OCP_RBC1919_n_22476 ( .a(n_22476), .o(FE_OCP_RBN1919_n_22476) );
in01f80 g772218 ( .a(n_8765), .o(n_8764) );
in01f80 newInst_3267 ( .a(newNet_2509), .o(newNet_3267) );
na02f80 g757812 ( .a(n_23183), .b(n_23116), .o(n_23184) );
in01f80 FE_RC_1413_0 ( .a(n_15688), .o(FE_RN_412_0) );
no02f80 g769933 ( .a(n_10948), .b(n_10891), .o(n_10971) );
no02f80 g740147 ( .a(n_39816), .b(n_39864), .o(n_39865) );
oa12f80 g766676 ( .a(n_14221), .b(n_14220), .c(n_14219), .o(n_15564) );
na02f80 g754865 ( .a(n_25668), .b(n_25667), .o(n_25723) );
no02f80 g769900 ( .a(n_10965), .b(n_10918), .o(n_10970) );
in01f80 g746957 ( .a(n_33246), .o(n_33247) );
na02f80 FE_RC_3996_0 ( .a(n_30178), .b(n_29969), .o(n_30283) );
in01f80 g747367 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .o(n_32637) );
na02f80 g749835 ( .a(FE_OCP_RBN3013_n_31117), .b(n_31116), .o(n_31536) );
no02f80 g739011 ( .a(n_41133), .b(n_46947), .o(n_41155) );
oa22f80 g780043 ( .a(n_1233), .b(n_896), .c(n_1232), .d(n_895), .o(n_1241) );
no02f80 g781171 ( .a(n_177), .b(n_264), .o(n_181) );
no02f80 g745585 ( .a(n_34297), .b(n_34292), .o(n_34377) );
in01f80 g764649 ( .a(n_15911), .o(n_15910) );
in01f80 g753100 ( .a(n_27465), .o(n_27466) );
oa12f80 g775894 ( .a(n_5209), .b(n_5208), .c(n_5207), .o(n_5363) );
in01f80 g750069 ( .a(n_30244), .o(n_30217) );
in01f80 g749946 ( .a(n_30239), .o(n_30240) );
na02f80 g766164 ( .a(n_14656), .b(n_14625), .o(n_14678) );
no02f80 g779639 ( .a(n_1512), .b(n_1420), .o(n_1497) );
in01f80 g770784 ( .a(n_10223), .o(n_10353) );
no02f80 FE_RC_1136_0 ( .a(FE_RN_342_0), .b(FE_RN_343_0), .o(FE_RN_344_0) );
oa22f80 g778756 ( .a(n_2170), .b(n_1772), .c(n_2171), .d(n_1771), .o(n_2620) );
oa12f80 g751854 ( .a(n_28919), .b(n_28921), .c(n_29026), .o(n_28990) );
in01f80 g738156 ( .a(n_42046), .o(n_42026) );
no02f80 g759989 ( .a(n_20539), .b(n_20491), .o(n_20582) );
oa22f80 FE_RC_617_0 ( .a(n_40598), .b(n_40579), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_44958), .o(n_40587) );
in01f80 g780869 ( .a(n_360), .o(n_361) );
na02f80 g738424 ( .a(n_41450), .b(n_41473), .o(n_41474) );
no02f80 g765790 ( .a(n_14923), .b(n_14956), .o(n_15018) );
no02f80 g766949 ( .a(n_14758), .b(n_14253), .o(n_14345) );
oa22f80 FE_RC_1677_0 ( .a(n_11181), .b(n_11222), .c(n_11221), .d(n_11217), .o(n_11308) );
ao12f80 g755244 ( .a(n_24842), .b(n_24975), .c(n_24803), .o(n_24990) );
ao12f80 g767629 ( .a(n_13020), .b(n_13019), .c(n_13018), .o(n_13134) );
in01f80 g742699 ( .a(n_37544), .o(n_37981) );
na02f80 g736315 ( .a(n_43859), .b(n_43641), .o(n_43876) );
in01f80 newInst_1677 ( .a(newNet_1676), .o(newNet_1677) );
in01f80 g771913 ( .a(n_8980), .o(n_8990) );
na02f80 g736750 ( .a(n_43553), .b(n_43186), .o(n_43285) );
in01f80 fopt783572 ( .a(n_40563), .o(n_45196) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_27_ ( .ck(newNet_2927), .d(n_6529), .o(delay_add_ln22_unr5_stage3_stallmux_q_27_) );
in01f80 g740451 ( .a(n_39776), .o(n_39777) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_25_ ( .ck(newNet_3612), .d(n_17759), .o(delay_add_ln22_unr11_stage5_stallmux_q_25_) );
no02f80 g756298 ( .a(n_24585), .b(n_23811), .o(n_24673) );
in01f80 FE_OCP_RBC2898_n_45484 ( .a(n_45484), .o(FE_OCP_RBN2898_n_45484) );
in01f80 newInst_3028 ( .a(newNet_1162), .o(newNet_3028) );
no02f80 g773424 ( .a(n_7565), .b(n_7564), .o(n_7566) );
ao22s80 FE_RC_3457_0 ( .a(FE_OCPN1410_n_27014), .b(n_30697), .c(n_30696), .d(FE_RN_1486_0), .o(n_30818) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_16_ ( .ck(newNet_1633), .d(n_27107), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_) );
na02f80 g762877 ( .a(n_17841), .b(delay_add_ln22_unr11_stage5_stallmux_q_8_), .o(n_17906) );
in01f80 g774028 ( .a(n_6874), .o(n_6875) );
in01f80 newInst_3618 ( .a(newNet_3617), .o(newNet_3618) );
ao12f80 g772613 ( .a(n_7697), .b(n_8289), .c(n_7827), .o(n_8557) );
ao12f80 g773512 ( .a(n_7471), .b(n_7470), .c(n_7469), .o(n_8568) );
na02f80 g781217 ( .a(n_143), .b(n_54), .o(n_160) );
na02f80 FE_RC_1847_0 ( .a(FE_RN_560_0), .b(FE_RN_562_0), .o(n_36272) );
in01f80 g777892 ( .a(n_3272), .o(n_3273) );
na02f80 g776971 ( .a(n_3743), .b(n_3813), .o(n_3849) );
na02f80 g769590 ( .a(n_11362), .b(n_11237), .o(n_11390) );
no02f80 g751046 ( .a(n_29822), .b(n_29819), .o(n_30003) );
na03f80 FE_RC_1213_0 ( .a(n_33367), .b(n_33851), .c(n_33852), .o(n_33876) );
no02f80 g763737 ( .a(n_17498), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n_17533) );
ao12f80 g784668 ( .a(n_5838), .b(n_5793), .c(n_5587), .o(n_46998) );
oa22f80 g779111 ( .a(n_1958), .b(n_1803), .c(n_1964), .d(n_1802), .o(n_2540) );
na02f80 g770096 ( .a(n_10861), .b(n_10822), .o(n_10959) );
ao12f80 g768562 ( .a(n_12243), .b(n_12242), .c(n_12241), .o(n_12850) );
ao12f80 g762054 ( .a(n_18589), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n_18629) );
no02f80 g768842 ( .a(n_45685), .b(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .o(n_12147) );
na02f80 g758241 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .o(n_22783) );
in01f80 g758641 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n_22456) );
ao12f80 g738546 ( .a(n_41387), .b(n_41407), .c(n_41406), .o(n_41453) );
no02f80 g762879 ( .a(n_17841), .b(delay_add_ln22_unr11_stage5_stallmux_q_8_), .o(n_17866) );
oa22f80 g739759 ( .a(n_40484), .b(n_40103), .c(n_40485), .d(n_40102), .o(n_40512) );
in01f80 g749801 ( .a(n_31534), .o(n_31535) );
no02f80 FE_RC_2790_0 ( .a(FE_RN_1190_0), .b(FE_RN_1192_0), .o(n_34261) );
na02f80 g775948 ( .a(n_5144), .b(n_5131), .o(n_5132) );
in01f80 newInst_457 ( .a(newNet_456), .o(newNet_457) );
in01f80 FE_OFC755_n_44461 ( .a(FE_OCP_RBN2616_n_44561), .o(FE_OFN755_n_44461) );
na02f80 g772885 ( .a(n_7929), .b(n_7635), .o(n_7971) );
na02f80 g777969 ( .a(n_3200), .b(n_3199), .o(n_3210) );
na02f80 g767818 ( .a(n_13065), .b(n_13041), .o(n_13761) );
in01f80 FE_RC_504_0 ( .a(n_22972), .o(FE_RN_153_0) );
no03m80 g747695 ( .a(n_33311), .b(n_33313), .c(n_33359), .o(n_33360) );
in01f80 g772316 ( .a(n_8760), .o(n_8690) );
na02f80 g767285 ( .a(n_13626), .b(n_13625), .o(n_13588) );
no02f80 g754575 ( .a(n_26308), .b(n_26311), .o(n_26743) );
na02f80 g753822 ( .a(n_26321), .b(FE_OCPN1488_n_23447), .o(n_26473) );
na02f80 g738419 ( .a(n_41814), .b(n_41632), .o(n_41963) );
in01f80 FE_RC_3458_0 ( .a(n_30790), .o(FE_RN_1487_0) );
na02f80 g773248 ( .a(n_7603), .b(n_7602), .o(n_7604) );
in01f80 newInst_3444 ( .a(newNet_3443), .o(newNet_3444) );
na02f80 FE_RC_4249_0 ( .a(FE_RN_1869_0), .b(n_26802), .o(n_26877) );
in01f80 newInst_2684 ( .a(newNet_2683), .o(newNet_2684) );
na02f80 g760685 ( .a(n_19638), .b(n_18032), .o(n_19705) );
na02f80 g770563 ( .a(FE_OCP_RBN2794_n_10106), .b(FE_OCP_RBN2529_n_9044), .o(n_10337) );
na02f80 g750884 ( .a(n_29054), .b(FE_OFN787_n_25834), .o(n_29110) );
na02f80 g742090 ( .a(FE_OCP_RBN3452_n_37945), .b(n_37760), .o(n_38181) );
ms00f80 sin_out_reg_9_ ( .ck(newNet_7), .d(n_43773), .o(sin_out_9) );
na02f80 g778767 ( .a(FE_OCP_RBN2289_n_2314), .b(n_2358), .o(n_2408) );
no02f80 g737477 ( .a(n_42564), .b(n_42662), .o(n_42701) );
in01f80 g763539 ( .a(n_16916), .o(n_16872) );
no02f80 g762042 ( .a(n_18226), .b(n_18075), .o(n_18227) );
in01f80 g769111 ( .a(n_11856), .o(n_11805) );
in01f80 newInst_3043 ( .a(newNet_3042), .o(newNet_3043) );
na02f80 g765208 ( .a(n_15338), .b(n_15337), .o(n_15378) );
in01f80 g738705 ( .a(n_41488), .o(n_41489) );
ao12f80 g784097 ( .a(n_45845), .b(n_45887), .c(FE_OCPN1754_n_7225), .o(n_45846) );
in01f80 newInst_2978 ( .a(newNet_385), .o(newNet_2978) );
no02f80 g761185 ( .a(n_19769), .b(n_19767), .o(n_19768) );
na02f80 g737589 ( .a(n_42663), .b(n_42584), .o(n_42683) );
no02f80 g763593 ( .a(n_17539), .b(n_17465), .o(n_17540) );
no02f80 g754510 ( .a(n_26740), .b(FE_OCP_RBN2966_n_26231), .o(n_26868) );
no02f80 g777704 ( .a(n_3340), .b(n_3152), .o(n_3360) );
ao12f80 g774198 ( .a(n_6998), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .o(n_7040) );
na02f80 g738551 ( .a(n_41448), .b(n_41382), .o(n_41506) );
no02f80 g762439 ( .a(n_18106), .b(delay_add_ln22_unr11_stage5_stallmux_q_14_), .o(n_18127) );
oa12f80 g749900 ( .a(n_30974), .b(n_30973), .c(n_30972), .o(n_31372) );
oa22f80 FE_RC_1540_0 ( .a(n_38201), .b(n_38506), .c(n_38460), .d(n_38202), .o(n_38537) );
in01f80 FE_OCPC1413_n_19715 ( .a(n_19715), .o(FE_OCPN1413_n_19715) );
na02f80 g778172 ( .a(n_2754), .b(n_2753), .o(n_2755) );
in01f80 g777835 ( .a(n_3264), .o(n_3265) );
na02f80 g773493 ( .a(n_45213), .b(n_8406), .o(n_7498) );
na02f80 g737719 ( .a(n_42367), .b(FE_OCP_RBN2443_n_42051), .o(n_42502) );
in01f80 g777422 ( .a(n_3596), .o(n_3705) );
no03m80 FE_RC_4141_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .c(n_32525), .o(FE_RN_1540_0) );
in01f80 g769419 ( .a(n_11582), .o(n_11575) );
na02f80 g744320 ( .a(n_35513), .b(n_34152), .o(n_35565) );
in01f80 FE_RC_1064_0 ( .a(n_37220), .o(FE_RN_313_0) );
oa22f80 g780058 ( .a(n_1229), .b(n_1062), .c(n_1228), .d(n_1063), .o(n_1237) );
ao12f80 g759135 ( .a(n_20838), .b(n_21018), .c(n_20815), .o(n_21090) );
na02f80 g737722 ( .a(n_42194), .b(n_41504), .o(n_42223) );
na02f80 g764689 ( .a(n_15703), .b(n_15409), .o(n_15774) );
in01f80 FE_OCP_RBC1700_n_19353 ( .a(FE_OCP_RBN1699_n_19353), .o(FE_OCP_RBN1700_n_19353) );
na02f80 g742373 ( .a(n_37768), .b(n_37799), .o(n_37819) );
no02f80 g780316 ( .a(n_964), .b(n_1079), .o(n_965) );
oa12f80 g746565 ( .a(n_34839), .b(n_34666), .c(n_34774), .o(n_35478) );
ao12f80 g762811 ( .a(n_17195), .b(n_17659), .c(n_17174), .o(n_17658) );
no02f80 g755480 ( .a(n_24778), .b(n_24518), .o(n_24782) );
in01f80 FE_OCP_RBC3734_n_31819 ( .a(FE_OCP_RBN3733_n_31819), .o(FE_OCP_RBN3734_n_31819) );
no02f80 g779622 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .o(n_2021) );
in01f80 g749975 ( .a(n_30275), .o(n_30276) );
no02f80 g763826 ( .a(n_17530), .b(n_17106), .o(n_17902) );
in01f80 g743397 ( .a(n_36703), .o(n_36704) );
no02f80 g754558 ( .a(n_26549), .b(n_26510), .o(n_26511) );
oa12f80 g756723 ( .a(n_23373), .b(n_23514), .c(n_23371), .o(n_23558) );
na02f80 g747599 ( .a(n_32241), .b(n_32221), .o(n_32305) );
no02f80 g763849 ( .a(n_16702), .b(FE_OCP_RBN2675_n_14991), .o(n_16751) );
no03m80 FE_RC_1529_0 ( .a(n_32635), .b(n_32754), .c(n_32731), .o(n_32772) );
no02f80 g755386 ( .a(n_25494), .b(n_24996), .o(n_25410) );
in01f80 FE_RC_1164_0 ( .a(n_28011), .o(FE_RN_351_0) );
no02f80 g777265 ( .a(n_3542), .b(FE_OCP_RBN2622_n_3601), .o(n_3672) );
na02f80 g773779 ( .a(n_7230), .b(n_7229), .o(n_7231) );
no02f80 g756081 ( .a(n_24183), .b(n_24182), .o(n_24184) );
ao12f80 g752733 ( .a(n_27192), .b(n_27193), .c(n_26958), .o(n_27237) );
no02f80 g775953 ( .a(n_4978), .b(n_4843), .o(n_4979) );
in01f80 g780885 ( .a(n_400), .o(n_401) );
in01f80 newInst_234 ( .a(newNet_233), .o(newNet_234) );
in01f80 g749017 ( .a(n_32312), .o(n_32313) );
in01f80 FE_RC_1936_0 ( .a(n_18848), .o(FE_RN_617_0) );
in01f80 FE_OCP_RBC2719_n_9182 ( .a(n_9182), .o(FE_OCP_RBN2719_n_9182) );
no02f80 g762398 ( .a(n_18421), .b(n_18417), .o(n_18499) );
in01f80 g749073 ( .a(n_31070), .o(n_31071) );
in01f80 g763131 ( .a(n_17294), .o(n_17290) );
na02f80 g740571 ( .a(FE_OCP_RBN2927_n_39614), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39657) );
no02f80 g755799 ( .a(n_24254), .b(n_21975), .o(n_24273) );
in01f80 g756610 ( .a(n_23629), .o(n_23656) );
na02f80 g746554 ( .a(n_34694), .b(n_34693), .o(n_34695) );
in01f80 g771518 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .o(n_9652) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_0_ ( .ck(newNet_602), .d(n_16619), .o(delay_xor_ln22_unr12_stage5_stallmux_q_0_) );
no02f80 g742514 ( .a(n_37515), .b(n_37514), .o(n_37516) );
in01f80 g760203 ( .a(n_20334), .o(n_20363) );
na02f80 g778366 ( .a(n_2790), .b(n_3594), .o(n_2809) );
na02f80 g775455 ( .a(n_5842), .b(n_47270), .o(n_5843) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_0_ ( .ck(newNet_765), .d(n_46165), .o(delay_xor_ln21_unr6_stage3_stallmux_q_0_) );
in01f80 newInst_2617 ( .a(newNet_2616), .o(newNet_2617) );
in01f80 g752695 ( .a(n_27440), .o(n_27441) );
in01f80 g773252 ( .a(n_7615), .o(n_7674) );
no02f80 g741819 ( .a(n_38341), .b(n_38220), .o(n_38418) );
na02f80 g771771 ( .a(n_9062), .b(FE_OCP_RBN3547_n_44575), .o(n_9119) );
oa22f80 g784357 ( .a(FE_OCP_RBN3075_FE_OFN807_n_46195), .b(n_5840), .c(FE_OFN86_n_46137), .d(n_5789), .o(n_46163) );
no02f80 g766733 ( .a(n_13725), .b(n_13690), .o(n_13731) );
in01f80 g748731 ( .a(n_31141), .o(n_31203) );
in01f80 newInst_368 ( .a(newNet_317), .o(newNet_368) );
no02f80 g780490 ( .a(n_743), .b(n_781), .o(n_1171) );
in01f80 g738681 ( .a(n_41685), .o(n_41686) );
na02f80 g749526 ( .a(n_30409), .b(n_30144), .o(n_30410) );
in01f80 g745608 ( .a(n_34704), .o(n_34651) );
in01f80 newInst_3610 ( .a(newNet_2007), .o(newNet_3610) );
oa22f80 g768715 ( .a(n_11922), .b(n_11799), .c(n_11923), .d(n_11800), .o(n_12068) );
na02f80 g745639 ( .a(n_34286), .b(n_33546), .o(n_34398) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_6_ ( .ck(newNet_401), .d(n_32594), .o(delay_xor_ln22_unr21_stage8_stallmux_q_6_) );
oa12f80 g746419 ( .a(n_33352), .b(n_33351), .c(n_33350), .o(n_34292) );
na02f80 g770626 ( .a(n_10425), .b(n_10424), .o(n_10426) );
no02f80 g760655 ( .a(n_19752), .b(FE_OCP_DRV_N1568_n_19751), .o(n_19837) );
ao22s80 g736321 ( .a(n_43808), .b(n_43619), .c(n_43807), .d(n_43620), .o(n_43858) );
in01f80 g755097 ( .a(n_25207), .o(n_25208) );
ao12f80 g779495 ( .a(n_1542), .b(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .o(n_1436) );
in01f80 FE_RC_1909_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(FE_RN_600_0) );
in01f80 g752273 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .o(n_28795) );
oa22f80 g751517 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_31_), .c(n_28460), .d(n_27824), .o(n_28824) );
in01f80 FE_RC_938_0 ( .a(n_22327), .o(FE_RN_276_0) );
in01f80 newInst_1285 ( .a(newNet_1242), .o(newNet_1285) );
na02f80 g763110 ( .a(n_17581), .b(n_17582), .o(n_17583) );
oa12f80 g742949 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36988), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .o(n_37252) );
in01f80 g776800 ( .a(n_4236), .o(n_4237) );
in01f80 newInst_2885 ( .a(newNet_372), .o(newNet_2885) );
oa22f80 g746456 ( .a(n_33291), .b(n_33265), .c(n_33255), .d(n_33266), .o(n_34293) );
no02f80 g736917 ( .a(FE_OCPN912_n_43022), .b(n_42748), .o(n_43538) );
in01f80 g755850 ( .a(n_24421), .o(n_24438) );
in01f80 g753377 ( .a(n_27110), .o(n_27287) );
oa12f80 g745040 ( .a(n_34851), .b(n_34873), .c(n_34850), .o(n_34924) );
oa22f80 FE_RC_1015_0 ( .a(n_29163), .b(n_25738), .c(FE_RN_1513_0), .d(FE_OCP_RBN3435_n_29163), .o(n_29271) );
in01f80 g745458 ( .a(n_34463), .o(n_34435) );
no02f80 g767307 ( .a(n_13549), .b(n_13548), .o(n_13550) );
in01f80 g751253 ( .a(n_29909), .o(n_29944) );
in01f80 newInst_379 ( .a(newNet_123), .o(newNet_379) );
in01f80 g738215 ( .a(n_41983), .o(n_41993) );
no02f80 g770338 ( .a(n_10720), .b(n_9875), .o(n_10718) );
no02f80 g767886 ( .a(n_13249), .b(n_13198), .o(n_13315) );
na02f80 g741063 ( .a(n_39048), .b(n_38996), .o(n_39134) );
oa22f80 g779265 ( .a(FE_OCP_RBN2173_n_1813), .b(n_1567), .c(n_1813), .d(n_1568), .o(n_1865) );
no02f80 g745641 ( .a(n_35477), .b(n_35463), .o(n_35931) );
in01f80 newInst_198 ( .a(newNet_115), .o(newNet_198) );
in01f80 g763706 ( .a(n_16712), .o(n_16713) );
na02f80 g777973 ( .a(n_3124), .b(n_3165), .o(n_3190) );
na02f80 g775492 ( .a(n_5770), .b(n_5581), .o(n_5793) );
in01f80 g763137 ( .a(n_17859), .o(n_17860) );
no02f80 g772675 ( .a(n_8480), .b(n_8479), .o(n_8481) );
no02f80 g767792 ( .a(n_12743), .b(delay_add_ln22_unr8_stage4_stallmux_q_22_), .o(n_12869) );
in01f80 newInst_1708 ( .a(newNet_1707), .o(newNet_1708) );
ao12f80 g739039 ( .a(n_40956), .b(n_41110), .c(n_40837), .o(n_41133) );
in01f80 newInst_3167 ( .a(newNet_3166), .o(newNet_3167) );
oa22f80 g779524 ( .a(n_1433), .b(n_607), .c(n_1403), .d(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n_2359) );
ao12f80 g754532 ( .a(n_26236), .b(n_26235), .c(n_26234), .o(n_26351) );
no02f80 g739288 ( .a(n_40770), .b(n_40769), .o(n_40934) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_29_ ( .ck(newNet_2537), .d(n_27784), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_) );
na02f80 g775761 ( .a(n_5304), .b(n_5251), .o(n_5409) );
no02f80 g766956 ( .a(n_14075), .b(n_14171), .o(n_14756) );
oa22f80 g739851 ( .a(n_40345), .b(n_39972), .c(n_40346), .d(n_39971), .o(n_40419) );
in01f80 FE_RC_3994_0 ( .a(FE_OCP_RBN1179_n_18981), .o(FE_RN_1732_0) );
in01f80 g737184 ( .a(n_42989), .o(n_43265) );
no02f80 g776927 ( .a(FE_OCP_RBN2646_n_47015), .b(n_3794), .o(n_3927) );
ao12f80 g774247 ( .a(n_6570), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .o(n_6660) );
in01f80 g764632 ( .a(n_16107), .o(n_16108) );
no02f80 g770995 ( .a(n_9798), .b(FE_OCP_RBN2558_n_44576), .o(n_9848) );
no02f80 g754178 ( .a(n_25943), .b(n_25970), .o(n_26098) );
in01f80 g737105 ( .a(FE_OCPN913_n_43022), .o(n_43120) );
na02f80 g752335 ( .a(n_27773), .b(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n_28098) );
na02f80 g748823 ( .a(n_32392), .b(n_32446), .o(n_32479) );
oa22f80 g752478 ( .a(n_27643), .b(n_24350), .c(n_27619), .d(n_27845), .o(n_27671) );
in01f80 fopt783798 ( .a(n_6214), .o(n_45479) );
in01f80 g739837 ( .a(n_40444), .o(n_40445) );
no02f80 g777869 ( .a(n_3133), .b(n_2450), .o(n_3141) );
ao22s80 g754609 ( .a(FE_OCP_RBN2960_n_26231), .b(n_25524), .c(FE_OCP_RBN3704_n_26231), .d(n_26419), .o(n_26937) );
in01f80 newInst_2213 ( .a(newNet_448), .o(newNet_2213) );
ao12f80 g782648 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32312), .c(n_32492), .o(n_44042) );
no02f80 g749918 ( .a(n_30172), .b(n_30171), .o(n_30200) );
oa22f80 FE_RC_87_0 ( .a(n_17192), .b(n_17072), .c(n_17020), .d(n_17073), .o(n_17340) );
in01f80 FE_RC_1674_0 ( .a(n_28310), .o(FE_RN_466_0) );
oa22f80 FE_RC_944_0 ( .a(n_20231), .b(n_22897), .c(n_22793), .d(n_22856), .o(n_22957) );
in01f80 FE_OCP_RBC2834_n_39586 ( .a(n_39586), .o(FE_OCP_RBN2834_n_39586) );
in01f80 newInst_1721 ( .a(newNet_1720), .o(newNet_1721) );
no02f80 g758306 ( .a(n_22288), .b(n_22331), .o(n_22438) );
na02f80 g741656 ( .a(FE_OCP_RBN2453_n_38537), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38576) );
no02f80 g765478 ( .a(n_15017), .b(n_15053), .o(n_15054) );
na02f80 g756765 ( .a(n_23472), .b(n_23512), .o(n_23537) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_17_ ( .ck(newNet_2399), .d(n_36415), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_) );
ao12f80 g754967 ( .a(n_25050), .b(n_25076), .c(n_25025), .o(n_25187) );
na02f80 g746791 ( .a(n_32911), .b(n_32916), .o(n_32947) );
in01f80 g743874 ( .a(n_36013), .o(n_36043) );
in01f80 g777408 ( .a(n_3450), .o(n_3485) );
in01f80 newInst_794 ( .a(newNet_793), .o(newNet_794) );
na02f80 g757722 ( .a(n_22623), .b(n_22529), .o(n_22740) );
no04s80 FE_RC_3309_0 ( .a(n_32599), .b(n_32600), .c(n_32601), .d(n_32602), .o(n_32617) );
no02f80 FE_RC_2243_0 ( .a(FE_RN_820_0), .b(FE_RN_821_0), .o(FE_RN_822_0) );
ao12f80 g774215 ( .a(n_6985), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .o(n_7034) );
in01f80 g771882 ( .a(n_8862), .o(n_8905) );
in01f80 g744959 ( .a(n_34999), .o(n_35897) );
na02f80 g752044 ( .a(n_28099), .b(n_28098), .o(n_28100) );
na02f80 g740163 ( .a(n_39812), .b(n_39548), .o(n_40013) );
in01f80 FE_RC_1925_0 ( .a(FE_RN_609_0), .o(n_35365) );
na02f80 g768038 ( .a(n_12914), .b(n_12965), .o(n_13115) );
in01f80 newInst_1660 ( .a(newNet_1659), .o(newNet_1660) );
no02f80 g772620 ( .a(n_8230), .b(n_8219), .o(n_8355) );
in01f80 newInst_2530 ( .a(newNet_2529), .o(newNet_2530) );
no02f80 g741328 ( .a(FE_OCP_RBN2546_n_44944), .b(n_38587), .o(n_39091) );
in01f80 FE_OCP_RBC3056_n_39913 ( .a(FE_OCP_RBN3053_n_39913), .o(FE_OCP_RBN3056_n_39913) );
no02f80 g740514 ( .a(n_39748), .b(n_39747), .o(n_39756) );
na04m80 FE_RC_1100_0 ( .a(n_37270), .b(n_37271), .c(n_37112), .d(n_37252), .o(n_37277) );
in01f80 g741167 ( .a(n_39244), .o(n_39245) );
no02f80 g763954 ( .a(n_16540), .b(n_17054), .o(n_17713) );
no02f80 g746880 ( .a(FE_OCP_RBN3387_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_28_), .o(n_33855) );
no02f80 g738569 ( .a(n_41533), .b(n_41571), .o(n_41572) );
na02f80 g778661 ( .a(n_2240), .b(n_2239), .o(n_2241) );
in01f80 g756130 ( .a(n_25026), .o(n_25188) );
in01f80 FE_OCP_RBC2216_FE_OCPN950_n_28595 ( .a(FE_OCP_RBN2214_FE_OCPN950_n_28595), .o(FE_OCP_RBN2216_FE_OCPN950_n_28595) );
in01f80 newInst_2379 ( .a(newNet_2378), .o(newNet_2379) );
na02f80 g757023 ( .a(n_23803), .b(n_23860), .o(n_24044) );
ao12f80 g774228 ( .a(n_6747), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .o(n_6852) );
no02f80 g760972 ( .a(n_19355), .b(n_19354), .o(n_19382) );
na02f80 g770909 ( .a(n_10129), .b(n_10070), .o(n_10169) );
na02f80 g749907 ( .a(n_30245), .b(n_30216), .o(n_30246) );
ao12f80 g738939 ( .a(n_41227), .b(n_41226), .c(n_41225), .o(n_41631) );
oa12f80 g777641 ( .a(n_3491), .b(n_3490), .c(n_3489), .o(n_5067) );
ao22s80 FE_RC_1346_0 ( .a(n_43544), .b(n_43826), .c(n_43543), .d(n_43825), .o(n_43863) );
no02f80 g774604 ( .a(n_6374), .b(n_6223), .o(n_6418) );
in01f80 FE_RC_3149_0 ( .a(n_20904), .o(FE_RN_1397_0) );
na02f80 g743595 ( .a(n_36400), .b(n_36045), .o(n_36447) );
na02f80 g761014 ( .a(n_19213), .b(n_19076), .o(n_19217) );
na02f80 g746798 ( .a(n_32915), .b(n_32912), .o(n_32946) );
in01f80 newInst_3103 ( .a(newNet_658), .o(newNet_3103) );
in01f80 newInst_58 ( .a(newNet_57), .o(newNet_58) );
in01f80 newInst_3601 ( .a(newNet_3600), .o(newNet_3601) );
no02f80 g766753 ( .a(n_14011), .b(n_14010), .o(n_14012) );
in01f80 newInst_1159 ( .a(newNet_1158), .o(newNet_1159) );
in01f80 newInst_622 ( .a(newNet_621), .o(newNet_622) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_22_ ( .ck(newNet_2748), .d(n_17550), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_) );
in01f80 g774161 ( .a(n_6669), .o(n_6948) );
in01f80 g754453 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_), .o(n_27050) );
in01f80 newInst_662 ( .a(newNet_661), .o(newNet_662) );
in01f80 newInst_3174 ( .a(newNet_1234), .o(newNet_3174) );
in01f80 g780234 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .o(n_1126) );
na02f80 g747299 ( .a(n_32690), .b(n_32855), .o(n_32853) );
in01f80 g780024 ( .a(n_1262), .o(n_1263) );
ao12f80 g755679 ( .a(n_24321), .b(n_24347), .c(n_21975), .o(n_24473) );
na02f80 g739863 ( .a(n_40265), .b(n_40046), .o(n_40263) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_6_ ( .ck(newNet_1899), .d(n_36874), .o(delay_sub_ln22_unr24_stage9_stallmux_q_6_) );
na02f80 g780822 ( .a(n_488), .b(n_464), .o(n_491) );
na02f80 g754746 ( .a(FE_OCP_RBN2959_n_26231), .b(n_25882), .o(n_26741) );
na02f80 g747412 ( .a(n_32687), .b(n_32632), .o(n_32649) );
in01f80 g772692 ( .a(n_8243), .o(n_8244) );
in01f80 g777937 ( .a(n_3167), .o(n_3168) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_8_ ( .ck(newNet_1564), .d(n_27001), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_) );
na02f80 g767031 ( .a(n_14758), .b(n_13649), .o(n_14296) );
no02f80 g739173 ( .a(n_40747), .b(FE_OCP_RBN2161_n_40687), .o(n_40896) );
oa12f80 g778181 ( .a(n_2175), .b(n_2645), .c(n_2149), .o(n_2805) );
no02f80 g745721 ( .a(n_44104), .b(n_34306), .o(n_34366) );
in01f80 FE_OCP_RBC2953_n_21538 ( .a(n_21538), .o(FE_OCP_RBN2953_n_21538) );
na02f80 g762137 ( .a(n_18703), .b(n_18667), .o(n_18668) );
in01f80 newInst_2647 ( .a(newNet_554), .o(newNet_2647) );
no02f80 g766762 ( .a(n_13722), .b(n_13721), .o(n_13805) );
na02f80 FE_RC_1732_0 ( .a(n_17864), .b(FE_RN_481_0), .o(n_17997) );
ao22s80 g757178 ( .a(n_23489), .b(n_23152), .c(n_23488), .d(n_23153), .o(n_23802) );
no02f80 g740076 ( .a(n_40110), .b(n_40112), .o(n_40137) );
na03f80 FE_RC_9_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .b(n_1551), .c(n_1393), .o(n_47027) );
na02f80 g760908 ( .a(n_20118), .b(n_20117), .o(n_20119) );
in01f80 g771709 ( .a(n_9387), .o(n_9388) );
na02f80 g744485 ( .a(n_35423), .b(n_35359), .o(n_35447) );
oa22f80 FE_RC_1376_0 ( .a(FE_OCPN1488_n_23447), .b(FE_OCP_RBN2852_n_26169), .c(n_23466), .d(n_26169), .o(n_26322) );
no02f80 g778668 ( .a(FE_OCP_RBN2290_n_2438), .b(n_2515), .o(n_2592) );
na02f80 g752289 ( .a(FE_OCP_RBN2179_FE_RN_526_0), .b(n_28498), .o(n_28499) );
in01f80 newInst_3222 ( .a(newNet_169), .o(newNet_3222) );
no02f80 g740602 ( .a(n_39559), .b(n_45840), .o(n_39579) );
na02f80 g738222 ( .a(n_41946), .b(n_41933), .o(n_41934) );
in01f80 FE_OCP_RBC1195_n_22542 ( .a(FE_OCP_RBN1193_n_22542), .o(FE_OCP_RBN1195_n_22542) );
in01f80 g751385 ( .a(n_28745), .o(n_28726) );
na02f80 g745592 ( .a(n_34286), .b(n_33540), .o(n_34460) );
na02f80 g742048 ( .a(FE_OCP_RBN2256_n_37844), .b(n_37587), .o(n_37984) );
na02f80 g764962 ( .a(n_16350), .b(n_16349), .o(n_16351) );
no02f80 g756539 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n_23735) );
in01f80 g759322 ( .a(n_21072), .o(n_21073) );
in01f80 g767066 ( .a(n_13793), .o(n_13794) );
no02f80 g748586 ( .a(n_31584), .b(n_31583), .o(n_31648) );
in01f80 FE_OCPC859_n_12880 ( .a(n_12739), .o(FE_OCPN859_n_12880) );
in01f80 FE_OCP_RBC1212_n_32142 ( .a(n_32142), .o(FE_OCP_RBN1212_n_32142) );
in01f80 g742572 ( .a(n_37535), .o(n_37534) );
ao12f80 g776666 ( .a(n_3970), .b(n_4213), .c(n_4035), .o(n_4305) );
no02f80 g740081 ( .a(n_39998), .b(n_39940), .o(n_40039) );
in01f80 FE_OCP_RBC1145_n_13098 ( .a(n_13098), .o(FE_OCP_RBN1145_n_13098) );
na02f80 g762887 ( .a(n_17523), .b(n_17282), .o(n_17659) );
oa12f80 g780851 ( .a(n_489), .b(n_521), .c(n_485), .o(n_637) );
oa12f80 g750347 ( .a(n_29592), .b(n_29666), .c(n_29632), .o(n_29674) );
in01f80 fopt783802 ( .a(n_5192), .o(n_45484) );
in01f80 g780727 ( .a(n_616), .o(n_617) );
no02f80 g758879 ( .a(n_21399), .b(FE_OCP_RBN1380_n_21240), .o(n_21442) );
na02f80 g773638 ( .a(n_7300), .b(n_7326), .o(n_7330) );
no02f80 FE_RC_1166_0 ( .a(FE_RN_351_0), .b(FE_RN_352_0), .o(FE_RN_353_0) );
oa22f80 g744584 ( .a(n_36598), .b(n_36052), .c(n_36619), .d(n_36053), .o(n_36680) );
na02f80 g758063 ( .a(n_22879), .b(n_22810), .o(n_23565) );
oa12f80 g746758 ( .a(FE_OCP_RBN3384_n_33108), .b(n_33253), .c(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n_33217) );
na02f80 g736932 ( .a(FE_OCPN910_n_43022), .b(n_46944), .o(n_43062) );
no02f80 g760780 ( .a(n_19653), .b(n_19685), .o(n_19686) );
oa12f80 g757889 ( .a(n_22065), .b(n_22113), .c(n_22035), .o(n_22237) );
no02f80 g749080 ( .a(n_30979), .b(n_29556), .o(n_31094) );
in01f80 g771633 ( .a(n_9017), .o(n_9018) );
no02f80 g778100 ( .a(n_2958), .b(FE_OCP_RBN3490_n_3390), .o(n_3003) );
na02f80 g773592 ( .a(n_7363), .b(n_7251), .o(n_7373) );
no02f80 g748126 ( .a(n_31905), .b(n_31819), .o(n_31968) );
no02f80 g770956 ( .a(n_9891), .b(FE_OCP_RBN3635_n_47260), .o(n_10047) );
in01f80 g743955 ( .a(n_35787), .o(n_35788) );
in01f80 g760022 ( .a(n_21691), .o(n_21714) );
in01f80 g777566 ( .a(n_4046), .o(n_4182) );
ao12f80 g743073 ( .a(n_37088), .b(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n_37345) );
oa22f80 FE_RC_3299_0 ( .a(n_17792), .b(n_17884), .c(n_17793), .d(n_17842), .o(n_17942) );
in01f80 newInst_648 ( .a(newNet_57), .o(newNet_648) );
in01f80 g740668 ( .a(n_39617), .o(n_39625) );
in01f80 g771386 ( .a(n_9266), .o(n_9267) );
in01f80 g770376 ( .a(n_10511), .o(n_10512) );
no02f80 g748940 ( .a(n_31013), .b(FE_OCP_DRV_N1588_n_31012), .o(n_31086) );
na02f80 g759649 ( .a(n_21799), .b(n_21798), .o(n_21800) );
in01f80 g748175 ( .a(n_32130), .o(n_32131) );
in01f80 g738970 ( .a(n_41190), .o(n_41484) );
na02f80 g737246 ( .a(n_42916), .b(n_42817), .o(n_42932) );
in01f80 FE_OCP_RBC2787_n_15079 ( .a(n_15079), .o(FE_OCP_RBN2787_n_15079) );
no02f80 g745876 ( .a(n_34134), .b(n_34110), .o(n_34189) );
na02f80 g759599 ( .a(n_20757), .b(n_20793), .o(n_20843) );
in01f80 FE_OCP_RBC2673_n_14991 ( .a(n_14991), .o(FE_OCP_RBN2673_n_14991) );
in01f80 g738503 ( .a(n_41638), .o(n_41587) );
in01f80 g771453 ( .a(n_9113), .o(n_9050) );
no02f80 g751375 ( .a(n_28705), .b(n_28649), .o(n_28727) );
in01f80 g743351 ( .a(n_36706), .o(n_36707) );
no02f80 g739703 ( .a(n_40501), .b(n_40374), .o(n_40521) );
no02f80 g749923 ( .a(n_30262), .b(n_30261), .o(n_30281) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_2_ ( .ck(newNet_1704), .d(n_21929), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_) );
na02f80 g740368 ( .a(n_39793), .b(n_39084), .o(n_39857) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_27_ ( .ck(newNet_3032), .d(n_1217), .o(delay_add_ln22_unr2_stage2_stallmux_q_27_) );
in01f80 g765285 ( .a(n_15926), .o(n_15927) );
na02f80 g781035 ( .a(sin_out_25), .b(FE_OFN4_n_43918), .o(n_331) );
na02f80 g764730 ( .a(n_15795), .b(FE_RN_473_0), .o(n_15850) );
in01f80 newInst_618 ( .a(newNet_510), .o(newNet_618) );
in01f80 g774134 ( .a(n_6739), .o(n_6700) );
oa12f80 g766404 ( .a(n_14622), .b(n_14621), .c(n_14620), .o(n_15718) );
na02f80 g754022 ( .a(n_26087), .b(FE_OCPN1440_n_23339), .o(n_26216) );
na02f80 g764439 ( .a(n_16159), .b(n_16157), .o(n_16277) );
in01f80 g748097 ( .a(n_32900), .o(n_32901) );
in01f80 FE_RC_2039_0 ( .a(n_25909), .o(FE_RN_682_0) );
na02f80 g784082 ( .a(n_8199), .b(n_45824), .o(n_45828) );
no02f80 g766186 ( .a(n_14544), .b(n_14543), .o(n_14572) );
na02f80 g760159 ( .a(n_20428), .b(n_20528), .o(n_20674) );
na02f80 g745305 ( .a(n_36118), .b(FE_OCP_RBN2987_n_35539), .o(n_36083) );
na02f80 g749933 ( .a(n_31065), .b(n_31041), .o(n_31042) );
oa22f80 g754801 ( .a(n_26006), .b(n_25710), .c(n_26005), .d(n_25711), .o(n_26680) );
in01f80 g753356 ( .a(n_27103), .o(n_27120) );
no02f80 g751752 ( .a(n_28309), .b(n_28308), .o(n_28310) );
no02f80 g751551 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_20_), .o(n_28550) );
in01f80 FE_OCPC1021_n_23195 ( .a(n_23195), .o(FE_OCPN1021_n_23195) );
in01f80 newInst_3137 ( .a(newNet_343), .o(newNet_3137) );
in01f80 FE_OCP_DRV_C1575_n_28829 ( .a(n_28829), .o(FE_OCP_DRV_N1575_n_28829) );
no02f80 g769189 ( .a(n_12083), .b(n_12014), .o(n_12610) );
in01f80 g747960 ( .a(n_31959), .o(n_32003) );
in01f80 newInst_1263 ( .a(newNet_1262), .o(newNet_1263) );
na02f80 g762366 ( .a(FE_OFN751_n_45003), .b(n_18492), .o(n_18839) );
in01f80 FE_OCP_RBC2581_n_3734 ( .a(n_3734), .o(FE_OCP_RBN2581_n_3734) );
in01f80 g776276 ( .a(n_4652), .o(n_4653) );
in01f80 newInst_2733 ( .a(newNet_2194), .o(newNet_2733) );
in01f80 newInst_2722 ( .a(newNet_1384), .o(newNet_2722) );
in01f80 FE_OCP_RBC3118_n_22755 ( .a(n_22755), .o(FE_OCP_RBN3118_n_22755) );
in01f80 newInst_1410 ( .a(newNet_1409), .o(newNet_1410) );
in01f80 newInst_2007 ( .a(newNet_2006), .o(newNet_2007) );
no02f80 g745649 ( .a(n_35453), .b(n_34842), .o(n_35463) );
oa12f80 g780191 ( .a(n_703), .b(n_837), .c(n_730), .o(n_1075) );
in01f80 newInst_2272 ( .a(newNet_1397), .o(newNet_2272) );
no02f80 g768696 ( .a(n_12108), .b(n_12071), .o(n_12072) );
in01f80 g770087 ( .a(n_10732), .o(n_10765) );
in01f80 FE_RC_2966_0 ( .a(FE_RN_1296_0), .o(n_11159) );
in01f80 FE_OCP_RBC2397_n_38586 ( .a(n_38586), .o(FE_OCP_RBN2397_n_38586) );
in01f80 newInst_3738 ( .a(newNet_1376), .o(newNet_3738) );
no02f80 g768596 ( .a(n_12261), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .o(n_12275) );
na02f80 g768083 ( .a(FE_OCPN860_n_12880), .b(n_13074), .o(n_13103) );
no02f80 g770421 ( .a(n_10607), .b(FE_OCP_RBN2568_n_8904), .o(n_10678) );
ao22s80 g768300 ( .a(n_44425), .b(n_12408), .c(n_44426), .d(n_12409), .o(n_13646) );
in01f80 g774150 ( .a(n_7168), .o(n_7169) );
no02f80 g754101 ( .a(n_26045), .b(FE_OCPN1494_n_23398), .o(n_26096) );
in01f80 newInst_1327 ( .a(newNet_58), .o(newNet_1327) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_6_ ( .ck(newNet_2997), .d(n_886), .o(delay_add_ln22_unr2_stage2_stallmux_q_6_) );
no02f80 g767560 ( .a(n_13051), .b(n_12284), .o(n_13224) );
in01f80 FE_RC_2242_0 ( .a(n_37253), .o(FE_RN_821_0) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_10_ ( .ck(newNet_986), .d(n_22894), .o(delay_xor_ln21_unr15_stage6_stallmux_q_10_) );
in01f80 FE_RC_3452_0 ( .a(n_26555), .o(FE_RN_1484_0) );
in01f80 FE_OCP_RBC2896_n_39575 ( .a(FE_OCP_RBN2895_n_39575), .o(FE_OCP_RBN2896_n_39575) );
in01f80 g780069 ( .a(n_1228), .o(n_1229) );
no02f80 g774341 ( .a(FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_5_), .o(n_6523) );
no02f80 g762460 ( .a(n_18327), .b(n_18326), .o(n_18328) );
na02f80 g769915 ( .a(n_10879), .b(n_44511), .o(n_10938) );
ms00f80 delay_sub_ln23_0_unr30_stage10_stallmux_q_reg ( .ck(newNet_1272), .d(n_45898), .o(delay_sub_ln23_0_unr30_stage10_stallmux_q) );
in01f80 g764116 ( .a(n_16624), .o(n_16625) );
in01f80 FE_RC_1118_0 ( .a(n_3127), .o(FE_RN_336_0) );
in01f80 newInst_1712 ( .a(newNet_1711), .o(newNet_1712) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_11_ ( .ck(newNet_1770), .d(n_22116), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_) );
na02f80 FE_RC_3071_0 ( .a(n_26319), .b(FE_RN_1350_0), .o(FE_RN_1351_0) );
in01f80 newInst_2431 ( .a(newNet_2430), .o(newNet_2431) );
na02f80 g750397 ( .a(n_30634), .b(n_30616), .o(n_30617) );
in01f80 g745807 ( .a(n_34128), .o(n_34116) );
in01f80 g737404 ( .a(n_42806), .o(n_42807) );
no02f80 FE_RC_3062_0 ( .a(FE_OCP_RBN1349_n_19270), .b(FE_RN_1343_0), .o(FE_RN_1344_0) );
no02f80 g763765 ( .a(n_16751), .b(n_16715), .o(n_16752) );
na02f80 g777250 ( .a(n_3504), .b(n_3518), .o(n_3616) );
ao12f80 g767588 ( .a(n_12555), .b(n_12802), .c(n_12583), .o(n_12875) );
in01f80 g742484 ( .a(n_37702), .o(n_37703) );
no02f80 g760468 ( .a(n_20005), .b(n_20029), .o(n_20046) );
oa22f80 FE_RC_31_0 ( .a(FE_OFN84_n_46137), .b(n_6519), .c(FE_OFN806_n_46196), .d(n_6529), .o(n_46184) );
in01f80 g776677 ( .a(n_3896), .o(n_3905) );
oa12f80 g755152 ( .a(n_25571), .b(n_25714), .c(n_25604), .o(n_25773) );
ao12f80 g781006 ( .a(n_52), .b(n_272), .c(n_103), .o(n_276) );
no02f80 g780620 ( .a(n_890), .b(n_905), .o(n_985) );
no02f80 g765832 ( .a(FE_OCP_RBN1185_n_14823), .b(FE_OCP_RBN2503_n_13896), .o(n_14888) );
ao22s80 g736502 ( .a(n_43696), .b(n_43590), .c(n_43697), .d(n_43589), .o(n_43724) );
no02f80 g778758 ( .a(n_2354), .b(n_2353), .o(n_2355) );
no02f80 g760865 ( .a(n_19334), .b(n_18539), .o(n_19391) );
in01f80 g737971 ( .a(n_42202), .o(n_42277) );
na02f80 g766201 ( .a(n_14414), .b(n_14377), .o(n_14556) );
oa22f80 FE_RC_889_0 ( .a(n_20633), .b(n_20926), .c(n_20632), .d(n_20861), .o(n_20984) );
na02f80 g769730 ( .a(n_11239), .b(n_11043), .o(n_11291) );
in01f80 g760595 ( .a(n_19961), .o(n_19962) );
no02f80 g757497 ( .a(n_22899), .b(n_22898), .o(n_22987) );
na02f80 g738861 ( .a(n_41310), .b(n_41309), .o(n_41322) );
in01f80 g780388 ( .a(n_950), .o(n_864) );
in01f80 fopt784300 ( .a(beta_31), .o(n_7) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_7_ ( .ck(newNet_484), .d(n_22777), .o(delay_xor_ln22_unr15_stage6_stallmux_q_7_) );
in01f80 g742996 ( .a(n_37012), .o(n_36963) );
na02f80 g777365 ( .a(n_5494), .b(n_4693), .o(n_4833) );
no02f80 g757983 ( .a(n_22048), .b(FE_OCP_RBN1337_n_20941), .o(n_22082) );
na02f80 g757601 ( .a(n_22795), .b(n_44061), .o(n_22816) );
in01f80 FE_OCP_DRV_C1605_n_31445 ( .a(n_31445), .o(FE_OCP_DRV_N1605_n_31445) );
in01f80 g779224 ( .a(n_1938), .o(n_1939) );
no02f80 g764360 ( .a(n_16234), .b(n_16233), .o(n_16235) );
no02f80 g743404 ( .a(n_36570), .b(n_36587), .o(n_36655) );
no02f80 g737430 ( .a(n_42690), .b(n_42707), .o(n_42780) );
oa22f80 FE_RC_962_0 ( .a(n_32124), .b(n_32365), .c(n_32125), .d(n_32364), .o(n_32519) );
in01f80 g773343 ( .a(FE_OCP_RBN3475_n_7886), .o(n_8189) );
in01f80 g765026 ( .a(n_15286), .o(n_15316) );
in01f80 newInst_1314 ( .a(newNet_1313), .o(newNet_1314) );
no02f80 g777876 ( .a(n_3241), .b(n_3161), .o(n_3242) );
in01f80 newInst_528 ( .a(newNet_527), .o(newNet_528) );
in01f80 g779362 ( .a(n_1616), .o(n_1617) );
na02f80 FE_RC_1162_0 ( .a(FE_RN_350_0), .b(n_41598), .o(n_41727) );
na02f80 g737889 ( .a(n_42201), .b(n_42323), .o(n_42416) );
na02f80 g777341 ( .a(n_4759), .b(FE_OFN822_n_4597), .o(n_4852) );
oa12f80 g767321 ( .a(n_13039), .b(n_13638), .c(n_13312), .o(n_13680) );
no02f80 g740265 ( .a(n_40133), .b(n_40132), .o(n_40173) );
in01f80 g765861 ( .a(n_14979), .o(n_14950) );
no02f80 g752964 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n_28200) );
na02f80 g777127 ( .a(n_3784), .b(FE_OCPN966_n_47020), .o(n_3928) );
no02f80 g776426 ( .a(FE_OCP_RBN2698_n_4238), .b(n_3106), .o(n_4381) );
no02f80 g746762 ( .a(n_33103), .b(n_33108), .o(n_33203) );
no02f80 g761195 ( .a(n_19187), .b(n_19186), .o(n_19188) );
oa12f80 g744714 ( .a(n_35121), .b(n_35107), .c(n_35106), .o(n_35210) );
oa22f80 FE_RC_913_0 ( .a(n_25318), .b(FE_OCP_RBN1060_n_24473), .c(n_24204), .d(n_24473), .o(n_24576) );
no02f80 g761340 ( .a(n_20084), .b(n_20112), .o(n_20599) );
ao12f80 g761644 ( .a(n_19490), .b(n_19489), .c(n_19488), .o(n_19928) );
in01f80 g759900 ( .a(n_21478), .o(n_21479) );
in01f80 FE_RC_2420_0 ( .a(n_6767), .o(FE_RN_957_0) );
in01f80 g745685 ( .a(n_34297), .o(n_34286) );
na02f80 g750272 ( .a(n_30838), .b(n_30837), .o(n_30839) );
no02f80 g753937 ( .a(n_26182), .b(n_26207), .o(n_26286) );
oa12f80 g781102 ( .a(n_238), .b(n_244), .c(n_237), .o(n_447) );
ao12f80 g763621 ( .a(n_17663), .b(n_17732), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .o(n_18385) );
no02f80 g750144 ( .a(n_30925), .b(n_30902), .o(n_30903) );
in01f80 newInst_1801 ( .a(newNet_1800), .o(newNet_1801) );
in01f80 newInst_971 ( .a(newNet_970), .o(newNet_971) );
in01f80 g776519 ( .a(FE_OCP_RBN2700_n_4238), .o(n_5422) );
no02f80 g771832 ( .a(n_9517), .b(n_9596), .o(n_9961) );
na02f80 g762218 ( .a(n_18663), .b(n_18586), .o(n_18739) );
in01f80 g766061 ( .a(n_14801), .o(n_14711) );
no02f80 g753570 ( .a(n_26673), .b(n_26699), .o(n_26804) );
oa12f80 g739272 ( .a(n_40877), .b(n_40876), .c(n_40875), .o(n_40929) );
oa12f80 g754599 ( .a(n_25462), .b(n_25461), .c(n_25460), .o(n_27040) );
na02f80 g759608 ( .a(n_20648), .b(n_20618), .o(n_20820) );
ao22s80 FE_RC_3821_0 ( .a(FE_OCPN1858_n_22207), .b(n_24797), .c(n_24828), .d(n_24918), .o(n_24967) );
oa12f80 g780767 ( .a(n_530), .b(n_558), .c(n_542), .o(n_565) );
na02f80 g778581 ( .a(n_2303), .b(n_1965), .o(n_2369) );
in01f80 g756181 ( .a(n_24245), .o(n_24332) );
no02f80 g749189 ( .a(n_30771), .b(n_27130), .o(n_30858) );
no02f80 g784131 ( .a(n_7136), .b(n_7135), .o(n_45878) );
in01f80 g763014 ( .a(n_17739), .o(n_17740) );
in01f80 newInst_2472 ( .a(newNet_242), .o(newNet_2472) );
na02f80 g765572 ( .a(n_15103), .b(FE_OCPN3767_n_14439), .o(n_15328) );
no02f80 g744672 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_36556) );
no02f80 g743032 ( .a(n_37100), .b(n_37111), .o(n_37153) );
oa12f80 g746323 ( .a(n_33526), .b(n_33525), .c(n_33524), .o(n_33583) );
in01f80 FE_RC_3083_0 ( .a(n_20429), .o(FE_RN_1360_0) );
in01f80 FE_RC_3612_0 ( .a(n_27014), .o(FE_RN_1580_0) );
na02f80 g758298 ( .a(FE_OCPN991_n_22249), .b(n_21011), .o(n_22465) );
no02f80 g757445 ( .a(n_22868), .b(n_22940), .o(n_22995) );
no02f80 g756740 ( .a(n_23513), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .o(n_23542) );
ao12f80 g768274 ( .a(n_12643), .b(n_12644), .c(n_12642), .o(n_12716) );
na02f80 g754482 ( .a(n_26351), .b(FE_OCP_RBN2961_n_26231), .o(n_26816) );
in01f80 g768633 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_26_), .o(n_12215) );
no02f80 g744457 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_36774) );
no02f80 g766328 ( .a(n_14701), .b(n_14700), .o(n_14702) );
in01f80 g780576 ( .a(n_1191), .o(n_752) );
in01f80 newInst_1651 ( .a(newNet_561), .o(newNet_1651) );
in01f80 newInst_47 ( .a(newNet_46), .o(newNet_47) );
na02f80 g779420 ( .a(n_1746), .b(n_1723), .o(n_1747) );
ao22s80 g762632 ( .a(n_18232), .b(n_17704), .c(n_18231), .d(n_17705), .o(n_18526) );
in01f80 newInst_3085 ( .a(newNet_3084), .o(newNet_3085) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_23_ ( .ck(newNet_1399), .d(n_36714), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_) );
oa22f80 g752515 ( .a(n_27632), .b(n_27497), .c(FE_OCP_RBN3126_n_27632), .d(n_27496), .o(n_27728) );
in01f80 g751077 ( .a(n_28894), .o(n_28868) );
in01f80 FE_RC_2954_0 ( .a(n_44490), .o(FE_RN_1290_0) );
na02f80 g766318 ( .a(n_14358), .b(n_14376), .o(n_14438) );
no02f80 g743827 ( .a(n_36071), .b(n_47264), .o(n_36105) );
oa22f80 g753439 ( .a(n_27559), .b(n_26906), .c(n_27560), .d(n_26905), .o(n_27588) );
in01f80 FE_OCP_DRV_C3741_n_29576 ( .a(FE_OCP_DRV_N3740_n_29576), .o(FE_OCP_DRV_N3741_n_29576) );
in01f80 newInst_3653 ( .a(newNet_3652), .o(newNet_3653) );
in01f80 newInst_925 ( .a(newNet_924), .o(newNet_925) );
in01f80 g758653 ( .a(n_21816), .o(n_21817) );
in01f80 g752244 ( .a(n_28056), .o(n_28057) );
in01f80 g778991 ( .a(n_2197), .o(n_2198) );
na02f80 g759473 ( .a(n_20913), .b(n_20608), .o(n_20973) );
ao12f80 g757173 ( .a(n_23531), .b(n_23530), .c(n_23529), .o(n_23860) );
in01f80 FE_OCP_RBC2168_n_32892 ( .a(FE_OCP_RBN2166_n_32892), .o(FE_OCP_RBN2168_n_32892) );
no02f80 g752148 ( .a(n_28064), .b(n_44735), .o(n_28066) );
oa12f80 g755914 ( .a(n_25141), .b(n_25160), .c(n_24844), .o(n_25883) );
na02f80 g749613 ( .a(n_30327), .b(n_30326), .o(n_30328) );
in01f80 newInst_577 ( .a(newNet_576), .o(newNet_577) );
na02f80 g778632 ( .a(n_2613), .b(n_2736), .o(n_3156) );
no02f80 g758179 ( .a(n_22435), .b(n_22292), .o(n_22501) );
in01f80 g780278 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .o(n_1031) );
in01f80 g766740 ( .a(n_13813), .o(n_13755) );
in01f80 g779502 ( .a(n_1485), .o(n_1486) );
no02f80 g778697 ( .a(n_2235), .b(n_1566), .o(n_2266) );
no03m80 FE_RC_1080_0 ( .a(FE_OCP_RBN3377_n_1675), .b(FE_RN_2_0), .c(n_1517), .o(n_1725) );
ao22s80 g784426 ( .a(n_36745), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .o(n_46238) );
oa12f80 g774525 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_6717) );
in01f80 FE_OCP_RBC3467_n_7886 ( .a(FE_OCP_RBN3462_n_7886), .o(FE_OCP_RBN3467_n_7886) );
oa22f80 FE_RC_1170_0 ( .a(n_11739), .b(n_11959), .c(n_11740), .d(n_11985), .o(n_12196) );
na02f80 g741130 ( .a(n_39326), .b(n_38976), .o(n_39360) );
na02f80 g740251 ( .a(n_40243), .b(n_40313), .o(n_40365) );
in01f80 g736773 ( .a(n_43055), .o(n_43056) );
in01f80 newInst_1096 ( .a(newNet_1095), .o(newNet_1096) );
in01f80 g767738 ( .a(n_12771), .o(n_12808) );
in01f80 g762700 ( .a(n_17944), .o(n_17945) );
na02f80 g762124 ( .a(n_18220), .b(n_18187), .o(n_18221) );
oa12f80 g757525 ( .a(n_22349), .b(n_22686), .c(n_22194), .o(n_22685) );
na02f80 g740916 ( .a(n_39257), .b(n_39299), .o(n_39340) );
in01f80 FE_OCP_RBC1179_n_18981 ( .a(FE_OCP_RBN1178_n_18981), .o(FE_OCP_RBN1179_n_18981) );
ao12f80 g746703 ( .a(n_34253), .b(n_34252), .c(n_34251), .o(n_34774) );
in01f80 FE_OCP_RBC3134_n_6567 ( .a(n_6567), .o(FE_OCP_RBN3134_n_6567) );
no02f80 g773070 ( .a(n_7839), .b(n_7858), .o(n_7859) );
na02f80 g758335 ( .a(n_22288), .b(n_21080), .o(n_22466) );
no02f80 g740060 ( .a(n_40118), .b(n_40011), .o(n_40012) );
in01f80 newInst_1957 ( .a(newNet_1956), .o(newNet_1957) );
no02f80 g776931 ( .a(n_3759), .b(n_3528), .o(n_3821) );
ao22s80 FE_RC_1574_0 ( .a(FE_OCP_RBN3313_delay_xor_ln22_unr18_stage7_stallmux_q_2_), .b(FE_OCP_RBN3308_n_44722), .c(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .d(n_44759), .o(n_27827) );
in01f80 FE_OCP_DRV_C1585_n_35594 ( .a(n_35594), .o(FE_OCP_DRV_N1585_n_35594) );
na02f80 g753152 ( .a(n_27380), .b(n_27329), .o(n_27486) );
ao12f80 g737614 ( .a(n_42298), .b(n_42311), .c(n_42202), .o(n_42373) );
na02f80 g762448 ( .a(n_18106), .b(delay_add_ln22_unr11_stage5_stallmux_q_14_), .o(n_18126) );
in01f80 g758103 ( .a(n_22261), .o(n_22262) );
in01f80 g751936 ( .a(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_34037) );
in01f80 newInst_2604 ( .a(newNet_2603), .o(newNet_2604) );
in01f80 FE_OCP_RBC1175_n_18981 ( .a(n_18981), .o(FE_OCP_RBN1175_n_18981) );
no02f80 g755432 ( .a(n_24687), .b(FE_OCPN1482_n_22207), .o(n_24808) );
no02f80 g748332 ( .a(n_31835), .b(n_30574), .o(n_31953) );
in01f80 newInst_2995 ( .a(newNet_2994), .o(newNet_2995) );
in01f80 g769868 ( .a(n_11134), .o(n_11164) );
no02f80 g768490 ( .a(FE_OCP_RBN3383_n_12365), .b(n_12043), .o(n_12423) );
no02f80 g780791 ( .a(n_528), .b(n_527), .o(n_529) );
na02f80 g752971 ( .a(n_27274), .b(n_27231), .o(n_27277) );
na02f80 g767761 ( .a(n_13025), .b(n_13024), .o(n_13099) );
no02f80 g777109 ( .a(n_3706), .b(n_3700), .o(n_3839) );
no02f80 g772285 ( .a(n_8576), .b(n_8545), .o(n_8666) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_18_ ( .ck(newNet_1240), .d(n_5929), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_) );
no02f80 g768590 ( .a(n_12232), .b(delay_add_ln22_unr8_stage4_stallmux_q_7_), .o(n_12262) );
in01f80 FE_OCP_RBC3384_n_33108 ( .a(n_33108), .o(FE_OCP_RBN3384_n_33108) );
in01f80 g771560 ( .a(n_10733), .o(n_9200) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_24_ ( .ck(newNet_1838), .d(n_16849), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_) );
ao22s80 FE_RC_1326_0 ( .a(n_20414), .b(n_20303), .c(n_20286), .d(n_20415), .o(n_20545) );
na02f80 g745186 ( .a(n_34594), .b(n_34763), .o(n_34818) );
in01f80 g775631 ( .a(n_5638), .o(n_5639) );
in01f80 newInst_754 ( .a(newNet_753), .o(newNet_754) );
na02f80 g765289 ( .a(n_16255), .b(n_16174), .o(n_16306) );
in01f80 newInst_519 ( .a(newNet_518), .o(newNet_519) );
in01f80 g763319 ( .a(n_17386), .o(n_17387) );
ao12f80 g775327 ( .a(n_5877), .b(n_5876), .c(n_5582), .o(n_5902) );
na02f80 g774321 ( .a(n_6580), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6801) );
in01f80 FE_OCP_DRV_C1611_n_21706 ( .a(n_21706), .o(FE_OCP_DRV_N1611_n_21706) );
no02f80 g774743 ( .a(n_6321), .b(n_6322), .o(n_6350) );
oa22f80 FE_RC_3875_0 ( .a(n_12961), .b(n_13816), .c(n_12962), .d(n_13815), .o(n_13927) );
no02f80 FE_RC_3858_0 ( .a(FE_RN_1683_0), .b(n_21046), .o(FE_RN_1684_0) );
oa12f80 g770192 ( .a(n_10842), .b(n_10869), .c(n_10841), .o(n_10913) );
no02f80 g776556 ( .a(n_4305), .b(n_4045), .o(n_4357) );
na02f80 g766385 ( .a(n_14125), .b(n_14062), .o(n_14158) );
in01f80 g739451 ( .a(n_40901), .o(n_40872) );
no02f80 FE_RC_2563_0 ( .a(FE_RN_1050_0), .b(FE_OCP_RBN1980_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_RN_1052_0) );
in01f80 g773663 ( .a(n_7358), .o(n_7343) );
no02f80 FE_RC_216_0 ( .a(FE_RN_71_0), .b(n_12478), .o(n_12523) );
oa12f80 g767246 ( .a(n_13588), .b(n_13626), .c(n_13625), .o(n_13639) );
in01f80 g778526 ( .a(n_2630), .o(n_2631) );
na02f80 g739119 ( .a(n_41014), .b(n_40865), .o(n_41048) );
na02f80 g769058 ( .a(FE_OCP_RBN3265_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(n_11650) );
no02f80 g762776 ( .a(n_17889), .b(n_17888), .o(n_17890) );
na02f80 g773667 ( .a(n_7238), .b(delay_add_ln22_unr5_stage3_stallmux_q_17_), .o(n_7300) );
no02f80 g738574 ( .a(n_41530), .b(n_41529), .o(n_41567) );
no02f80 g771970 ( .a(FE_OCPN955_n_44460), .b(n_9768), .o(n_9876) );
in01f80 newInst_702 ( .a(newNet_701), .o(newNet_702) );
in01f80 newInst_3560 ( .a(newNet_3559), .o(newNet_3560) );
na02f80 g771696 ( .a(n_8964), .b(FE_OCP_RBN2385_n_8342), .o(n_9027) );
na02f80 g743187 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_3_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .o(n_36897) );
in01f80 FE_OCP_RBC2508_n_13896 ( .a(FE_OCP_RBN2503_n_13896), .o(FE_OCP_RBN2508_n_13896) );
in01f80 g773865 ( .a(n_7053), .o(n_7054) );
in01f80 FE_RC_2260_0 ( .a(n_25032), .o(FE_RN_836_0) );
no02f80 g750952 ( .a(n_30039), .b(n_30038), .o(n_30040) );
in01f80 newInst_878 ( .a(newNet_877), .o(newNet_878) );
no02f80 g761140 ( .a(n_19063), .b(n_18391), .o(n_19115) );
in01f80 FE_RC_4099_0 ( .a(n_31518), .o(FE_RN_1793_0) );
oa12f80 g766813 ( .a(n_13942), .b(n_13943), .c(n_13941), .o(n_15482) );
in01f80 newInst_3226 ( .a(newNet_3225), .o(newNet_3226) );
oa12f80 g749748 ( .a(n_31121), .b(n_31120), .c(n_31119), .o(n_31417) );
no02f80 g756554 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23818) );
na02f80 g776187 ( .a(n_4891), .b(n_4890), .o(n_4892) );
no02f80 g747003 ( .a(n_32990), .b(n_32989), .o(n_33012) );
na02f80 g744489 ( .a(n_35428), .b(FE_OCP_DRV_N1540_n_35427), .o(n_35536) );
in01f80 g768985 ( .a(n_11900), .o(n_11901) );
in01f80 g741521 ( .a(n_38709), .o(n_38705) );
in01f80 g768283 ( .a(n_12558), .o(n_12559) );
in01f80 g744133 ( .a(n_36240), .o(n_36241) );
no02f80 g756750 ( .a(n_23514), .b(n_23498), .o(n_23499) );
in01f80 FE_OCP_RBC3048_n_6013 ( .a(n_6013), .o(FE_OCP_RBN3048_n_6013) );
in01f80 g737584 ( .a(n_42769), .o(n_42770) );
in01f80 newInst_2375 ( .a(newNet_759), .o(newNet_2375) );
na02f80 g773098 ( .a(n_7739), .b(n_7841), .o(n_8371) );
in01f80 FE_OFC756_n_44461 ( .a(FE_OCP_RBN2616_n_44561), .o(FE_RN_1433_0) );
na02f80 g749846 ( .a(n_31044), .b(n_31043), .o(n_31066) );
no02f80 g751447 ( .a(n_28736), .b(n_28723), .o(n_28724) );
in01f80 FE_RC_3426_0 ( .a(FE_RN_1482_0), .o(n_30708) );
in01f80 g762622 ( .a(n_18124), .o(n_18125) );
no02f80 g745005 ( .a(n_34796), .b(n_34831), .o(n_34905) );
no02f80 g739449 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .o(n_40769) );
oa22f80 g744973 ( .a(n_34878), .b(FE_OFN627_n_34445), .c(n_34879), .d(n_34446), .o(n_34978) );
oa22f80 g770666 ( .a(FE_OCP_RBN2822_n_10023), .b(FE_OCP_RBN3597_FE_OCPN1243_n_44460), .c(n_10023), .d(FE_RN_1433_0), .o(n_10192) );
no02f80 g778672 ( .a(FE_OCP_RBN2294_n_2438), .b(n_2611), .o(n_2660) );
no02f80 g759191 ( .a(n_21382), .b(n_21456), .o(n_21527) );
in01f80 g766433 ( .a(n_14125), .o(n_14126) );
oa12f80 g737958 ( .a(n_42183), .b(n_42182), .c(n_42181), .o(n_43025) );
in01f80 newInst_1783 ( .a(newNet_1782), .o(newNet_1783) );
no02f80 g751169 ( .a(n_29944), .b(n_29942), .o(n_29977) );
in01f80 FE_OCP_RBC2800_n_15706 ( .a(n_15706), .o(FE_OCP_RBN2800_n_15706) );
in01f80 g762675 ( .a(n_18251), .o(n_18252) );
no02f80 FE_RC_632_0 ( .a(FE_RN_195_0), .b(FE_RN_196_0), .o(FE_RN_197_0) );
na02f80 g738009 ( .a(n_42129), .b(n_42174), .o(n_42189) );
in01f80 g763009 ( .a(n_17622), .o(n_17623) );
na02f80 g738924 ( .a(n_41249), .b(n_41248), .o(n_41250) );
oa12f80 g737847 ( .a(n_42197), .b(n_42178), .c(n_42196), .o(n_42198) );
na02f80 g772696 ( .a(n_8259), .b(n_8268), .o(n_8368) );
ao12f80 g765380 ( .a(n_15874), .b(n_15958), .c(n_15957), .o(n_16016) );
na02f80 FE_RC_3901_0 ( .a(FE_RN_1693_0), .b(FE_RN_1694_0), .o(FE_RN_1695_0) );
no02f80 g775378 ( .a(n_5575), .b(n_5605), .o(n_5717) );
na02f80 g737033 ( .a(n_43030), .b(n_43083), .o(n_43529) );
in01f80 g773751 ( .a(n_8174), .o(n_7327) );
oa12f80 g773225 ( .a(n_7625), .b(n_7624), .c(n_7623), .o(n_8150) );
ao22s80 FE_RC_3221_0 ( .a(n_7591), .b(n_8788), .c(n_7590), .d(n_8769), .o(n_8915) );
in01f80 g747302 ( .a(n_32597), .o(n_32598) );
in01f80 g761732 ( .a(n_18681), .o(n_18714) );
na02f80 g744497 ( .a(n_35405), .b(n_35401), .o(n_35475) );
no02f80 g776489 ( .a(n_4407), .b(n_4140), .o(n_4470) );
oa12f80 g769241 ( .a(n_11570), .b(n_11707), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n_12198) );
no02f80 g763805 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .o(n_17310) );
ao22s80 g780855 ( .a(n_457), .b(n_375), .c(n_420), .d(n_501), .o(n_527) );
no02f80 g757221 ( .a(n_44995), .b(n_23184), .o(n_23569) );
na02f80 g756738 ( .a(n_23423), .b(n_22203), .o(n_23503) );
in01f80 g737351 ( .a(n_42839), .o(n_42840) );
no02f80 g775302 ( .a(n_5798), .b(n_5516), .o(n_5811) );
na02f80 g747083 ( .a(n_32762), .b(n_32792), .o(n_32862) );
na02f80 g778271 ( .a(n_2676), .b(n_3058), .o(n_2677) );
no02f80 g748971 ( .a(n_31097), .b(n_30988), .o(n_31133) );
no02f80 g770341 ( .a(n_10590), .b(n_10587), .o(n_10647) );
no02f80 g759163 ( .a(n_21018), .b(n_20754), .o(n_21093) );
in01f80 newInst_997 ( .a(newNet_968), .o(newNet_997) );
no02f80 g780416 ( .a(n_846), .b(n_845), .o(n_955) );
no02f80 g774477 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n_6850) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_25_ ( .ck(newNet_3037), .d(n_1206), .o(delay_add_ln22_unr2_stage2_stallmux_q_25_) );
in01f80 g772589 ( .a(n_8369), .o(n_8433) );
in01f80 g769748 ( .a(n_11297), .o(n_11265) );
no02f80 g751736 ( .a(n_28319), .b(n_28091), .o(n_28331) );
no02f80 g777271 ( .a(n_3629), .b(n_3571), .o(n_3670) );
in01f80 g739177 ( .a(n_40897), .o(n_40833) );
no02f80 g736756 ( .a(n_43202), .b(n_43204), .o(n_43222) );
in01f80 FE_RC_970_0 ( .a(n_26158), .o(FE_RN_279_0) );
na02f80 g780502 ( .a(n_733), .b(n_753), .o(n_1012) );
na02f80 g779302 ( .a(n_1730), .b(n_1729), .o(n_1846) );
no02f80 g776608 ( .a(n_4315), .b(n_4259), .o(n_4479) );
na02f80 g755144 ( .a(n_25074), .b(n_25073), .o(n_25075) );
na02f80 g765333 ( .a(FE_OCP_RBN3621_n_15135), .b(n_14157), .o(n_15486) );
na02f80 g762420 ( .a(n_45002), .b(n_18688), .o(n_18810) );
ao12f80 g746421 ( .a(n_33457), .b(n_33456), .c(n_33455), .o(n_34123) );
in01f80 newInst_3067 ( .a(newNet_3066), .o(newNet_3067) );
no02f80 g759244 ( .a(n_20975), .b(n_20942), .o(n_21094) );
no02f80 g741302 ( .a(n_38830), .b(n_38146), .o(n_38853) );
no02f80 g759716 ( .a(n_20542), .b(n_45066), .o(n_20682) );
in01f80 g772259 ( .a(n_8812), .o(n_8831) );
no02f80 g780442 ( .a(n_855), .b(n_46055), .o(n_788) );
no02f80 g784069 ( .a(n_802), .b(n_45812), .o(n_45815) );
in01f80 FE_OCP_RBC2595_n_25181 ( .a(FE_OCP_RBN2592_n_25181), .o(FE_OCP_RBN2595_n_25181) );
na02f80 g740397 ( .a(n_39787), .b(n_39910), .o(n_39994) );
in01f80 g758067 ( .a(n_22761), .o(n_22762) );
in01f80 FE_OCPC1464_n_29630 ( .a(FE_OCPN1463_n_29630), .o(FE_OCPN1464_n_29630) );
oa12f80 g743687 ( .a(n_36188), .b(n_36279), .c(n_35619), .o(n_36347) );
in01f80 FE_RC_3548_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .o(FE_RN_1538_0) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_12_ ( .ck(newNet_2975), .d(n_5724), .o(delay_add_ln22_unr5_stage3_stallmux_q_12_) );
no02f80 g763414 ( .a(n_16839), .b(n_17118), .o(n_17213) );
no02f80 g763398 ( .a(n_16919), .b(n_16191), .o(n_16996) );
in01f80 g771058 ( .a(n_9461), .o(n_9465) );
no02f80 g743302 ( .a(n_36736), .b(n_36755), .o(n_36767) );
no02f80 g754758 ( .a(n_25366), .b(n_25333), .o(n_25334) );
na02f80 g759518 ( .a(n_20850), .b(n_20495), .o(n_20851) );
in01f80 newInst_1922 ( .a(newNet_1921), .o(newNet_1922) );
in01f80 g781161 ( .a(n_199), .o(n_194) );
in01f80 g739081 ( .a(n_41126), .o(n_41415) );
in01f80 FE_OCPC908_n_23227 ( .a(FE_OCPN907_n_23227), .o(FE_OCPN908_n_23227) );
no02f80 g748811 ( .a(n_32603), .b(n_32486), .o(n_32823) );
in01f80 g773791 ( .a(n_7204), .o(n_7205) );
oa22f80 g740228 ( .a(n_39788), .b(n_39804), .c(n_39789), .d(n_39805), .o(n_39896) );
oa12f80 g756091 ( .a(n_24100), .b(n_24161), .c(n_21852), .o(n_24207) );
ao22s80 g740817 ( .a(n_39468), .b(n_39423), .c(n_39381), .d(n_39424), .o(n_39947) );
in01f80 g770571 ( .a(n_10195), .o(n_10196) );
oa12f80 g738931 ( .a(n_41170), .b(n_41169), .c(n_41168), .o(n_41613) );
oa22f80 g751278 ( .a(n_28708), .b(n_28463), .c(n_28748), .d(n_28464), .o(n_29844) );
na02f80 g762108 ( .a(n_18246), .b(n_18222), .o(n_18261) );
oa22f80 g744878 ( .a(n_46953), .b(n_36210), .c(n_36402), .d(n_36209), .o(n_36452) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_18_ ( .ck(newNet_2107), .d(n_46995), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_) );
in01f80 g777236 ( .a(n_3650), .o(n_3686) );
in01f80 g757541 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_31_), .o(n_22929) );
oa12f80 g749488 ( .a(n_31350), .b(n_31782), .c(n_31286), .o(n_31888) );
in01f80 FE_RC_2744_0 ( .a(n_12432), .o(FE_RN_1165_0) );
oa12f80 g762710 ( .a(n_17155), .b(n_18210), .c(n_17309), .o(n_18231) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_30_ ( .ck(newNet_3115), .d(FE_OCP_RBN3108_n_40586), .o(delay_add_ln22_unr27_stage10_stallmux_q_30_) );
oa22f80 g784353 ( .a(FE_OCP_RBN3077_FE_OFN807_n_46195), .b(n_6154), .c(FE_OFN774_n_46137), .d(n_6124), .o(n_46159) );
in01f80 g765114 ( .a(n_15084), .o(n_15163) );
no02f80 g772410 ( .a(n_8332), .b(n_8440), .o(n_8441) );
in01f80 g738465 ( .a(n_41472), .o(n_41548) );
na02f80 g774003 ( .a(n_6891), .b(n_6842), .o(n_6970) );
no02f80 g776247 ( .a(n_4698), .b(n_4194), .o(n_4851) );
in01f80 g743000 ( .a(n_37070), .o(n_36962) );
na02f80 g742074 ( .a(FE_OCP_RBN3441_n_37945), .b(n_38315), .o(n_38328) );
na02f80 g739199 ( .a(n_40701), .b(n_45181), .o(n_40792) );
no02f80 g779040 ( .a(n_2119), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .o(n_2149) );
no02f80 g774354 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_7_), .o(n_6570) );
in01f80 FE_OCPC1794_n_30612 ( .a(FE_OCPN1793_n_30612), .o(FE_OCPN1794_n_30612) );
no02f80 g760122 ( .a(n_20309), .b(n_20269), .o(n_20310) );
in01f80 g755118 ( .a(n_25350), .o(n_25351) );
na02f80 g752991 ( .a(n_27186), .b(n_27120), .o(n_27273) );
in01f80 g755195 ( .a(n_25712), .o(n_25713) );
in01f80 newInst_3274 ( .a(newNet_3273), .o(newNet_3274) );
no02f80 g742795 ( .a(n_37281), .b(n_37014), .o(n_37298) );
in01f80 g773836 ( .a(n_7153), .o(n_7131) );
no02f80 g756893 ( .a(n_23314), .b(n_23387), .o(n_23452) );
in01f80 g750789 ( .a(n_29192), .o(n_29215) );
no02f80 g747627 ( .a(n_33420), .b(n_33418), .o(n_33445) );
no02f80 g764402 ( .a(n_16195), .b(n_16223), .o(n_16398) );
no02f80 g765836 ( .a(n_14865), .b(n_13656), .o(n_14909) );
in01f80 g771457 ( .a(n_9633), .o(n_9634) );
no02f80 g763359 ( .a(n_17026), .b(n_17125), .o(n_17227) );
in01f80 FE_OCPC1753_n_7225 ( .a(n_7225), .o(FE_OCPN1753_n_7225) );
in01f80 g777361 ( .a(n_4721), .o(n_4722) );
na02f80 g776457 ( .a(n_4643), .b(n_4642), .o(n_4673) );
na02f80 g758294 ( .a(n_22249), .b(n_20614), .o(n_22507) );
in01f80 g754390 ( .a(n_25869), .o(n_25870) );
no02f80 g746060 ( .a(n_33901), .b(n_33921), .o(n_34010) );
na02f80 g743625 ( .a(n_36483), .b(n_36271), .o(n_36484) );
in01f80 newInst_453 ( .a(newNet_348), .o(newNet_453) );
no02f80 g757990 ( .a(n_22342), .b(n_22221), .o(n_22343) );
in01f80 FE_RC_2607_0 ( .a(n_17897), .o(FE_RN_1084_0) );
no02f80 g736856 ( .a(n_43362), .b(n_43510), .o(n_43617) );
ao12f80 g737084 ( .a(n_43097), .b(n_43083), .c(n_43121), .o(n_43162) );
in01f80 g763463 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .o(n_16990) );
oa12f80 g751351 ( .a(n_29458), .b(n_29457), .c(n_29456), .o(n_29851) );
ao12f80 g742664 ( .a(n_37498), .b(n_37497), .c(n_37496), .o(n_37948) );
oa22f80 FE_RC_764_0 ( .a(n_8381), .b(n_7546), .c(n_7545), .d(n_8382), .o(n_8498) );
in01f80 FE_RC_4204_0 ( .a(FE_RN_1840_0), .o(n_19589) );
no02f80 g758728 ( .a(n_22285), .b(n_21629), .o(n_22395) );
na02f80 g741466 ( .a(n_38746), .b(n_38721), .o(n_38770) );
in01f80 fopt783260 ( .a(n_44829), .o(n_44828) );
in01f80 newInst_3202 ( .a(newNet_3017), .o(newNet_3202) );
in01f80 g773387 ( .a(n_7732), .o(n_7733) );
na02f80 g737668 ( .a(FE_OCPN887_n_42367), .b(n_42065), .o(n_42726) );
na02f80 g765355 ( .a(n_15226), .b(n_15225), .o(n_15227) );
oa22f80 FE_RC_3407_0 ( .a(n_33643), .b(FE_OCP_RBN1353_n_33584), .c(n_33584), .d(n_33660), .o(n_33757) );
in01f80 g748292 ( .a(n_31685), .o(n_31686) );
in01f80 g737047 ( .a(n_43127), .o(n_43311) );
no02f80 FE_RC_2787_0 ( .a(n_34224), .b(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(FE_RN_1190_0) );
na02f80 g776840 ( .a(n_3855), .b(n_3765), .o(n_3856) );
in01f80 g745329 ( .a(n_36215), .o(n_36216) );
oa12f80 g736560 ( .a(n_345), .b(n_43656), .c(FE_OFN2_n_43918), .o(n_43694) );
no02f80 g768027 ( .a(n_12914), .b(n_12985), .o(n_13079) );
oa12f80 g757668 ( .a(n_22330), .b(n_22705), .c(n_22461), .o(n_22706) );
ao12f80 g739570 ( .a(n_40636), .b(n_40638), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n_41343) );
na02f80 g737565 ( .a(n_42442), .b(FE_OCPN885_n_42216), .o(n_42491) );
na02f80 FE_RC_2329_0 ( .a(FE_RN_888_0), .b(n_33382), .o(FE_RN_889_0) );
in01f80 g766282 ( .a(n_14334), .o(n_14335) );
in01f80 g769645 ( .a(n_47182), .o(n_11419) );
na02f80 g739436 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_), .o(n_40822) );
na02f80 g737930 ( .a(n_42201), .b(n_42321), .o(n_42413) );
in01f80 FE_RC_1304_0 ( .a(n_20343), .o(FE_RN_382_0) );
no02f80 g776309 ( .a(n_4680), .b(n_4246), .o(n_4752) );
ao12f80 g779457 ( .a(n_2126), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .o(n_2145) );
na02f80 g773710 ( .a(n_7236), .b(n_7122), .o(n_7267) );
ao12f80 g761628 ( .a(n_19525), .b(n_19524), .c(n_19523), .o(n_19607) );
no02f80 g746341 ( .a(n_33506), .b(n_33505), .o(n_33507) );
in01f80 newInst_965 ( .a(newNet_964), .o(newNet_965) );
na02f80 g752352 ( .a(n_27738), .b(n_27802), .o(n_27825) );
oa22f80 FE_RC_3759_0 ( .a(n_5389), .b(n_5250), .c(n_5249), .d(n_5361), .o(n_5531) );
oa22f80 g739737 ( .a(n_40509), .b(n_40174), .c(n_40510), .d(n_40173), .o(n_40549) );
na02f80 g779214 ( .a(n_1906), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .o(n_1968) );
in01f80 newInst_3698 ( .a(newNet_3697), .o(newNet_3698) );
in01f80 newInst_2593 ( .a(newNet_2592), .o(newNet_2593) );
ao12f80 g751433 ( .a(n_28407), .b(n_28428), .c(n_28406), .o(n_29644) );
na02f80 g768259 ( .a(n_12576), .b(n_12559), .o(n_12599) );
in01f80 FE_OCP_RBC1371_n_20763 ( .a(FE_OCP_RBN1370_n_20763), .o(FE_OCP_RBN1371_n_20763) );
in01f80 g775295 ( .a(n_5832), .o(n_5833) );
no02f80 g749090 ( .a(n_30963), .b(n_30911), .o(n_30987) );
oa12f80 g767423 ( .a(n_13396), .b(n_13395), .c(n_13394), .o(n_13476) );
oa12f80 g750540 ( .a(n_29497), .b(n_29496), .c(n_29495), .o(n_29555) );
in01f80 g763933 ( .a(n_17152), .o(n_17153) );
no02f80 g770250 ( .a(n_46989), .b(FE_OCP_RBN2613_n_9075), .o(n_10891) );
oa22f80 g744710 ( .a(n_36495), .b(n_36172), .c(n_36494), .d(n_36173), .o(n_36573) );
na02f80 g780585 ( .a(n_745), .b(n_783), .o(n_829) );
in01f80 g761582 ( .a(n_22580), .o(n_22907) );
oa12f80 g773567 ( .a(n_7410), .b(n_7409), .c(n_7408), .o(n_7812) );
no02f80 g745227 ( .a(n_36025), .b(n_35930), .o(n_36125) );
no02f80 g753528 ( .a(n_26846), .b(n_26799), .o(n_26839) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_14_ ( .ck(newNet_3442), .d(n_27472), .o(delay_add_ln22_unr17_stage7_stallmux_q_14_) );
oa12f80 g780527 ( .a(n_710), .b(n_890), .c(n_701), .o(n_1084) );
in01f80 g759666 ( .a(n_20553), .o(n_20548) );
in01f80 g756711 ( .a(n_23517), .o(n_23518) );
no02f80 FE_RC_1617_0 ( .a(FE_RN_450_0), .b(FE_RN_451_0), .o(FE_RN_452_0) );
oa12f80 g779336 ( .a(n_1627), .b(n_1635), .c(n_1626), .o(n_2276) );
ao22s80 g761848 ( .a(n_18360), .b(n_18198), .c(n_18318), .d(n_18199), .o(n_18515) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_21_ ( .ck(newNet_3528), .d(n_22750), .o(delay_add_ln22_unr14_stage6_stallmux_q_21_) );
in01f80 g767040 ( .a(n_13821), .o(n_13822) );
na02f80 g771373 ( .a(n_9345), .b(n_9376), .o(n_9425) );
na02f80 g750140 ( .a(n_29845), .b(n_29844), .o(n_29925) );
in01f80 g769169 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_6_), .o(n_11689) );
ao12f80 g778989 ( .a(n_1561), .b(n_2074), .c(n_1516), .o(n_2129) );
in01f80 g764372 ( .a(n_16390), .o(n_16391) );
na02f80 g762092 ( .a(FE_OCP_RBN2205_n_18242), .b(n_17806), .o(n_18460) );
no02f80 g773071 ( .a(n_7997), .b(n_7918), .o(n_7998) );
na02f80 g765406 ( .a(n_15050), .b(n_15054), .o(n_15151) );
no02f80 g759298 ( .a(n_21214), .b(n_21175), .o(n_21261) );
no02f80 g761696 ( .a(n_19404), .b(n_18571), .o(n_19494) );
in01f80 FE_OFC823_n_15791 ( .a(FE_OFN841_n_15791), .o(FE_OFN823_n_15791) );
no02f80 g772939 ( .a(n_7884), .b(n_7883), .o(n_7987) );
na02f80 g780614 ( .a(n_713), .b(n_757), .o(n_842) );
na02f80 g765794 ( .a(FE_OCP_RBN1165_n_13726), .b(n_14921), .o(n_15035) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_2_ ( .ck(newNet_2532), .d(n_26491), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_) );
in01f80 g737022 ( .a(n_43133), .o(n_43174) );
oa22f80 FE_RC_907_0 ( .a(n_25824), .b(n_25729), .c(FE_OFN738_n_22641), .d(n_25728), .o(n_25847) );
na02f80 g771585 ( .a(n_8884), .b(n_8309), .o(n_8979) );
na02f80 FE_RC_44_0 ( .a(n_2539), .b(FE_RN_11_0), .o(n_47026) );
in01f80 FE_RC_1400_0 ( .a(n_15999), .o(FE_RN_409_0) );
in01f80 g774313 ( .a(n_6716), .o(n_6547) );
in01f80 FE_OCPC1443_n_45050 ( .a(n_45050), .o(FE_OCPN1443_n_45050) );
na02f80 g765134 ( .a(n_15204), .b(FE_OCP_RBN2507_n_13896), .o(n_15205) );
no02f80 FE_RC_2445_0 ( .a(n_13034), .b(n_13035), .o(FE_RN_976_0) );
in01f80 g772861 ( .a(n_8102), .o(n_8103) );
in01f80 FE_OCP_RBC3798_delay_xor_ln22_unr12_stage5_stallmux_q_0_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(FE_OCP_RBN3798_delay_xor_ln22_unr12_stage5_stallmux_q_0_) );
in01f80 FE_OCPC1768_n_29715 ( .a(FE_OCPN1767_n_29715), .o(FE_OCPN1768_n_29715) );
na02f80 g761344 ( .a(n_18924), .b(n_47247), .o(n_19002) );
na02f80 g754939 ( .a(n_25149), .b(n_24054), .o(n_25242) );
na02f80 g743646 ( .a(n_36410), .b(n_36103), .o(n_36483) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_16_ ( .ck(newNet_1128), .d(n_10717), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_) );
oa22f80 g769742 ( .a(n_11267), .b(n_10296), .c(n_11233), .d(n_10297), .o(n_11305) );
in01f80 g780286 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_), .o(n_2483) );
no03m80 FE_RC_834_0 ( .a(n_9495), .b(FE_RN_1198_0), .c(FE_OCP_RBN2587_n_9492), .o(n_9577) );
in01f80 g756565 ( .a(n_23664), .o(n_23634) );
oa22f80 g768852 ( .a(n_11833), .b(n_11773), .c(n_11927), .d(n_11772), .o(n_12021) );
no02f80 g763400 ( .a(FE_OCPN1756_n_16923), .b(n_15992), .o(n_17388) );
na02f80 FE_RC_2019_0 ( .a(n_20321), .b(FE_RN_664_0), .o(FE_RN_669_0) );
in01f80 newInst_2332 ( .a(newNet_2331), .o(newNet_2332) );
in01f80 g748868 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n_32357) );
oa22f80 FE_RC_3191_0 ( .a(n_18259), .b(n_18654), .c(n_18653), .d(n_18260), .o(n_18866) );
in01f80 newInst_2579 ( .a(newNet_2578), .o(newNet_2579) );
in01f80 g761494 ( .a(n_20082), .o(n_20083) );
na02f80 g758581 ( .a(n_22034), .b(n_22065), .o(n_22094) );
na02f80 g775093 ( .a(n_6012), .b(n_6006), .o(n_6119) );
oa22f80 g771331 ( .a(n_8942), .b(n_7764), .c(n_8941), .d(n_7765), .o(n_9090) );
in01f80 g768665 ( .a(n_12197), .o(n_12116) );
no02f80 g760455 ( .a(n_20026), .b(n_19969), .o(n_20048) );
oa22f80 FE_RC_3744_0 ( .a(n_14889), .b(n_14852), .c(n_14874), .d(n_14890), .o(n_14991) );
na02f80 g748640 ( .a(n_31421), .b(n_31441), .o(n_31442) );
in01f80 g737278 ( .a(n_42902), .o(n_42916) );
in01f80 g757056 ( .a(n_23722), .o(n_23697) );
in01f80 g748513 ( .a(n_31700), .o(n_31701) );
in01f80 newInst_3328 ( .a(newNet_476), .o(newNet_3328) );
oa12f80 g780330 ( .a(n_686), .b(n_739), .c(n_689), .o(n_786) );
no02f80 g748282 ( .a(FE_OCP_RBN3084_n_31819), .b(FE_OCP_RBN2888_n_46957), .o(n_31967) );
in01f80 g745712 ( .a(n_34367), .o(n_34368) );
no02f80 g737767 ( .a(n_42283), .b(n_42306), .o(n_42721) );
in01f80 FE_RC_3562_0 ( .a(FE_RN_1547_0), .o(n_25066) );
in01f80 g770398 ( .a(n_10405), .o(n_10406) );
no02f80 g757356 ( .a(n_23100), .b(delay_add_ln22_unr14_stage6_stallmux_q_3_), .o(n_23124) );
no02f80 g755694 ( .a(n_24403), .b(n_24053), .o(n_24467) );
in01f80 FE_RC_4022_0 ( .a(FE_OFN738_n_22641), .o(FE_RN_1747_0) );
na02f80 g757028 ( .a(n_23803), .b(n_23802), .o(n_23864) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_27_ ( .ck(newNet_2457), .d(n_32546), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_) );
in01f80 g777896 ( .a(n_4022), .o(n_3301) );
in01f80 g764463 ( .a(n_16653), .o(n_16673) );
no02f80 g748967 ( .a(n_30919), .b(n_30858), .o(n_30967) );
in01f80 FE_OCPC3180_FE_OCP_RBN2744_n_15319 ( .a(FE_OCPN3179_FE_OCP_RBN2744_n_15319), .o(FE_OCPN3180_FE_OCP_RBN2744_n_15319) );
no02f80 g771161 ( .a(n_9739), .b(n_9702), .o(n_9907) );
ao12f80 g754588 ( .a(n_26551), .b(n_26856), .c(n_26510), .o(n_26892) );
in01f80 FE_OCP_RBC2882_n_26318 ( .a(n_26318), .o(FE_OCP_RBN2882_n_26318) );
oa22f80 g784559 ( .a(FE_OFN800_n_46285), .b(n_10680), .c(FE_OCP_RBN3709_n_46337), .d(n_10631), .o(n_46380) );
na02f80 g749574 ( .a(n_30486), .b(n_30485), .o(n_30487) );
na02f80 g750550 ( .a(n_29475), .b(n_29477), .o(n_29478) );
no02f80 g766535 ( .a(n_14090), .b(n_14057), .o(n_14233) );
in01f80 g761004 ( .a(n_19327), .o(n_19328) );
no02f80 g750080 ( .a(n_29896), .b(n_29442), .o(n_30318) );
no02f80 g743338 ( .a(n_36660), .b(n_36614), .o(n_36677) );
ao22s80 g784753 ( .a(n_7687), .b(n_7310), .c(n_7686), .d(n_7309), .o(n_47235) );
in01f80 newInst_1655 ( .a(newNet_1654), .o(newNet_1655) );
in01f80 g744370 ( .a(n_46216), .o(n_36814) );
ao12f80 g776073 ( .a(n_4557), .b(n_4558), .c(n_4296), .o(n_4605) );
na02f80 g755320 ( .a(n_24810), .b(n_24754), .o(n_24842) );
oa12f80 g746113 ( .a(n_35112), .b(n_35111), .c(n_35110), .o(n_35675) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_1_ ( .ck(newNet_238), .d(n_46169), .o(delay_xor_ln22_unr6_stage3_stallmux_q_1_) );
in01f80 g779293 ( .a(n_1760), .o(n_1761) );
ms00f80 sin_out_reg_11_ ( .ck(newNet_88), .d(n_43805), .o(sin_out_11) );
na02f80 g773181 ( .a(n_7615), .b(n_7630), .o(n_7665) );
no02f80 g752188 ( .a(FE_OCP_RBN2126_n_44734), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .o(n_28226) );
in01f80 newInst_1880 ( .a(newNet_1879), .o(newNet_1880) );
na02f80 FE_RC_2416_0 ( .a(n_7134), .b(FE_RN_954_0), .o(n_7470) );
in01f80 g767310 ( .a(n_13569), .o(n_13525) );
no02f80 g742914 ( .a(n_36971), .b(n_37016), .o(n_37301) );
na02f80 g769094 ( .a(n_11459), .b(n_11007), .o(n_11499) );
oa12f80 g754595 ( .a(n_26690), .b(FE_OCP_RBN3704_n_26231), .c(n_25605), .o(n_26943) );
in01f80 FE_OCP_RBC3524_n_8242 ( .a(FE_OCP_RBN3523_n_8242), .o(FE_OCP_RBN3524_n_8242) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_13_ ( .ck(newNet_1873), .d(n_16616), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_) );
in01f80 FE_OCP_RBC2180_FE_RN_526_0 ( .a(FE_RN_526_0), .o(FE_OCP_RBN2180_FE_RN_526_0) );
no02f80 g770807 ( .a(n_10050), .b(n_10092), .o(n_10093) );
na02f80 g776595 ( .a(n_4438), .b(n_4437), .o(n_4594) );
na02f80 g767783 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_28_), .o(n_13101) );
no02f80 g753985 ( .a(n_26277), .b(n_26205), .o(n_26316) );
oa12f80 g742818 ( .a(n_36967), .b(n_37223), .c(n_37013), .o(n_37245) );
in01f80 g776731 ( .a(n_4165), .o(n_4240) );
in01f80 g767397 ( .a(n_13478), .o(n_13479) );
no02f80 g775129 ( .a(n_5693), .b(n_4759), .o(n_5734) );
in01f80 g780251 ( .a(n_1088), .o(n_1127) );
na02f80 g776625 ( .a(n_4011), .b(n_3029), .o(n_4092) );
no02f80 g774821 ( .a(n_6228), .b(n_5780), .o(n_6330) );
in01f80 g740357 ( .a(n_39753), .o(n_39754) );
in01f80 FE_OCP_RBC2318_n_2367 ( .a(n_2367), .o(FE_OCP_RBN2318_n_2367) );
na02f80 g740376 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39465), .o(n_40270) );
in01f80 g741607 ( .a(n_38658), .o(n_38659) );
na02f80 g753730 ( .a(n_26526), .b(n_26525), .o(n_26527) );
in01f80 g760346 ( .a(n_20894), .o(n_20895) );
in01f80 g738851 ( .a(n_41349), .o(n_41348) );
in01f80 g748962 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n_32318) );
no02f80 FE_RC_1845_0 ( .a(n_35755), .b(n_35754), .o(FE_RN_561_0) );
in01f80 g762112 ( .a(n_18309), .o(n_18310) );
in01f80 g737256 ( .a(n_42907), .o(n_42908) );
ao12f80 g777747 ( .a(n_3061), .b(n_3232), .c(n_3109), .o(n_3303) );
oa12f80 g752016 ( .a(n_28165), .b(n_28164), .c(n_28163), .o(n_29187) );
no02f80 g765637 ( .a(n_15481), .b(n_15442), .o(n_15443) );
na02f80 g764577 ( .a(n_15992), .b(n_14650), .o(n_16044) );
in01f80 g745689 ( .a(n_34291), .o(n_34315) );
na02f80 g777036 ( .a(n_3608), .b(n_3632), .o(n_3746) );
na03f80 FE_RC_1683_0 ( .a(n_6187), .b(n_6162), .c(n_6188), .o(n_6189) );
in01f80 g741553 ( .a(n_38678), .o(n_38679) );
oa22f80 g758561 ( .a(n_22523), .b(n_21853), .c(n_22524), .d(n_21854), .o(n_22587) );
na02f80 g750120 ( .a(FE_OCP_RBN2572_n_29922), .b(n_30136), .o(n_30170) );
na02f80 g740235 ( .a(n_39835), .b(n_39894), .o(n_39895) );
in01f80 FE_OCP_RBC2747_n_9584 ( .a(n_9584), .o(FE_OCP_RBN2747_n_9584) );
na02f80 g760217 ( .a(n_20249), .b(FE_OCP_RBN1688_n_18986), .o(n_20311) );
na02f80 g741960 ( .a(n_47336), .b(n_38120), .o(n_38166) );
na02f80 g779006 ( .a(n_2180), .b(n_2142), .o(n_2192) );
na02f80 g761884 ( .a(n_18405), .b(FE_OFN778_n_17093), .o(n_18433) );
in01f80 newInst_3393 ( .a(newNet_3392), .o(newNet_3393) );
in01f80 newInst_1965 ( .a(newNet_1964), .o(newNet_1965) );
oa12f80 g772541 ( .a(n_7928), .b(n_8337), .c(n_7914), .o(n_8649) );
na02f80 FE_RC_1009_0 ( .a(FE_RN_291_0), .b(FE_RN_292_0), .o(FE_RN_293_0) );
ao22s80 FE_RC_1358_0 ( .a(n_5136), .b(n_5532), .c(n_5137), .d(n_5533), .o(n_5627) );
in01f80 FE_OCP_RBC2910_n_26394 ( .a(n_26394), .o(FE_OCP_RBN2910_n_26394) );
na02f80 g760508 ( .a(n_20451), .b(n_19821), .o(n_20513) );
na02f80 g750812 ( .a(n_29095), .b(n_28718), .o(n_29120) );
na02f80 g748985 ( .a(n_31149), .b(n_31148), .o(n_31150) );
in01f80 FE_RC_532_0 ( .a(n_22560), .o(FE_RN_166_0) );
in01f80 newInst_177 ( .a(newNet_176), .o(newNet_177) );
in01f80 FE_OCP_RBC3132_n_27736 ( .a(n_27736), .o(FE_OCP_RBN3132_n_27736) );
no02f80 g776903 ( .a(n_3877), .b(FE_OCP_RBN3577_n_4528), .o(n_3965) );
na02f80 g758079 ( .a(n_22005), .b(FE_OCPN1416_FE_OCP_RBN1362_n_20504), .o(n_22085) );
na02f80 g740161 ( .a(FE_OCP_RBN3055_n_39913), .b(n_39900), .o(n_39980) );
oa12f80 g738824 ( .a(n_41298), .b(n_44429), .c(n_41349), .o(n_41359) );
na02f80 g764873 ( .a(n_15551), .b(n_15545), .o(n_15620) );
in01f80 g762336 ( .a(n_18075), .o(n_18076) );
na02f80 g759632 ( .a(n_20719), .b(n_45012), .o(n_20842) );
oa12f80 g747948 ( .a(n_33090), .b(n_33089), .c(n_33088), .o(n_33169) );
na03f80 FE_RC_3792_0 ( .a(n_29952), .b(n_29956), .c(n_30021), .o(n_30022) );
in01f80 newInst_981 ( .a(newNet_980), .o(newNet_981) );
in01f80 g758929 ( .a(n_21430), .o(n_21661) );
in01f80 g740321 ( .a(n_39770), .o(n_39781) );
na02f80 g761931 ( .a(n_18969), .b(n_18968), .o(n_18970) );
na02f80 g775425 ( .a(n_5820), .b(n_4700), .o(n_6001) );
oa12f80 g741705 ( .a(n_38482), .b(n_38481), .c(n_38480), .o(n_39040) );
oa12f80 g781276 ( .a(n_7), .b(beta_20), .c(beta_19), .o(n_104) );
in01f80 g775849 ( .a(n_5350), .o(n_5408) );
in01f80 FE_OCP_RBC2865_n_39640 ( .a(n_39640), .o(FE_OCP_RBN2865_n_39640) );
ao12f80 g746353 ( .a(n_33235), .b(n_33559), .c(n_33200), .o(n_33638) );
in01f80 newInst_719 ( .a(newNet_150), .o(newNet_719) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_5_ ( .ck(newNet_1949), .d(n_10213), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_) );
in01f80 newInst_1524 ( .a(newNet_1523), .o(newNet_1524) );
in01f80 g751656 ( .a(n_28438), .o(n_28467) );
na02f80 g758946 ( .a(n_21640), .b(FE_OCP_DRV_N1602_n_21639), .o(n_21727) );
in01f80 FE_OCP_RBC1325_n_29056 ( .a(FE_OCP_RBN1324_n_29056), .o(FE_OCP_RBN1325_n_29056) );
oa12f80 g750605 ( .a(n_28784), .b(n_29353), .c(n_28828), .o(n_29383) );
in01f80 g773616 ( .a(n_7363), .o(n_7348) );
na02f80 g768681 ( .a(n_12039), .b(n_12038), .o(n_12040) );
na02f80 g752506 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(n_27642) );
oa22f80 g784556 ( .a(FE_OFN800_n_46285), .b(n_11177), .c(FE_OCP_RBN3710_n_46337), .d(n_11151), .o(n_46377) );
no02f80 g755633 ( .a(n_24546), .b(n_24633), .o(n_24635) );
in01f80 g770002 ( .a(n_10991), .o(n_10978) );
na02f80 g769032 ( .a(FE_OCP_RBN2006_n_45209), .b(n_45224), .o(n_11786) );
ao12f80 g756632 ( .a(n_23508), .b(n_23507), .c(n_23506), .o(n_24893) );
na02f80 g766467 ( .a(n_14068), .b(n_14095), .o(n_14176) );
in01f80 newInst_137 ( .a(newNet_136), .o(newNet_137) );
oa12f80 g741821 ( .a(n_38367), .b(n_38366), .c(n_38365), .o(n_38890) );
in01f80 newInst_1204 ( .a(newNet_1203), .o(newNet_1204) );
oa22f80 g753471 ( .a(n_27537), .b(n_26790), .c(n_27538), .d(n_26791), .o(n_27574) );
in01f80 newInst_3575 ( .a(newNet_684), .o(newNet_3575) );
no03m80 FE_RC_1404_0 ( .a(n_44158), .b(n_21030), .c(n_21153), .o(n_46967) );
in01f80 g745656 ( .a(n_35461), .o(n_35462) );
no02f80 g765059 ( .a(n_15977), .b(n_15926), .o(n_16384) );
na02f80 FE_RC_2546_0 ( .a(FE_RN_1042_0), .b(n_39165), .o(FE_RN_1043_0) );
in01f80 newInst_3469 ( .a(newNet_3468), .o(newNet_3469) );
in01f80 g748616 ( .a(n_31544), .o(n_31545) );
no02f80 g751794 ( .a(n_28299), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .o(n_28341) );
no02f80 g756360 ( .a(n_24417), .b(n_24383), .o(n_24384) );
na02f80 g777923 ( .a(n_3194), .b(n_3175), .o(n_3275) );
no02f80 FE_RC_2128_0 ( .a(FE_RN_742_0), .b(n_25732), .o(n_25786) );
oa12f80 g749597 ( .a(n_30055), .b(n_30483), .c(n_30022), .o(n_30302) );
in01f80 g736869 ( .a(n_43609), .o(n_43610) );
in01f80 FE_OCP_RBC3579_n_44944 ( .a(FE_OCP_RBN2545_n_44944), .o(FE_OCP_RBN3579_n_44944) );
ao12f80 g762660 ( .a(n_17929), .b(FE_OCP_RBN2145_FE_OCPN861_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_15_), .o(n_17950) );
oa22f80 g739730 ( .a(n_40462), .b(n_40077), .c(n_40463), .d(n_40076), .o(n_40498) );
na02f80 FE_RC_506_0 ( .a(FE_RN_153_0), .b(FE_RN_154_0), .o(FE_RN_155_0) );
na02f80 g768420 ( .a(n_12361), .b(n_12059), .o(n_12362) );
in01f80 FE_RC_411_0 ( .a(n_14194), .o(FE_RN_121_0) );
na02f80 g745961 ( .a(n_34031), .b(n_34063), .o(n_34088) );
na02f80 g754421 ( .a(n_25636), .b(n_25402), .o(n_25702) );
na02f80 g753230 ( .a(n_27207), .b(n_26165), .o(n_27382) );
na02f80 g749247 ( .a(n_30652), .b(n_30537), .o(n_30683) );
in01f80 g771536 ( .a(n_9398), .o(n_9399) );
ao22s80 FE_RC_1469_0 ( .a(n_17213), .b(n_17275), .c(n_17287), .d(n_17214), .o(n_17475) );
in01f80 newInst_2086 ( .a(newNet_2085), .o(newNet_2086) );
na02f80 FE_RC_1808_0 ( .a(n_11983), .b(n_12026), .o(FE_RN_536_0) );
in01f80 g770690 ( .a(n_10322), .o(n_10323) );
na02f80 g762230 ( .a(n_18092), .b(n_18136), .o(n_18149) );
oa12f80 g743666 ( .a(n_36072), .b(n_36411), .c(n_35911), .o(n_36437) );
no02f80 g755177 ( .a(n_25020), .b(n_25049), .o(n_25021) );
na02f80 g747953 ( .a(n_33089), .b(n_33088), .o(n_33090) );
no02f80 g771748 ( .a(n_8790), .b(n_8189), .o(n_8791) );
in01f80 g752325 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_), .o(n_28646) );
na02f80 g759179 ( .a(n_21188), .b(n_21222), .o(n_21272) );
na02f80 g755726 ( .a(n_24325), .b(n_23820), .o(n_24326) );
in01f80 FE_OCP_DRV_C1555_n_19384 ( .a(n_19384), .o(FE_OCP_DRV_N1555_n_19384) );
in01f80 FE_OCP_RBC2126_n_44734 ( .a(FE_OCP_RBN3367_n_44722), .o(FE_OCP_RBN2126_n_44734) );
na02f80 g761465 ( .a(n_19647), .b(n_19790), .o(n_19905) );
na02f80 g747217 ( .a(n_32829), .b(delay_add_ln22_unr20_stage8_stallmux_q_4_), .o(n_32884) );
in01f80 g758783 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .o(n_22208) );
na02f80 g760676 ( .a(n_19706), .b(n_19672), .o(n_19808) );
na02f80 g738542 ( .a(n_41761), .b(n_41723), .o(n_41784) );
no02f80 g753919 ( .a(n_26222), .b(n_26260), .o(n_26358) );
na02f80 g763458 ( .a(n_17171), .b(n_17114), .o(n_17311) );
ao12f80 g739392 ( .a(n_40771), .b(FE_OCPN897_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n_41303) );
in01f80 g736841 ( .a(n_43028), .o(n_43040) );
no02f80 g750617 ( .a(n_29397), .b(n_29443), .o(n_29496) );
in01f80 FE_RC_666_0 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .o(FE_RN_210_0) );
in01f80 newInst_3246 ( .a(newNet_3245), .o(newNet_3246) );
ao22s80 FE_RC_3032_0 ( .a(FE_RN_1327_0), .b(n_11870), .c(n_11850), .d(n_11810), .o(n_12060) );
na02f80 g751738 ( .a(n_28304), .b(n_28222), .o(n_28363) );
in01f80 g743144 ( .a(n_37104), .o(n_37028) );
in01f80 FE_OCP_RBC3410_n_45120 ( .a(n_45120), .o(FE_OCP_RBN3410_n_45120) );
na02f80 g773235 ( .a(n_7633), .b(n_7621), .o(n_7657) );
in01f80 g740338 ( .a(n_40390), .o(n_40391) );
in01f80 newInst_1977 ( .a(newNet_1976), .o(newNet_1977) );
in01f80 newInst_852 ( .a(newNet_851), .o(newNet_852) );
no02f80 g747194 ( .a(n_32849), .b(n_32848), .o(n_32850) );
na02f80 g742474 ( .a(n_37715), .b(n_37688), .o(n_37732) );
oa12f80 g737546 ( .a(n_42449), .b(n_42422), .c(n_42367), .o(n_42510) );
na02f80 g742447 ( .a(n_37717), .b(n_37691), .o(n_37718) );
in01f80 g777026 ( .a(n_3583), .o(n_3584) );
oa12f80 g740991 ( .a(n_38926), .b(n_38963), .c(n_39002), .o(n_39106) );
ao12f80 g747991 ( .a(n_32456), .b(n_33000), .c(n_32487), .o(n_33089) );
no02f80 g747543 ( .a(n_33375), .b(n_33758), .o(n_33793) );
in01f80 g775882 ( .a(n_5233), .o(n_5276) );
na02f80 g764345 ( .a(n_16482), .b(n_16451), .o(n_16575) );
in01f80 g779480 ( .a(n_1996), .o(n_1997) );
in01f80 g772525 ( .a(n_8487), .o(n_8509) );
na02f80 g758208 ( .a(n_22407), .b(n_22375), .o(n_22490) );
na02f80 g770498 ( .a(n_10332), .b(n_10104), .o(n_10368) );
in01f80 FE_OCP_RBC2009_n_45622 ( .a(n_45622), .o(FE_OCP_RBN2009_n_45622) );
ao22s80 FE_RC_2958_0 ( .a(n_11370), .b(FE_OCP_RBN3049_n_11329), .c(FE_RN_1291_0), .d(n_11329), .o(n_11475) );
na02f80 g738858 ( .a(n_41332), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41333) );
in01f80 g761558 ( .a(n_18950), .o(n_18859) );
oa12f80 g739512 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .b(FE_OCP_RBN2134_n_45508), .c(FE_OCP_RBN3337_n_44610), .o(n_40662) );
na02f80 g745126 ( .a(n_34663), .b(n_34662), .o(n_34664) );
in01f80 newInst_2948 ( .a(newNet_2947), .o(newNet_2948) );
in01f80 FE_RC_647_0 ( .a(n_37078), .o(FE_RN_205_0) );
in01f80 g776226 ( .a(n_4860), .o(n_4861) );
no02f80 g768389 ( .a(n_12463), .b(n_12462), .o(n_12479) );
oa12f80 g749722 ( .a(n_31311), .b(n_31411), .c(n_31410), .o(n_31412) );
no03m80 FE_RC_661_0 ( .a(n_43692), .b(n_43256), .c(n_43664), .o(n_43721) );
ao12f80 g774207 ( .a(n_6951), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .o(n_7113) );
no02f80 g770885 ( .a(n_9892), .b(FE_RN_1433_0), .o(n_9937) );
na02f80 g764220 ( .a(n_16462), .b(n_16436), .o(n_16527) );
in01f80 FE_OCPC1767_n_29715 ( .a(n_29715), .o(FE_OCPN1767_n_29715) );
in01f80 newInst_2787 ( .a(newNet_2786), .o(newNet_2787) );
in01f80 g756463 ( .a(n_23925), .o(n_23926) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_13_ ( .ck(newNet_1135), .d(n_10632), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_) );
in01f80 newInst_2058 ( .a(newNet_2057), .o(newNet_2058) );
in01f80 newInst_2204 ( .a(newNet_2203), .o(newNet_2204) );
na02f80 g776918 ( .a(n_3948), .b(n_3884), .o(n_4005) );
no02f80 g779056 ( .a(FE_OCP_RBN3412_n_2100), .b(n_1861), .o(n_2163) );
na02f80 g754729 ( .a(n_26541), .b(n_26033), .o(n_26898) );
in01f80 newInst_419 ( .a(newNet_418), .o(newNet_419) );
in01f80 g776102 ( .a(n_4975), .o(n_4976) );
in01f80 g760693 ( .a(n_19703), .o(n_19975) );
na02f80 g760798 ( .a(n_19537), .b(n_19468), .o(n_19637) );
in01f80 g744208 ( .a(n_36254), .o(n_36255) );
na02f80 g760921 ( .a(n_19286), .b(n_19285), .o(n_19287) );
ao12f80 g751502 ( .a(n_28490), .b(n_28817), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .o(n_28912) );
na02f80 g753094 ( .a(n_27426), .b(n_27425), .o(n_27467) );
no02f80 g766139 ( .a(n_14868), .b(n_14387), .o(n_14948) );
na02f80 g779755 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .o(n_1715) );
ao12f80 g775840 ( .a(n_4676), .b(n_5364), .c(n_4716), .o(n_5452) );
no02f80 g742394 ( .a(n_37745), .b(FE_OCPN1778_n_37744), .o(n_37767) );
na02f80 g748123 ( .a(n_31783), .b(n_31874), .o(n_31933) );
in01f80 g779541 ( .a(n_1519), .o(n_1520) );
in01f80 g763205 ( .a(n_17395), .o(n_17396) );
na02f80 g748039 ( .a(n_31935), .b(n_31766), .o(n_31974) );
na02f80 g764926 ( .a(n_15585), .b(n_15538), .o(n_15645) );
no02f80 g758036 ( .a(n_22846), .b(n_22845), .o(n_22847) );
in01f80 g744678 ( .a(n_35272), .o(n_35288) );
oa12f80 g755666 ( .a(n_24448), .b(n_24447), .c(n_24446), .o(n_26248) );
oa22f80 FE_RC_1630_0 ( .a(n_22801), .b(n_22818), .c(n_22793), .d(n_22791), .o(n_22894) );
in01f80 newInst_2131 ( .a(newNet_1355), .o(newNet_2131) );
ao12f80 g777715 ( .a(n_3436), .b(n_3435), .c(n_3434), .o(n_4760) );
in01f80 newInst_205 ( .a(newNet_164), .o(newNet_205) );
na02f80 g772363 ( .a(n_8627), .b(n_8626), .o(n_8657) );
no02f80 g771942 ( .a(n_8803), .b(FE_OCP_RBN2305_n_7817), .o(n_8805) );
oa12f80 g752162 ( .a(n_28560), .b(n_28559), .c(n_28558), .o(n_28982) );
na02f80 g745831 ( .a(n_44104), .b(n_33844), .o(n_34241) );
na02f80 g738268 ( .a(n_41846), .b(n_41641), .o(n_41896) );
ao12f80 g782637 ( .a(n_44875), .b(n_38270), .c(n_37595), .o(n_44030) );
no02f80 g745530 ( .a(n_34403), .b(n_34322), .o(n_34789) );
in01f80 newInst_2092 ( .a(newNet_2091), .o(newNet_2092) );
in01f80 g777631 ( .a(n_3648), .o(n_3649) );
in01f80 g747579 ( .a(n_33498), .o(n_33556) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_13_ ( .ck(newNet_2413), .d(n_36371), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_) );
oa12f80 g761838 ( .a(n_18202), .b(n_18269), .c(n_18171), .o(n_18322) );
oa12f80 g736541 ( .a(n_341), .b(n_43660), .c(FE_OFN2_n_43918), .o(n_43695) );
in01f80 g758049 ( .a(n_23116), .o(n_22952) );
oa12f80 g768773 ( .a(n_11598), .b(n_11914), .c(n_11520), .o(n_11986) );
in01f80 g764792 ( .a(n_15804), .o(n_15851) );
na02f80 g759009 ( .a(n_21391), .b(n_21470), .o(n_21392) );
oa12f80 g777215 ( .a(n_3527), .b(n_3526), .c(n_3525), .o(n_3605) );
na02f80 g759398 ( .a(n_20974), .b(n_20998), .o(n_21118) );
no02f80 g775586 ( .a(n_5746), .b(FE_OCP_RBN2788_n_4294), .o(n_5891) );
no02f80 g757342 ( .a(n_44068), .b(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .o(n_23131) );
in01f80 FE_OCP_RBC2247_n_13017 ( .a(FE_OCP_RBN2243_n_13017), .o(FE_OCP_RBN2247_n_13017) );
in01f80 g747447 ( .a(n_32630), .o(n_32661) );
na02f80 g776776 ( .a(n_3933), .b(n_3106), .o(n_4133) );
na02f80 FE_RC_2583_0 ( .a(FE_RN_1058_0), .b(FE_RN_1066_0), .o(n_3456) );
in01f80 g775100 ( .a(n_6076), .o(n_6096) );
no02f80 g772577 ( .a(n_8296), .b(FE_OCPN890_n_7802), .o(n_8306) );
na02f80 FE_RC_2298_0 ( .a(n_25135), .b(FE_RN_865_0), .o(FE_RN_866_0) );
no02f80 FE_RC_2180_0 ( .a(FE_RN_778_0), .b(n_26920), .o(n_26879) );
no02f80 g752617 ( .a(n_28206), .b(n_27959), .o(n_28298) );
no02f80 g764446 ( .a(FE_OCP_RBN3690_n_16146), .b(FE_OCPN3775_n_14730), .o(n_16223) );
ao22s80 g756704 ( .a(n_23463), .b(n_23141), .c(n_23482), .d(n_23140), .o(n_23561) );
no02f80 g740670 ( .a(n_39569), .b(n_39588), .o(n_39628) );
in01f80 newInst_1215 ( .a(newNet_1214), .o(newNet_1215) );
in01f80 g770481 ( .a(n_10369), .o(n_10542) );
no02f80 g769191 ( .a(n_11974), .b(n_11973), .o(n_12567) );
in01f80 newInst_2783 ( .a(newNet_2719), .o(newNet_2783) );
no02f80 g746399 ( .a(n_33501), .b(n_33203), .o(n_33536) );
in01f80 FE_OCP_RBC2155_n_1602 ( .a(n_1602), .o(FE_OCP_RBN2155_n_1602) );
na02f80 g740105 ( .a(n_40002), .b(n_40181), .o(n_40283) );
in01f80 FE_OCP_RBC3121_n_32239 ( .a(n_32239), .o(FE_OCP_RBN3121_n_32239) );
na02f80 g770201 ( .a(n_10594), .b(n_10622), .o(n_10730) );
in01f80 g763554 ( .a(n_16923), .o(n_16975) );
in01f80 g764120 ( .a(n_16960), .o(n_16961) );
no02f80 g740860 ( .a(n_39399), .b(n_39047), .o(n_39400) );
in01f80 FE_OCP_RBC2832_n_26081 ( .a(n_26081), .o(FE_OCP_RBN2832_n_26081) );
in01f80 newInst_2952 ( .a(newNet_2951), .o(newNet_2952) );
in01f80 FE_RC_1779_0 ( .a(n_1936), .o(FE_RN_518_0) );
in01f80 g757879 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .o(n_22354) );
na02f80 g744983 ( .a(n_34946), .b(n_30545), .o(n_34975) );
na02f80 g778459 ( .a(n_2372), .b(n_2347), .o(n_2467) );
ao12f80 g740946 ( .a(n_38821), .b(n_39065), .c(n_38864), .o(n_39338) );
na02f80 g754838 ( .a(n_25564), .b(n_25973), .o(n_25565) );
in01f80 newInst_949 ( .a(newNet_948), .o(newNet_949) );
in01f80 g755100 ( .a(n_25206), .o(n_25231) );
no02f80 g747804 ( .a(n_33372), .b(n_33170), .o(n_33990) );
no02f80 g755234 ( .a(n_25038), .b(n_25036), .o(n_25068) );
in01f80 g749316 ( .a(n_30735), .o(n_30736) );
na02f80 g766485 ( .a(n_14023), .b(n_13441), .o(n_14068) );
in01f80 FE_RC_2193_0 ( .a(n_31234), .o(FE_RN_786_0) );
in01f80 g760542 ( .a(n_19921), .o(n_19946) );
na02f80 g774883 ( .a(n_6282), .b(n_6203), .o(n_6343) );
no02f80 g778373 ( .a(n_2751), .b(n_2114), .o(n_2947) );
in01f80 g738723 ( .a(n_41399), .o(n_41400) );
no02f80 g777256 ( .a(n_3533), .b(n_3532), .o(n_3534) );
in01f80 FE_OCP_DRV_C1572_n_29860 ( .a(FE_OCP_DRV_N1571_n_29860), .o(FE_OCP_DRV_N1572_n_29860) );
in01f80 FE_OCP_RBC2110_n_6616 ( .a(n_6616), .o(FE_OCP_RBN2110_n_6616) );
na02f80 g765276 ( .a(FE_OCP_RBN2776_n_15110), .b(n_15195), .o(n_15231) );
no02f80 g764152 ( .a(n_16499), .b(n_16446), .o(n_16500) );
in01f80 g738734 ( .a(n_41531), .o(n_41662) );
na02f80 g743766 ( .a(n_37284), .b(n_36824), .o(n_37294) );
ao12f80 g779646 ( .a(n_1570), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n_1790) );
na02f80 g765650 ( .a(n_14911), .b(FE_OCP_RBN2507_n_13896), .o(n_14943) );
in01f80 g753649 ( .a(n_27319), .o(n_27320) );
oa12f80 g747237 ( .a(n_33465), .b(n_33725), .c(n_33462), .o(n_33890) );
in01f80 g740934 ( .a(n_39256), .o(n_39257) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_8_ ( .ck(newNet_1920), .d(n_36896), .o(delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
no02f80 g745241 ( .a(n_35968), .b(n_35892), .o(n_35969) );
na02f80 g740581 ( .a(n_39678), .b(n_39660), .o(n_39691) );
na02f80 g743083 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_6_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .o(n_36935) );
no02f80 g759748 ( .a(n_21600), .b(n_21104), .o(n_21601) );
in01f80 g747389 ( .a(n_32651), .o(n_32652) );
na02f80 FE_RC_1103_0 ( .a(FE_RN_327_0), .b(FE_RN_328_0), .o(FE_RN_329_0) );
na02f80 g781025 ( .a(sin_out_5), .b(FE_OFN3_n_43918), .o(n_311) );
na02f80 FE_RC_1956_0 ( .a(FE_RN_629_0), .b(n_19388), .o(n_19517) );
no02f80 FE_RC_2211_0 ( .a(n_20345), .b(n_20914), .o(FE_RN_797_0) );
in01f80 g767650 ( .a(n_12802), .o(n_12827) );
in01f80 g758964 ( .a(n_21609), .o(n_21636) );
in01f80 newInst_1002 ( .a(newNet_1001), .o(newNet_1002) );
ao22s80 g774769 ( .a(n_6328), .b(n_6226), .c(n_45216), .d(n_6225), .o(n_6379) );
no02f80 g780514 ( .a(n_726), .b(n_751), .o(n_1096) );
na02f80 g750518 ( .a(n_29481), .b(n_29428), .o(n_29482) );
in01f80 g749512 ( .a(n_30575), .o(n_30595) );
in01f80 g768345 ( .a(n_12947), .o(n_12617) );
in01f80 FE_OCP_RBC3500_n_8187 ( .a(FE_OCP_RBN3499_n_8187), .o(FE_OCP_RBN3500_n_8187) );
na02f80 g774608 ( .a(n_6320), .b(FE_OCP_RBN3105_n_6358), .o(n_6404) );
na02f80 g744703 ( .a(n_35198), .b(n_34055), .o(n_35251) );
na02f80 g748505 ( .a(n_31476), .b(n_30803), .o(n_31683) );
no02f80 g748757 ( .a(n_31112), .b(n_27366), .o(n_31202) );
na02f80 g766271 ( .a(n_14245), .b(n_14243), .o(n_14248) );
na02f80 g773019 ( .a(n_7752), .b(n_7672), .o(n_7766) );
no02f80 g767354 ( .a(n_13507), .b(n_13480), .o(n_13549) );
na02f80 g742792 ( .a(n_37344), .b(n_37157), .o(n_37389) );
in01f80 g776207 ( .a(n_4558), .o(n_4530) );
na02f80 g773901 ( .a(n_7007), .b(n_6771), .o(n_7052) );
in01f80 g767852 ( .a(n_13069), .o(n_13317) );
na02f80 g751315 ( .a(n_29597), .b(n_28961), .o(n_29651) );
in01f80 newInst_2077 ( .a(newNet_2076), .o(newNet_2077) );
na02f80 g759572 ( .a(n_20729), .b(n_20687), .o(n_20853) );
no02f80 FE_RC_3665_0 ( .a(n_24848), .b(n_26440), .o(FE_RN_1609_0) );
in01f80 g771491 ( .a(n_9137), .o(n_9138) );
na02f80 FE_RC_3093_0 ( .a(FE_RN_1365_0), .b(FE_RN_1366_0), .o(n_21786) );
ao22s80 g736375 ( .a(n_43772), .b(n_43561), .c(n_43759), .d(n_43560), .o(n_43823) );
in01f80 g745233 ( .a(n_34492), .o(n_34573) );
oa12f80 g753146 ( .a(n_26912), .b(n_26993), .c(n_26837), .o(n_27047) );
in01f80 g740872 ( .a(n_39374), .o(n_39375) );
in01f80 g778517 ( .a(n_2594), .o(n_2595) );
na02f80 g771214 ( .a(n_9884), .b(n_9815), .o(n_9816) );
na02f80 g756568 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_22_), .o(n_23711) );
oa12f80 g748019 ( .a(n_32075), .b(n_31954), .c(n_32077), .o(n_32184) );
in01f80 g739646 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_31_), .o(n_40594) );
in01f80 newInst_433 ( .a(newNet_432), .o(newNet_433) );
no02f80 g777336 ( .a(n_3690), .b(n_3721), .o(n_3883) );
na02f80 g775383 ( .a(n_5537), .b(n_5495), .o(n_5644) );
in01f80 g751960 ( .a(n_29305), .o(n_29306) );
oa12f80 g748781 ( .a(n_30962), .b(n_31241), .c(n_31081), .o(n_31242) );
na02f80 g766631 ( .a(n_13862), .b(n_13842), .o(n_14027) );
in01f80 newInst_3750 ( .a(newNet_1108), .o(newNet_3750) );
na02f80 g766996 ( .a(n_13798), .b(n_13797), .o(n_13799) );
in01f80 FE_OCP_RBC2243_n_13017 ( .a(FE_OCP_RBN2242_n_13017), .o(FE_OCP_RBN2243_n_13017) );
in01f80 g742397 ( .a(n_37775), .o(n_37776) );
na02f80 g762831 ( .a(n_18104), .b(n_17470), .o(n_18123) );
na02f80 g779375 ( .a(n_1552), .b(n_1395), .o(n_1635) );
na02f80 g742826 ( .a(n_37215), .b(n_37130), .o(n_37233) );
in01f80 newInst_924 ( .a(newNet_767), .o(newNet_924) );
na02f80 g765480 ( .a(n_15077), .b(n_14758), .o(n_15195) );
in01f80 newInst_1484 ( .a(newNet_602), .o(newNet_1484) );
na02f80 g771378 ( .a(n_9400), .b(FE_OCP_RBN3546_n_44575), .o(n_9531) );
no02f80 g758688 ( .a(n_21946), .b(n_20275), .o(n_21960) );
in01f80 g746581 ( .a(n_34615), .o(n_34549) );
na02f80 g741939 ( .a(n_38117), .b(n_38115), .o(n_38169) );
in01f80 g775507 ( .a(n_5433), .o(n_5434) );
in01f80 newInst_2924 ( .a(newNet_1082), .o(newNet_2924) );
in01f80 g771695 ( .a(n_9027), .o(n_9070) );
no02f80 g743072 ( .a(n_37090), .b(n_37089), .o(n_37248) );
na02f80 FE_RC_642_0 ( .a(n_28682), .b(FE_RN_203_0), .o(n_28705) );
na02f80 g752953 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_8_), .o(n_27875) );
in01f80 g747966 ( .a(n_32186), .o(n_32187) );
in01f80 newInst_1905 ( .a(newNet_1904), .o(newNet_1905) );
na02f80 g762650 ( .a(n_18038), .b(delay_add_ln22_unr11_stage5_stallmux_q_12_), .o(n_18105) );
in01f80 g777402 ( .a(n_3651), .o(n_3652) );
na02f80 g781303 ( .a(beta_31), .b(beta_5), .o(n_44) );
no02f80 g745266 ( .a(n_35803), .b(FE_OCP_RBN2988_n_35539), .o(n_35892) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_18_ ( .ck(newNet_2200), .d(n_1092), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_) );
no02f80 g765782 ( .a(n_14933), .b(n_14956), .o(n_15009) );
in01f80 g765349 ( .a(n_15374), .o(n_15375) );
in01f80 g755917 ( .a(n_25739), .o(n_25740) );
in01f80 g757562 ( .a(n_22771), .o(n_22772) );
na02f80 g762408 ( .a(n_45002), .b(n_18689), .o(n_18722) );
in01f80 g773132 ( .a(n_7710), .o(n_7711) );
na02f80 g741915 ( .a(n_38145), .b(n_38208), .o(n_38320) );
in01f80 newInst_1335 ( .a(newNet_1334), .o(newNet_1335) );
ao12f80 g777710 ( .a(n_3383), .b(n_3335), .c(n_2913), .o(n_3473) );
in01f80 newInst_1609 ( .a(newNet_521), .o(newNet_1609) );
na02f80 FE_RC_2267_0 ( .a(n_25528), .b(FE_RN_842_0), .o(FE_RN_843_0) );
ao12f80 g778284 ( .a(n_2835), .b(n_2947), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n_2911) );
oa12f80 g780143 ( .a(n_881), .b(n_1139), .c(n_802), .o(n_1160) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_15_ ( .ck(newNet_2114), .d(n_46997), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_) );
in01f80 FE_RC_3077_0 ( .a(n_27361), .o(FE_RN_1356_0) );
in01f80 g765847 ( .a(n_14886), .o(n_14887) );
no02f80 g736726 ( .a(n_43072), .b(n_43027), .o(n_43073) );
in01f80 g761388 ( .a(n_19678), .o(n_19679) );
oa22f80 g737865 ( .a(n_42270), .b(n_42160), .c(n_42547), .d(n_42151), .o(n_42708) );
ao12f80 g768321 ( .a(n_12487), .b(n_12486), .c(n_12485), .o(n_13073) );
no02f80 g738577 ( .a(n_41688), .b(n_41722), .o(n_42023) );
ao12f80 g738183 ( .a(n_41863), .b(n_41973), .c(n_41694), .o(n_42011) );
na02f80 g773983 ( .a(n_6874), .b(n_5103), .o(n_6992) );
in01f80 FE_OCP_RBC1157_n_18375 ( .a(FE_OCP_RBN1155_n_18375), .o(FE_OCP_RBN1157_n_18375) );
na02f80 g764451 ( .a(n_16630), .b(n_15964), .o(n_16655) );
na02f80 FE_RC_2611_0 ( .a(FE_OCP_RBN3247_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .o(FE_RN_1086_0) );
no02f80 g759692 ( .a(n_20591), .b(n_20611), .o(n_20719) );
in01f80 newInst_2075 ( .a(newNet_2074), .o(newNet_2075) );
oa12f80 g752021 ( .a(n_28694), .b(n_28693), .c(n_28692), .o(n_29026) );
na02f80 FE_RC_2898_0 ( .a(FE_RN_1255_0), .b(n_9633), .o(n_9921) );
no02f80 g771163 ( .a(n_9491), .b(n_9462), .o(n_9621) );
in01f80 newInst_2674 ( .a(newNet_2673), .o(newNet_2674) );
no02f80 g751901 ( .a(n_29004), .b(n_28957), .o(n_29510) );
na02f80 g770960 ( .a(n_10040), .b(n_8428), .o(n_10127) );
na02f80 FE_RC_1071_0 ( .a(FE_RN_315_0), .b(FE_RN_316_0), .o(FE_RN_317_0) );
na02f80 g768738 ( .a(n_12130), .b(n_12042), .o(n_12204) );
in01f80 g752343 ( .a(n_27910), .o(n_28163) );
in01f80 g769063 ( .a(n_11769), .o(n_11718) );
na02f80 g766690 ( .a(n_13849), .b(n_12798), .o(n_13945) );
na02f80 g749962 ( .a(n_29925), .b(n_29863), .o(n_30151) );
no02f80 g742492 ( .a(n_37578), .b(n_37709), .o(n_37645) );
in01f80 g744715 ( .a(n_35231), .o(n_35232) );
ao22s80 g779451 ( .a(n_1373), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n_1438) );
oa12f80 g743934 ( .a(n_35647), .b(n_35646), .c(n_35645), .o(n_35705) );
in01f80 newInst_2049 ( .a(newNet_2048), .o(newNet_2049) );
in01f80 g766198 ( .a(n_14450), .o(n_14484) );
oa12f80 g749323 ( .a(n_30673), .b(n_30672), .c(n_30671), .o(n_30734) );
in01f80 g769960 ( .a(n_11024), .o(n_11025) );
in01f80 g736589 ( .a(n_43627), .o(n_43628) );
in01f80 newInst_1196 ( .a(newNet_1195), .o(newNet_1196) );
no02f80 g748187 ( .a(n_31607), .b(FE_OCP_RBN3714_n_31466), .o(n_31687) );
na02f80 g754743 ( .a(n_26231), .b(n_25687), .o(n_26415) );
na02f80 g771061 ( .a(n_9419), .b(n_8362), .o(n_9422) );
no02f80 g779124 ( .a(n_1940), .b(n_2343), .o(n_1963) );
na02f80 g772322 ( .a(n_8619), .b(FE_OCPN1011_n_7802), .o(n_8663) );
in01f80 g743333 ( .a(n_36753), .o(n_36754) );
na02f80 g777306 ( .a(n_3562), .b(n_3580), .o(n_3581) );
in01f80 g745882 ( .a(n_35354), .o(n_35408) );
in01f80 newInst_3033 ( .a(newNet_880), .o(newNet_3033) );
in01f80 g756517 ( .a(n_24050), .o(n_24051) );
na02f80 g737678 ( .a(n_42392), .b(n_42069), .o(n_42519) );
in01f80 newInst_1575 ( .a(newNet_1574), .o(newNet_1575) );
in01f80 g771707 ( .a(n_9306), .o(n_9307) );
no02f80 g766111 ( .a(n_14539), .b(n_13514), .o(n_14581) );
in01f80 FE_RC_3941_0 ( .a(n_16972), .o(FE_RN_1705_0) );
no02f80 g756171 ( .a(n_24176), .b(n_24098), .o(n_24201) );
na02f80 g751034 ( .a(n_29853), .b(n_186), .o(n_29855) );
no02f80 g776409 ( .a(n_4324), .b(n_4293), .o(n_4458) );
na02f80 g752919 ( .a(n_27733), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .o(n_27790) );
in01f80 g738508 ( .a(n_41632), .o(n_41585) );
no02f80 g780214 ( .a(n_1089), .b(n_883), .o(n_1125) );
no02f80 g778359 ( .a(n_2462), .b(n_2475), .o(n_2517) );
no02f80 g736413 ( .a(n_43791), .b(n_43678), .o(n_43834) );
na02f80 g779401 ( .a(n_1590), .b(n_1549), .o(n_1550) );
na02f80 g745701 ( .a(n_35435), .b(n_35434), .o(n_35436) );
na02f80 FE_RC_3987_0 ( .a(n_29903), .b(n_29815), .o(n_30056) );
in01f80 g768997 ( .a(n_11767), .o(n_11768) );
in01f80 g773068 ( .a(n_8014), .o(n_8015) );
no02f80 g739284 ( .a(n_40771), .b(n_40723), .o(n_40772) );
ao22s80 FE_RC_761_0 ( .a(n_8764), .b(FE_OCPN1011_n_7802), .c(FE_OCP_RBN3467_n_7886), .d(n_8765), .o(n_8879) );
in01f80 newInst_2181 ( .a(newNet_419), .o(newNet_2181) );
na02f80 g749501 ( .a(n_30410), .b(n_30429), .o(n_30465) );
na02f80 g771960 ( .a(n_44463), .b(n_9631), .o(n_9730) );
in01f80 newInst_2737 ( .a(newNet_1905), .o(newNet_2737) );
no02f80 g748411 ( .a(FE_OCP_RBN3088_FE_OCPN1052_n_31674), .b(FE_OCP_RBN2807_n_30643), .o(n_32149) );
no02f80 g742001 ( .a(n_37979), .b(n_37896), .o(n_38125) );
no02f80 g772398 ( .a(n_8517), .b(n_8550), .o(n_8613) );
na02f80 g763667 ( .a(n_16891), .b(FE_OCP_RBN3209_n_44365), .o(n_16892) );
in01f80 g750841 ( .a(n_29228), .o(n_29229) );
no02f80 g758802 ( .a(n_21550), .b(n_21505), .o(n_21955) );
in01f80 g756312 ( .a(n_24079), .o(n_24117) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_24_ ( .ck(newNet_3519), .d(n_22789), .o(delay_add_ln22_unr14_stage6_stallmux_q_24_) );
na02f80 g764809 ( .a(n_15625), .b(n_15192), .o(n_15739) );
no02f80 g756941 ( .a(n_24169), .b(n_23779), .o(n_24240) );
na02f80 g770743 ( .a(n_10100), .b(FE_OCPN3771_n_8669), .o(n_10145) );
in01f80 g739583 ( .a(n_40617), .o(n_40619) );
oa22f80 FE_RC_945_0 ( .a(n_22801), .b(FE_OCP_RBN3116_n_22710), .c(n_22833), .d(n_22710), .o(n_22802) );
oa12f80 g775696 ( .a(n_5414), .b(n_5432), .c(n_5413), .o(n_5498) );
ao12f80 g761509 ( .a(n_19647), .b(n_19793), .c(n_19291), .o(n_19820) );
na02f80 g772858 ( .a(n_8051), .b(n_8050), .o(n_8158) );
in01f80 g747445 ( .a(n_32525), .o(n_32432) );
na02f80 g772902 ( .a(n_7843), .b(n_7720), .o(n_7948) );
no02f80 g753595 ( .a(n_26753), .b(n_26752), .o(n_26774) );
no02f80 g778597 ( .a(n_2609), .b(n_2620), .o(n_2621) );
in01f80 g754487 ( .a(n_25545), .o(n_25568) );
no02f80 g777870 ( .a(n_3120), .b(n_2451), .o(n_3166) );
na02f80 g744883 ( .a(n_34996), .b(FE_OCPN1434_n_30614), .o(n_35033) );
no02f80 g772814 ( .a(n_8100), .b(n_8099), .o(n_8123) );
in01f80 g743184 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_6_), .o(n_36946) );
in01f80 g741255 ( .a(n_39267), .o(n_39268) );
in01f80 FE_OCP_RBC1330_n_18866 ( .a(FE_OCP_RBN1329_n_18866), .o(FE_OCP_RBN1330_n_18866) );
in01f80 newInst_1118 ( .a(newNet_938), .o(newNet_1118) );
na02f80 g760740 ( .a(n_20201), .b(n_20200), .o(n_20202) );
na02f80 g773138 ( .a(FE_OCP_RBN3461_n_7886), .b(n_7945), .o(n_8018) );
na02f80 g742026 ( .a(n_38010), .b(n_37943), .o(n_38011) );
na02f80 g754971 ( .a(n_25148), .b(n_25241), .o(n_25463) );
na02f80 g760575 ( .a(n_20329), .b(n_20328), .o(n_20330) );
na02f80 g759791 ( .a(n_21824), .b(n_21693), .o(n_21859) );
no02f80 g767778 ( .a(n_12777), .b(n_12766), .o(n_12862) );
no02f80 g739459 ( .a(n_44800), .b(n_40454), .o(n_40816) );
in01f80 g777685 ( .a(n_3334), .o(n_3372) );
no02f80 g757294 ( .a(n_44084), .b(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .o(n_23023) );
in01f80 g754580 ( .a(n_26233), .o(n_26930) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_18_ ( .ck(newNet_3235), .d(n_36455), .o(delay_add_ln22_unr23_stage9_stallmux_q_18_) );
na02f80 g745200 ( .a(n_35648), .b(FE_OCP_DRV_N1592_n_34327), .o(n_34629) );
oa22f80 g744583 ( .a(n_36599), .b(n_36155), .c(n_36600), .d(n_36156), .o(n_36666) );
oa12f80 g739041 ( .a(n_41113), .b(n_41112), .c(n_41111), .o(n_41156) );
oa22f80 FE_RC_3380_0 ( .a(n_21645), .b(n_21927), .c(n_21678), .d(n_21895), .o(n_21983) );
in01f80 g777315 ( .a(n_3756), .o(n_3757) );
na02f80 g776499 ( .a(n_4322), .b(n_4393), .o(n_4441) );
in01f80 FE_RC_4198_0 ( .a(n_19184), .o(n_19178) );
na02f80 g762419 ( .a(n_45120), .b(n_18064), .o(n_18535) );
ao12f80 g749898 ( .a(FE_OCP_RBN3010_n_31117), .b(n_31275), .c(n_31213), .o(n_31346) );
no02f80 g745451 ( .a(n_34649), .b(n_34704), .o(n_34705) );
oa12f80 g747592 ( .a(n_31681), .b(n_32223), .c(n_32197), .o(n_32225) );
in01f80 g776124 ( .a(FE_OCP_RBN2840_n_4692), .o(n_5940) );
no02f80 g747096 ( .a(n_32794), .b(n_32793), .o(n_32800) );
no02f80 g737897 ( .a(n_42202), .b(n_41911), .o(n_42247) );
na03f80 FE_RC_3419_0 ( .a(n_27026), .b(FE_RN_1356_0), .c(n_27194), .o(FE_RN_1357_0) );
ao22s80 FE_RC_1596_0 ( .a(n_45319), .b(FE_OCP_RBN3687_n_5105), .c(n_5105), .d(n_45318), .o(n_5284) );
oa12f80 g781158 ( .a(n_190), .b(n_189), .c(n_188), .o(n_516) );
no02f80 g764280 ( .a(n_16207), .b(n_16234), .o(n_16337) );
in01f80 g777676 ( .a(n_3481), .o(n_3482) );
in01f80 g759238 ( .a(n_20945), .o(n_20946) );
in01f80 g746026 ( .a(n_35243), .o(n_35218) );
in01f80 g758401 ( .a(FE_OCPN1488_n_23447), .o(n_23509) );
no02f80 g765091 ( .a(n_15492), .b(n_15491), .o(n_15493) );
oa22f80 g752647 ( .a(n_27473), .b(n_27546), .c(n_27442), .d(n_27547), .o(n_27576) );
ao22s80 g745210 ( .a(n_34573), .b(n_34378), .c(n_34518), .d(n_34379), .o(n_35521) );
no02f80 g736641 ( .a(n_43035), .b(n_43075), .o(n_43156) );
in01f80 g761080 ( .a(n_19207), .o(n_19208) );
in01f80 FE_OCP_RBC2224_n_12902 ( .a(n_12902), .o(FE_OCP_RBN2224_n_12902) );
no02f80 g771657 ( .a(n_8851), .b(n_8669), .o(n_8938) );
no02f80 g763036 ( .a(n_17489), .b(n_17488), .o(n_17490) );
na02f80 g772941 ( .a(n_7847), .b(n_7844), .o(n_7939) );
na02f80 g775923 ( .a(n_5218), .b(n_4647), .o(n_5279) );
in01f80 g747513 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .o(n_32542) );
in01f80 g767897 ( .a(n_13168), .o(n_13271) );
no02f80 g762694 ( .a(n_17996), .b(n_17995), .o(n_18016) );
ao12f80 g779437 ( .a(n_1764), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .o(n_1829) );
no03m80 g746389 ( .a(FE_OCP_RBN2178_n_33022), .b(n_33433), .c(n_32972), .o(n_33525) );
oa12f80 g770714 ( .a(n_10204), .b(n_10334), .c(n_10125), .o(n_10425) );
na02f80 g748901 ( .a(n_32356), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(n_32423) );
oa22f80 FE_RC_953_0 ( .a(n_32131), .b(n_32346), .c(n_32130), .d(n_32330), .o(n_32471) );
na02f80 g757574 ( .a(n_22602), .b(n_22474), .o(n_22682) );
no02f80 FE_RC_2170_0 ( .a(n_26555), .b(FE_OCP_RBN2910_n_26394), .o(FE_RN_772_0) );
ao12f80 g741531 ( .a(n_38690), .b(n_45623), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38719) );
in01f80 g748452 ( .a(n_31765), .o(n_31783) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_10_ ( .ck(newNet_197), .d(n_46366), .o(delay_xor_ln22_unr9_stage4_stallmux_q_10_) );
oa12f80 g767630 ( .a(n_12939), .b(n_12938), .c(n_12937), .o(n_13787) );
no02f80 g778329 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_29_), .o(n_2920) );
in01f80 FE_OCP_RBC3856_FE_RN_779_0 ( .a(FE_RN_779_0), .o(FE_OCP_RBN3856_FE_RN_779_0) );
no02f80 g740388 ( .a(FE_OCP_RBN3028_n_39942), .b(n_39889), .o(n_40245) );
no02f80 g768373 ( .a(n_12443), .b(n_12442), .o(n_12444) );
na02f80 g765846 ( .a(n_15212), .b(n_14492), .o(n_15287) );
oa22f80 FE_RC_3801_0 ( .a(n_38778), .b(n_38654), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .d(n_38628), .o(n_38673) );
no02f80 FE_RC_2459_0 ( .a(n_13904), .b(n_13895), .o(FE_RN_986_0) );
na02f80 g750916 ( .a(n_28976), .b(n_28600), .o(n_29020) );
no02f80 g752761 ( .a(n_27437), .b(n_27276), .o(n_27438) );
in01f80 FE_OCP_RBC3337_n_44610 ( .a(n_44610), .o(FE_OCP_RBN3337_n_44610) );
na02f80 FE_RC_1726_0 ( .a(n_23373), .b(n_23374), .o(FE_RN_477_0) );
in01f80 g769715 ( .a(n_11271), .o(n_11272) );
in01f80 FE_OCP_RBC1714_n_20734 ( .a(n_20734), .o(FE_OCP_RBN1714_n_20734) );
no02f80 g743971 ( .a(n_47266), .b(n_47264), .o(n_36009) );
in01f80 newInst_339 ( .a(newNet_68), .o(newNet_339) );
na02f80 g749131 ( .a(n_30958), .b(n_27246), .o(n_31050) );
in01f80 g747320 ( .a(n_32706), .o(n_32712) );
no02f80 g757191 ( .a(n_23210), .b(n_23039), .o(n_23231) );
no02f80 g755298 ( .a(n_24971), .b(n_24964), .o(n_24970) );
na02f80 g740664 ( .a(n_39476), .b(n_39503), .o(n_39556) );
in01f80 g776874 ( .a(FE_OCP_RBN2626_n_3848), .o(n_3922) );
no02f80 g757869 ( .a(n_22237), .b(n_22063), .o(n_22389) );
in01f80 newInst_3749 ( .a(newNet_3748), .o(newNet_3749) );
na02f80 g754084 ( .a(n_26014), .b(n_26059), .o(n_26103) );
ao22s80 g780357 ( .a(n_1079), .b(FE_OFN761_n_45813), .c(n_853), .d(n_1203), .o(n_949) );
in01f80 g771630 ( .a(n_8817), .o(n_8796) );
in01f80 FE_OCP_RBC1715_n_20734 ( .a(n_20734), .o(FE_OCP_RBN1715_n_20734) );
na02f80 g769841 ( .a(n_11162), .b(n_11016), .o(n_11189) );
na02f80 g736874 ( .a(n_43453), .b(n_43092), .o(n_43536) );
no02f80 g753907 ( .a(n_26389), .b(n_26281), .o(n_26421) );
in01f80 g744541 ( .a(n_35399), .o(n_35400) );
no02f80 g766647 ( .a(n_13918), .b(FE_OCP_RBN2243_n_13017), .o(n_13947) );
in01f80 g756063 ( .a(n_25119), .o(n_25120) );
no02f80 g741594 ( .a(n_38633), .b(n_38778), .o(n_38650) );
no02f80 g768311 ( .a(n_12530), .b(delay_add_ln22_unr8_stage4_stallmux_q_15_), .o(n_12549) );
in01f80 FE_OCP_RBC2531_n_38693 ( .a(n_38693), .o(FE_OCP_RBN2531_n_38693) );
no02f80 g750179 ( .a(n_29810), .b(n_29848), .o(n_29811) );
in01f80 g759339 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_2_), .o(n_22941) );
oa22f80 FE_RC_3398_0 ( .a(n_24350), .b(n_27835), .c(n_27796), .d(FE_OCP_RBN1220_n_27835), .o(n_27894) );
na02f80 FE_RC_2296_0 ( .a(FE_RN_864_0), .b(n_44827), .o(n_28634) );
no02f80 g751702 ( .a(n_28368), .b(n_28367), .o(n_28389) );
na02f80 g747485 ( .a(n_33446), .b(n_33363), .o(n_33746) );
na02f80 g760974 ( .a(n_19355), .b(n_19354), .o(n_19422) );
in01f80 newInst_3634 ( .a(newNet_2637), .o(newNet_3634) );
oa22f80 g769662 ( .a(n_11288), .b(n_10381), .c(n_11287), .d(n_10382), .o(n_11344) );
na02f80 g741245 ( .a(FE_OCP_RBN2637_n_38806), .b(n_38527), .o(n_38984) );
in01f80 newInst_1430 ( .a(newNet_962), .o(newNet_1430) );
ao22s80 FE_RC_1365_0 ( .a(n_5172), .b(n_5129), .c(n_5171), .d(n_5128), .o(n_5307) );
in01f80 newInst_1745 ( .a(newNet_1683), .o(newNet_1745) );
no02f80 g762173 ( .a(n_18814), .b(n_18618), .o(n_18884) );
na02f80 FE_RC_2068_0 ( .a(n_35059), .b(FE_RN_703_0), .o(n_35078) );
no02f80 g769675 ( .a(n_11229), .b(n_11230), .o(n_11258) );
na02f80 g757927 ( .a(n_22852), .b(n_22652), .o(n_22853) );
in01f80 g761180 ( .a(n_19062), .o(n_19063) );
na02f80 g758807 ( .a(n_21784), .b(n_21842), .o(n_21869) );
ao12f80 g748579 ( .a(n_31300), .b(n_31270), .c(n_31272), .o(n_31426) );
no02f80 g741209 ( .a(n_39033), .b(n_39032), .o(n_39034) );
no02f80 g777970 ( .a(n_3090), .b(n_3089), .o(n_3091) );
no02f80 g737775 ( .a(n_42283), .b(n_41955), .o(n_42284) );
no02f80 g780489 ( .a(n_925), .b(n_913), .o(n_926) );
in01f80 FE_OCP_RBC2439_n_8402 ( .a(FE_OCP_RBN2438_n_8402), .o(FE_OCP_RBN2439_n_8402) );
na02f80 g755395 ( .a(n_25573), .b(n_25572), .o(n_25574) );
na02f80 g754290 ( .a(n_25924), .b(n_25911), .o(n_26037) );
na02f80 g742902 ( .a(n_37008), .b(n_37006), .o(n_37009) );
na02f80 g743297 ( .a(n_37922), .b(n_46247), .o(n_37923) );
no02f80 g775285 ( .a(n_5555), .b(n_4875), .o(n_5574) );
na02f80 g759414 ( .a(n_20771), .b(n_45066), .o(n_20825) );
oa12f80 g760409 ( .a(n_20027), .b(n_20079), .c(n_19859), .o(n_20127) );
na02f80 g756804 ( .a(n_23377), .b(n_23376), .o(n_23427) );
na02f80 g770050 ( .a(n_10856), .b(n_10456), .o(n_10909) );
no02f80 g775780 ( .a(n_5508), .b(FE_OCP_RBN2647_n_47014), .o(n_5626) );
na02f80 g775448 ( .a(n_5524), .b(n_5568), .o(n_5587) );
in01f80 g750260 ( .a(n_29839), .o(n_29840) );
no02f80 g741133 ( .a(n_39318), .b(n_38942), .o(n_39433) );
no02f80 g750597 ( .a(n_30192), .b(FE_OFN788_n_25834), .o(n_29424) );
oa12f80 g761895 ( .a(n_18970), .b(n_18969), .c(n_18968), .o(n_19650) );
in01f80 g756263 ( .a(n_24157), .o(n_24173) );
oa22f80 FE_RC_3168_0 ( .a(n_17336), .b(n_17686), .c(n_16338), .d(n_44153), .o(n_17755) );
na02f80 g743024 ( .a(n_37210), .b(n_37106), .o(n_37107) );
in01f80 g739764 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n_40471) );
na02f80 g773706 ( .a(n_7335), .b(n_7085), .o(n_7336) );
na02f80 g763852 ( .a(n_16702), .b(FE_OCP_RBN2675_n_14991), .o(n_16726) );
in01f80 FE_OCP_RBC3119_n_22755 ( .a(n_22755), .o(FE_OCP_RBN3119_n_22755) );
ao12f80 g738907 ( .a(n_41268), .b(n_41267), .c(n_41266), .o(n_41695) );
oa22f80 FE_RC_196_0 ( .a(n_17320), .b(n_17522), .c(n_17319), .d(n_17566), .o(n_17697) );
in01f80 g739898 ( .a(n_40377), .o(n_40378) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_29_ ( .ck(newNet_3204), .d(n_36651), .o(delay_add_ln22_unr23_stage9_stallmux_q_29_) );
ao12f80 g778390 ( .a(n_2751), .b(n_2684), .c(n_2683), .o(n_2796) );
no02f80 g776417 ( .a(n_4405), .b(n_4385), .o(n_4445) );
in01f80 g764640 ( .a(n_15915), .o(n_16007) );
in01f80 g742787 ( .a(n_37393), .o(n_37364) );
no02f80 g765266 ( .a(n_15521), .b(n_15520), .o(n_15522) );
no02f80 g740890 ( .a(n_39369), .b(n_39297), .o(n_39429) );
na02f80 g781345 ( .a(n_7), .b(beta_11), .o(n_127) );
na02f80 g756231 ( .a(n_24057), .b(n_23661), .o(n_24083) );
in01f80 newInst_2828 ( .a(newNet_2827), .o(newNet_2828) );
na02f80 g771436 ( .a(n_9190), .b(n_9012), .o(n_9318) );
in01f80 g742778 ( .a(n_37409), .o(n_37365) );
no02f80 g744104 ( .a(n_36064), .b(n_44180), .o(n_36141) );
no02f80 FE_RC_1881_0 ( .a(n_11919), .b(FE_RN_584_0), .o(n_11772) );
in01f80 newInst_689 ( .a(newNet_688), .o(newNet_689) );
no02f80 g768769 ( .a(n_11925), .b(n_11654), .o(n_11987) );
na02f80 g765479 ( .a(FE_OCP_RBN2736_n_14985), .b(FE_OCPN1007_n_13962), .o(n_15052) );
in01f80 g758391 ( .a(n_23509), .o(n_23486) );
na02f80 g753959 ( .a(n_26188), .b(FE_OCPN1440_n_23339), .o(n_26218) );
oa12f80 g756883 ( .a(n_23803), .b(n_24088), .c(n_24087), .o(n_24090) );
ao22s80 FE_RC_2672_0 ( .a(n_3015), .b(n_3935), .c(n_3014), .d(n_3859), .o(n_4158) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_2_ ( .ck(newNet_1293), .d(n_729), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_) );
na02f80 g738194 ( .a(n_41962), .b(n_41978), .o(n_41979) );
no02f80 g754711 ( .a(FE_OCP_RBN2955_n_26231), .b(n_25712), .o(n_26549) );
no02f80 g773855 ( .a(n_7127), .b(n_7126), .o(n_7128) );
no02f80 g763376 ( .a(FE_OCPN1756_n_16923), .b(n_15479), .o(n_17391) );
in01f80 FE_OCP_RBC3338_n_44610 ( .a(n_44610), .o(FE_OCP_RBN3338_n_44610) );
ao12f80 g745277 ( .a(n_34272), .b(n_34326), .c(n_34245), .o(n_34465) );
no02f80 g741499 ( .a(n_38747), .b(n_38736), .o(n_38737) );
in01f80 newInst_1289 ( .a(newNet_906), .o(newNet_1289) );
in01f80 newInst_1718 ( .a(newNet_1717), .o(newNet_1718) );
no02f80 g737488 ( .a(n_42635), .b(n_42645), .o(n_42685) );
oa22f80 FE_RC_3912_0 ( .a(n_36236), .b(n_36517), .c(n_36237), .d(n_36516), .o(n_36615) );
in01f80 g762190 ( .a(n_18240), .o(n_18241) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_10_ ( .ck(newNet_1548), .d(n_31976), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_) );
oa12f80 g762002 ( .a(n_18355), .b(n_18461), .c(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n_18508) );
ao12f80 g751201 ( .a(n_29128), .b(n_29771), .c(n_29124), .o(n_29805) );
na02f80 g740887 ( .a(n_39396), .b(n_39428), .o(n_40183) );
na02f80 g737928 ( .a(n_42202), .b(n_42035), .o(n_42302) );
no02f80 g762916 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_20_), .b(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n_17568) );
in01f80 g776795 ( .a(n_4248), .o(n_4249) );
in01f80 g760229 ( .a(n_20395), .o(n_20396) );
na02f80 FE_RC_1835_0 ( .a(n_13913), .b(FE_RN_552_0), .o(FE_RN_553_0) );
na02f80 g738135 ( .a(n_42040), .b(n_42028), .o(n_42107) );
na02f80 g775629 ( .a(n_47001), .b(n_5603), .o(n_5710) );
no02f80 g767814 ( .a(n_13118), .b(n_12914), .o(n_13160) );
oa22f80 g739825 ( .a(n_40347), .b(n_40327), .c(n_40348), .d(n_40326), .o(n_40421) );
in01f80 newInst_2012 ( .a(newNet_2011), .o(newNet_2012) );
na02f80 g747132 ( .a(n_33953), .b(n_33464), .o(n_33995) );
no02f80 g774500 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_), .o(n_6641) );
na02f80 g752134 ( .a(n_46961), .b(delay_add_ln22_unr17_stage7_stallmux_q_3_), .o(n_28142) );
in01f80 FE_OCP_RBC1680_n_33491 ( .a(n_33491), .o(FE_OCP_RBN1680_n_33491) );
na02f80 g771849 ( .a(n_44516), .b(n_10078), .o(n_10158) );
na02f80 g779281 ( .a(n_1762), .b(n_1789), .o(n_1763) );
no02f80 g773413 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .o(n_7669) );
in01f80 g755812 ( .a(n_24443), .o(n_24444) );
na02f80 g746919 ( .a(n_33108), .b(n_32303), .o(n_33198) );
in01f80 g744915 ( .a(n_35980), .o(n_35006) );
in01f80 g741677 ( .a(FE_OCP_RBN3504_n_38592), .o(n_39095) );
ao12f80 g740777 ( .a(n_39511), .b(n_39510), .c(n_39509), .o(n_39561) );
in01f80 newInst_3259 ( .a(newNet_300), .o(newNet_3259) );
no02f80 g745525 ( .a(n_34353), .b(n_34324), .o(n_34378) );
in01f80 g780349 ( .a(n_899), .o(n_973) );
na02f80 g740436 ( .a(n_39787), .b(n_39471), .o(n_39914) );
oa22f80 FE_RC_3516_0 ( .a(FE_OCPN1017_n_23307), .b(FE_RN_555_0), .c(FE_RN_557_0), .d(FE_RN_556_0), .o(n_23363) );
oa22f80 g777952 ( .a(n_3163), .b(n_3178), .c(n_3218), .d(n_3217), .o(n_3248) );
in01f80 FE_RC_3218_0 ( .a(n_11747), .o(FE_RN_1429_0) );
ao12f80 g780684 ( .a(n_656), .b(n_657), .c(n_655), .o(n_660) );
ao22s80 g759140 ( .a(n_21014), .b(n_20711), .c(n_21015), .d(n_20710), .o(n_21163) );
in01f80 g777587 ( .a(n_3564), .o(n_3562) );
no02f80 g755171 ( .a(n_25023), .b(n_25022), .o(n_25046) );
in01f80 g737592 ( .a(n_42524), .o(n_42525) );
in01f80 g757248 ( .a(n_23492), .o(n_23493) );
in01f80 g741343 ( .a(n_38828), .o(n_39032) );
in01f80 g766376 ( .a(n_14318), .o(n_14319) );
in01f80 fopt782887 ( .a(n_26407), .o(n_44325) );
in01f80 g764779 ( .a(n_15736), .o(n_15737) );
na02f80 g766002 ( .a(n_14667), .b(n_14695), .o(n_14798) );
na02f80 g750850 ( .a(n_29056), .b(FE_OFN788_n_25834), .o(n_29115) );
na02f80 g742710 ( .a(n_37326), .b(n_37325), .o(n_37327) );
in01f80 newInst_1840 ( .a(newNet_1839), .o(newNet_1840) );
in01f80 g750446 ( .a(n_29604), .o(n_29605) );
in01f80 FE_OCP_RBC3849_n_20290 ( .a(n_20290), .o(FE_OCP_RBN3849_n_20290) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_14_ ( .ck(newNet_362), .d(n_1348), .o(delay_xor_ln22_unr3_stage2_stallmux_q_14_) );
na02f80 g777626 ( .a(n_3586), .b(n_3540), .o(n_3613) );
na02f80 g748316 ( .a(n_31553), .b(n_30757), .o(n_31558) );
na02f80 g763279 ( .a(n_17194), .b(n_17193), .o(n_17231) );
na02f80 g759765 ( .a(n_21447), .b(n_21519), .o(n_21518) );
no02f80 g774015 ( .a(n_6802), .b(n_6610), .o(n_6800) );
ao12f80 g771899 ( .a(FE_OCP_RBN2493_n_8508), .b(FE_OCP_RBN2517_n_8762), .c(n_8561), .o(n_8836) );
in01f80 g758824 ( .a(n_21794), .o(n_21733) );
na02f80 g745410 ( .a(FE_OCP_RBN2984_n_35539), .b(n_35583), .o(n_35584) );
no02f80 g776351 ( .a(n_4465), .b(n_4543), .o(n_4560) );
in01f80 g758117 ( .a(n_22098), .o(n_22129) );
in01f80 g779386 ( .a(n_1577), .o(n_1578) );
in01f80 g774983 ( .a(n_6243), .o(n_6217) );
in01f80 FE_RC_3931_0 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .o(FE_RN_1700_0) );
no02f80 g778931 ( .a(n_2151), .b(n_1841), .o(n_2168) );
in01f80 g757101 ( .a(n_23142), .o(n_23143) );
na02f80 g748286 ( .a(FE_OCP_RBN3732_n_31819), .b(n_31034), .o(n_32015) );
no02f80 g755479 ( .a(n_24694), .b(n_22484), .o(n_24695) );
na02f80 g777696 ( .a(n_3503), .b(FE_OCP_RBN2382_n_3502), .o(n_3568) );
in01f80 g737163 ( .a(n_43097), .o(n_43230) );
in01f80 newInst_906 ( .a(newNet_838), .o(newNet_906) );
no02f80 g768890 ( .a(n_11726), .b(n_11661), .o(n_11736) );
na02f80 FE_RC_2419_0 ( .a(n_7165), .b(FE_RN_956_0), .o(n_7534) );
ao12f80 g758130 ( .a(n_22844), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n_23152) );
no02f80 g770373 ( .a(n_10659), .b(n_10637), .o(n_10638) );
na02f80 g756997 ( .a(n_23346), .b(n_23213), .o(n_23367) );
na02f80 g765069 ( .a(n_15383), .b(n_15422), .o(n_15644) );
ao12f80 g757679 ( .a(n_22291), .b(FE_OCPN3184_n_22294), .c(n_44322), .o(n_22743) );
in01f80 g772821 ( .a(n_8042), .o(n_8074) );
na02f80 g750422 ( .a(n_29620), .b(n_29494), .o(n_29642) );
in01f80 g737261 ( .a(n_42927), .o(n_42938) );
oa22f80 FE_RC_796_0 ( .a(n_8452), .b(n_8657), .c(FE_OCP_RBN2442_n_8402), .d(FE_OCP_RBN2516_n_8657), .o(n_8776) );
na02f80 g768578 ( .a(n_12233), .b(n_11900), .o(n_12236) );
na02f80 g766169 ( .a(n_14547), .b(FE_OCP_RBN3533_n_13765), .o(n_14549) );
in01f80 g759702 ( .a(n_21752), .o(n_21753) );
in01f80 g769092 ( .a(n_11638), .o(n_11639) );
no02f80 g749795 ( .a(n_31311), .b(n_31372), .o(n_31408) );
in01f80 g737706 ( .a(n_42420), .o(n_42437) );
ao12f80 g741945 ( .a(n_38063), .b(FE_OCP_RBN2256_n_37844), .c(n_37982), .o(n_38064) );
na03f80 FE_RC_2587_0 ( .a(FE_RN_1067_0), .b(FE_RN_1068_0), .c(n_17827), .o(FE_RN_1069_0) );
na02f80 g781072 ( .a(sin_out_24), .b(FE_OFN4_n_43918), .o(n_296) );
in01f80 newInst_2249 ( .a(newNet_2248), .o(newNet_2249) );
no02f80 g748892 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n_32445) );
oa22f80 FE_RC_3822_0 ( .a(n_15453), .b(n_15858), .c(n_15454), .d(n_15815), .o(n_16053) );
in01f80 newInst_3468 ( .a(newNet_3467), .o(newNet_3468) );
in01f80 newInst_2023 ( .a(newNet_2022), .o(newNet_2023) );
no02f80 g744738 ( .a(n_35102), .b(n_30614), .o(n_35152) );
in01f80 g739912 ( .a(n_40124), .o(n_40199) );
na02f80 g776370 ( .a(n_4661), .b(n_4267), .o(n_4664) );
no02f80 g748389 ( .a(n_31518), .b(n_30553), .o(n_31664) );
in01f80 FE_RC_495_0 ( .a(n_28229), .o(FE_RN_147_0) );
na02f80 g742976 ( .a(n_37082), .b(n_36503), .o(n_37133) );
in01f80 FE_OCP_RBC1355_n_44259 ( .a(n_44259), .o(FE_OCP_RBN1355_n_44259) );
in01f80 g781297 ( .a(n_62), .o(n_111) );
no02f80 g779623 ( .a(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .o(n_1705) );
na02f80 g776757 ( .a(n_3830), .b(n_2791), .o(n_3872) );
na02f80 g771472 ( .a(n_9519), .b(n_8024), .o(n_9603) );
in01f80 FE_OCPC1518_n_26752 ( .a(FE_OCPN1517_n_26752), .o(FE_OCPN1518_n_26752) );
in01f80 newInst_1688 ( .a(newNet_1687), .o(newNet_1688) );
ao22s80 FE_RC_3866_0 ( .a(FE_OCP_RBN3220_n_21358), .b(n_22288), .c(FE_OCP_RBN3219_n_21358), .d(FE_OCPN991_n_22249), .o(FE_RN_1689_0) );
ms00f80 sin_out_reg_6_ ( .ck(newNet_17), .d(n_43677), .o(sin_out_6) );
oa22f80 g749630 ( .a(n_30204), .b(n_30015), .c(n_30250), .d(n_30014), .o(n_31740) );
no02f80 FE_RC_4187_0 ( .a(FE_RN_1834_0), .b(n_24389), .o(FE_RN_1833_0) );
in01f80 g747667 ( .a(n_33760), .o(n_33761) );
no02f80 g740245 ( .a(n_39882), .b(n_39939), .o(n_39996) );
oa22f80 FE_RC_3249_0 ( .a(n_10757), .b(n_10790), .c(n_10789), .d(n_10758), .o(n_10906) );
na02f80 g746895 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_22_), .o(n_33199) );
oa12f80 g747769 ( .a(n_33600), .b(n_33571), .c(n_33554), .o(n_34021) );
no02f80 g752508 ( .a(n_28339), .b(n_28338), .o(n_28340) );
in01f80 fopt783587 ( .a(n_6328), .o(n_45216) );
na02f80 g766871 ( .a(n_14385), .b(n_14390), .o(n_14349) );
na02f80 g768307 ( .a(n_12579), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .o(n_12621) );
no02f80 g757093 ( .a(n_23248), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .o(n_23264) );
ao12f80 g772715 ( .a(n_8193), .b(n_8192), .c(n_8204), .o(n_9906) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_22_ ( .ck(newNet_1735), .d(n_22522), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_) );
oa12f80 g781091 ( .a(n_250), .b(n_258), .c(n_249), .o(n_437) );
na02f80 g774109 ( .a(FE_OCP_RBN2128_n_6745), .b(n_6547), .o(n_6729) );
in01f80 g769664 ( .a(n_11356), .o(n_11334) );
in01f80 newInst_3732 ( .a(newNet_3731), .o(newNet_3732) );
in01f80 fopt783655 ( .a(n_45301), .o(n_45300) );
in01f80 g743105 ( .a(n_37046), .o(n_37047) );
no02f80 g738243 ( .a(n_41928), .b(n_41927), .o(n_41929) );
in01f80 g753555 ( .a(n_27451), .o(n_27452) );
oa12f80 g780097 ( .a(n_725), .b(n_1119), .c(n_751), .o(n_1153) );
no02f80 g757905 ( .a(n_22313), .b(FE_OCPN3787_n_22156), .o(n_22353) );
no02f80 g764365 ( .a(n_16201), .b(n_16168), .o(n_16324) );
oa12f80 g759818 ( .a(n_21598), .b(FE_OCP_RBN3678_n_21051), .c(n_21597), .o(n_21722) );
no02f80 g751485 ( .a(n_28801), .b(n_28800), .o(n_28826) );
oa12f80 g746305 ( .a(n_33205), .b(n_33475), .c(n_33474), .o(n_33508) );
oa12f80 g776009 ( .a(n_5054), .b(n_5107), .c(n_5053), .o(n_5244) );
no02f80 g763146 ( .a(n_17348), .b(n_17347), .o(n_17406) );
no02f80 g754551 ( .a(n_26308), .b(n_26348), .o(n_26349) );
in01f80 newInst_83 ( .a(newNet_82), .o(newNet_83) );
in01f80 g769609 ( .a(n_11426), .o(n_11427) );
in01f80 g762983 ( .a(n_17594), .o(n_17565) );
no02f80 g748164 ( .a(n_47272), .b(n_47271), .o(n_32134) );
in01f80 g760297 ( .a(n_20281), .o(n_20282) );
na02f80 g740798 ( .a(n_39470), .b(n_40202), .o(n_39471) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_17_ ( .ck(newNet_2205), .d(n_1040), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_) );
in01f80 g747609 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n_32348) );
in01f80 g741123 ( .a(n_38991), .o(n_38992) );
na02f80 g745730 ( .a(n_34428), .b(n_34429), .o(n_34430) );
no02f80 g777232 ( .a(n_3417), .b(n_3424), .o(n_3557) );
no02f80 g763749 ( .a(n_46978), .b(FE_OCP_RBN2735_n_14985), .o(n_16762) );
in01f80 g771951 ( .a(n_9206), .o(n_9207) );
no02f80 g755056 ( .a(n_25647), .b(n_25535), .o(n_25536) );
oa12f80 g772754 ( .a(n_7360), .b(n_8042), .c(n_7307), .o(n_8106) );
in01f80 g751085 ( .a(n_30288), .o(n_30289) );
in01f80 newInst_568 ( .a(newNet_567), .o(newNet_568) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_7_ ( .ck(newNet_544), .d(n_17337), .o(delay_xor_ln22_unr12_stage5_stallmux_q_7_) );
in01f80 newInst_1295 ( .a(newNet_1294), .o(newNet_1295) );
in01f80 g770569 ( .a(n_10277), .o(n_10314) );
oa22f80 g778971 ( .a(n_2186), .b(n_1961), .c(n_2201), .d(n_1960), .o(n_2246) );
oa12f80 g765073 ( .a(n_16348), .b(n_16347), .c(n_16346), .o(n_16410) );
na02f80 g761785 ( .a(n_19158), .b(n_18884), .o(n_19293) );
na02f80 g760885 ( .a(n_19431), .b(n_17881), .o(n_19528) );
na02f80 g755872 ( .a(n_25306), .b(n_25166), .o(n_26072) );
in01f80 g757611 ( .a(FE_OCPN1780_n_24097), .o(n_22752) );
no02f80 g743820 ( .a(n_35878), .b(n_34918), .o(n_35879) );
no02f80 g736823 ( .a(n_43223), .b(n_43216), .o(n_43261) );
na02f80 g738208 ( .a(n_41977), .b(n_41963), .o(n_41964) );
in01f80 FE_OCP_RBC2639_n_38806 ( .a(FE_OCP_RBN2636_n_38806), .o(FE_OCP_RBN2639_n_38806) );
na02f80 g779186 ( .a(n_2494), .b(n_1909), .o(n_1910) );
in01f80 g752107 ( .a(n_28793), .o(n_28836) );
oa22f80 g781126 ( .a(n_219), .b(n_114), .c(n_220), .d(n_113), .o(n_402) );
na02f80 g770503 ( .a(n_10319), .b(n_10332), .o(n_10402) );
in01f80 newInst_1267 ( .a(newNet_1266), .o(newNet_1267) );
in01f80 g755130 ( .a(n_25500), .o(n_25556) );
in01f80 FE_OCPC3748_n_34296 ( .a(n_34296), .o(FE_OCPN3748_n_34296) );
in01f80 newInst_634 ( .a(newNet_633), .o(newNet_634) );
na02f80 g780085 ( .a(n_1198), .b(n_1195), .o(n_1196) );
in01f80 newInst_975 ( .a(newNet_974), .o(newNet_975) );
na02f80 g738383 ( .a(n_41513), .b(n_41472), .o(n_41514) );
na02f80 g773516 ( .a(n_7507), .b(n_7116), .o(n_7508) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_15_ ( .ck(newNet_2966), .d(n_6047), .o(delay_add_ln22_unr5_stage3_stallmux_q_15_) );
na02f80 g761063 ( .a(n_19117), .b(n_18427), .o(n_19183) );
no02f80 g777998 ( .a(n_3067), .b(n_2558), .o(n_3123) );
ao12f80 g743204 ( .a(n_36751), .b(n_36894), .c(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36896) );
ao12f80 g779449 ( .a(n_2026), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .o(n_2070) );
in01f80 g743061 ( .a(n_37142), .o(n_37143) );
na02f80 g776431 ( .a(n_4538), .b(n_4254), .o(n_4539) );
na02f80 g752987 ( .a(n_27274), .b(n_27187), .o(n_27275) );
in01f80 g766390 ( .a(n_14133), .o(n_14199) );
in01f80 fopt784012 ( .a(n_30263), .o(n_45744) );
in01f80 g755214 ( .a(n_25201), .o(n_25374) );
oa22f80 FE_RC_1692_0 ( .a(n_30401), .b(n_30886), .c(n_30402), .d(n_30885), .o(n_31010) );
na02f80 g756859 ( .a(n_23379), .b(n_23178), .o(n_23362) );
in01f80 FE_OCPC1025_n_25481 ( .a(n_25481), .o(FE_OCPN1025_n_25481) );
no02f80 g755530 ( .a(n_24528), .b(n_22111), .o(n_24580) );
na02f80 g753724 ( .a(n_26531), .b(n_26530), .o(n_26764) );
in01f80 newInst_1731 ( .a(newNet_1730), .o(newNet_1731) );
no02f80 g764740 ( .a(n_15700), .b(n_14524), .o(n_15741) );
na02f80 g777731 ( .a(FE_OCP_RBN2488_n_3338), .b(n_2913), .o(n_3359) );
ao12f80 g738959 ( .a(n_41060), .b(n_41155), .c(n_41208), .o(n_41222) );
in01f80 FE_OFC818_n_4575 ( .a(FE_OFN836_n_4575), .o(FE_OFN818_n_4575) );
na02f80 g740131 ( .a(n_39816), .b(n_39371), .o(n_39846) );
no02f80 g770737 ( .a(n_10146), .b(FE_OFN755_n_44461), .o(n_10190) );
na02f80 g780873 ( .a(n_457), .b(n_495), .o(n_515) );
in01f80 g761744 ( .a(n_18822), .o(n_18998) );
no02f80 g742249 ( .a(n_37864), .b(n_37863), .o(n_37865) );
na02f80 g776718 ( .a(n_3993), .b(n_3872), .o(n_4080) );
in01f80 g769232 ( .a(n_11675), .o(n_11676) );
in01f80 FE_OCPC1495_n_26528 ( .a(n_26528), .o(FE_OCPN1495_n_26528) );
no02f80 g776987 ( .a(n_3852), .b(FE_OCP_RBN2649_n_3840), .o(n_3979) );
na02f80 g748356 ( .a(n_31721), .b(n_31757), .o(n_31827) );
in01f80 newInst_1067 ( .a(newNet_971), .o(newNet_1067) );
na02f80 g739799 ( .a(n_40470), .b(n_40225), .o(n_40484) );
no02f80 g771295 ( .a(n_9513), .b(n_8185), .o(n_9555) );
in01f80 g757013 ( .a(n_24045), .o(n_24086) );
in01f80 g756280 ( .a(n_24072), .o(n_24043) );
no02f80 g737079 ( .a(n_43120), .b(n_43004), .o(n_43383) );
na02f80 g768651 ( .a(n_12253), .b(n_12252), .o(n_12377) );
in01f80 fopt784288 ( .a(n_7), .o(n_46055) );
na02f80 g749773 ( .a(n_31339), .b(n_31289), .o(n_31369) );
no02f80 g738398 ( .a(n_41580), .b(n_41640), .o(n_41641) );
in01f80 newInst_2712 ( .a(newNet_1077), .o(newNet_2712) );
ao12f80 g774060 ( .a(n_6834), .b(n_6833), .c(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n_6949) );
na02f80 g769268 ( .a(n_11556), .b(n_10802), .o(n_11752) );
na02f80 g762973 ( .a(n_17981), .b(n_17980), .o(n_17982) );
in01f80 FE_OCP_RBC3104_n_40561 ( .a(n_40561), .o(FE_OCP_RBN3104_n_40561) );
in01f80 newInst_1363 ( .a(newNet_1362), .o(newNet_1363) );
in01f80 newInst_1229 ( .a(newNet_1228), .o(newNet_1229) );
na03f80 FE_RC_1095_0 ( .a(n_17930), .b(FE_RN_323_0), .c(n_17827), .o(n_17971) );
na02f80 g746889 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_20_), .o(n_33097) );
ao12f80 g773037 ( .a(n_8118), .b(n_8362), .c(n_8150), .o(n_8961) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_9_ ( .ck(newNet_283), .d(n_1294), .o(delay_xor_ln22_unr3_stage2_stallmux_q_9_) );
in01f80 g774440 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .o(n_6512) );
no02f80 FE_RC_1742_0 ( .a(FE_RN_488_0), .b(n_12418), .o(n_12413) );
na02f80 g739035 ( .a(n_41073), .b(n_40757), .o(n_41098) );
na02f80 FE_RC_2702_0 ( .a(FE_RN_1134_0), .b(FE_RN_1133_0), .o(FE_RN_1135_0) );
ao12f80 g761817 ( .a(n_18398), .b(n_18406), .c(n_18284), .o(n_18516) );
in01f80 g749089 ( .a(n_30987), .o(n_30988) );
in01f80 g756523 ( .a(n_24009), .o(n_24010) );
no02f80 g777290 ( .a(n_4606), .b(FE_OFN821_n_4632), .o(n_5548) );
na02f80 g774805 ( .a(n_45474), .b(n_5609), .o(n_6326) );
in01f80 newInst_1105 ( .a(newNet_1104), .o(newNet_1105) );
in01f80 newInst_804 ( .a(newNet_803), .o(newNet_804) );
ms00f80 cos_out_reg_12_ ( .ck(newNet_3749), .d(n_43776), .o(cos_out_12) );
na02f80 g740356 ( .a(n_39739), .b(n_39738), .o(n_39771) );
in01f80 g745110 ( .a(n_34786), .o(n_34822) );
ao12f80 g771170 ( .a(n_9532), .b(n_9720), .c(n_9586), .o(n_9761) );
in01f80 g758452 ( .a(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .o(n_23259) );
no02f80 FE_RC_2241_0 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(FE_RN_819_0), .o(FE_RN_820_0) );
no02f80 g765871 ( .a(n_15128), .b(n_14486), .o(n_15212) );
ao12f80 g777750 ( .a(n_3455), .b(n_3454), .c(n_3453), .o(n_4777) );
in01f80 newInst_1568 ( .a(newNet_1567), .o(newNet_1568) );
in01f80 g765890 ( .a(n_14877), .o(n_14899) );
ao22s80 g742727 ( .a(n_37409), .b(n_37179), .c(n_37365), .d(n_37178), .o(n_38279) );
in01f80 FE_RC_2083_0 ( .a(n_27062), .o(FE_RN_713_0) );
no02f80 g779846 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .o(n_1632) );
na02f80 g755490 ( .a(n_24577), .b(n_23360), .o(n_24698) );
na02f80 g771853 ( .a(n_9283), .b(n_9380), .o(n_9435) );
in01f80 g744902 ( .a(n_36463), .o(n_36450) );
no02f80 g775393 ( .a(n_5526), .b(n_5529), .o(n_5554) );
no02f80 g748876 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .o(n_32418) );
in01f80 FE_OCP_RBC2112_n_22650 ( .a(n_22650), .o(FE_OCP_RBN2112_n_22650) );
no02f80 g741585 ( .a(n_38617), .b(n_38631), .o(n_38680) );
oa12f80 g738278 ( .a(n_41502), .b(n_41865), .c(n_41807), .o(n_41894) );
na02f80 FE_RC_4144_0 ( .a(n_16900), .b(n_16936), .o(FE_RN_1800_0) );
no02f80 g741147 ( .a(n_38981), .b(n_38568), .o(n_39039) );
na02f80 g769308 ( .a(n_11440), .b(n_10623), .o(n_11664) );
no02f80 g770999 ( .a(n_9928), .b(n_9763), .o(n_9963) );
na02f80 g769211 ( .a(n_11548), .b(n_11590), .o(n_11834) );
in01f80 g737362 ( .a(n_42847), .o(n_42862) );
in01f80 g745547 ( .a(n_34375), .o(n_34436) );
na03f80 g743313 ( .a(n_36855), .b(n_37855), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_37897) );
in01f80 newInst_2178 ( .a(newNet_2177), .o(newNet_2178) );
in01f80 FE_OCP_RBC2457_n_13765 ( .a(n_13765), .o(FE_OCP_RBN2457_n_13765) );
no02f80 g773969 ( .a(n_6937), .b(n_6651), .o(n_6960) );
na02f80 g742200 ( .a(n_44877), .b(n_37869), .o(n_37972) );
na02f80 g777815 ( .a(n_3206), .b(n_2386), .o(n_3318) );
in01f80 newInst_262 ( .a(newNet_261), .o(newNet_262) );
ao22s80 g773849 ( .a(n_7073), .b(n_6929), .c(FE_OCP_RBN3379_n_7073), .d(n_6928), .o(n_7129) );
na02f80 g769790 ( .a(n_11195), .b(n_11228), .o(n_11236) );
na02f80 g765156 ( .a(n_15413), .b(n_15412), .o(n_15414) );
na02f80 g767356 ( .a(n_13435), .b(FE_OCPN1472_n_13434), .o(n_13500) );
na02f80 g758167 ( .a(n_21973), .b(FE_OCP_RBN3853_n_20848), .o(n_22083) );
no02f80 g777184 ( .a(n_3769), .b(n_3883), .o(n_3984) );
ao12f80 g747892 ( .a(n_33120), .b(n_33119), .c(n_33118), .o(n_33651) );
no02f80 g775913 ( .a(n_4960), .b(n_4182), .o(n_5087) );
in01f80 g753277 ( .a(n_27294), .o(n_27395) );
no02f80 g754354 ( .a(n_25765), .b(n_25791), .o(n_25874) );
no02f80 g744239 ( .a(n_46220), .b(n_36808), .o(n_37381) );
in01f80 FE_OCP_RBC2932_n_5307 ( .a(n_5307), .o(FE_OCP_RBN2932_n_5307) );
in01f80 newInst_285 ( .a(newNet_284), .o(newNet_285) );
in01f80 g777228 ( .a(n_3899), .o(n_3900) );
in01f80 newInst_98 ( .a(newNet_97), .o(newNet_98) );
na02f80 g780569 ( .a(n_713), .b(n_734), .o(n_742) );
no02f80 g756615 ( .a(n_23606), .b(n_23653), .o(n_23738) );
in01f80 g758658 ( .a(n_21898), .o(n_21913) );
no02f80 g756003 ( .a(n_25160), .b(n_25000), .o(n_25436) );
na02f80 g752004 ( .a(n_28897), .b(n_28555), .o(n_29285) );
oa22f80 g775700 ( .a(n_5365), .b(n_4160), .c(n_5335), .d(n_5529), .o(n_5499) );
in01f80 g760852 ( .a(n_19470), .o(n_19471) );
in01f80 g737138 ( .a(n_43082), .o(n_43228) );
ao12f80 g763543 ( .a(n_16667), .b(n_16690), .c(n_16708), .o(n_16793) );
in01f80 g759945 ( .a(n_21772), .o(n_21773) );
na02f80 g777354 ( .a(FE_OCP_RBN2583_n_3734), .b(n_3771), .o(n_3940) );
oa22f80 FE_RC_1623_0 ( .a(n_17336), .b(n_17759), .c(n_17753), .d(n_44334), .o(n_17832) );
no02f80 g738539 ( .a(n_41379), .b(n_41388), .o(n_41431) );
no02f80 g762274 ( .a(n_18723), .b(n_18769), .o(n_19295) );
oa22f80 g757858 ( .a(n_22239), .b(n_22018), .c(n_22238), .d(n_22019), .o(n_22425) );
in01f80 newInst_1995 ( .a(newNet_1994), .o(newNet_1995) );
na02f80 g760835 ( .a(n_20265), .b(n_18140), .o(n_19583) );
in01f80 g780050 ( .a(n_1242), .o(n_1243) );
na02f80 g764783 ( .a(FE_OCP_RBN2777_n_15595), .b(n_14524), .o(n_15658) );
na02f80 g763243 ( .a(n_17273), .b(n_17393), .o(n_17473) );
oa12f80 g738868 ( .a(n_41232), .b(n_41231), .c(n_41230), .o(n_41481) );
in01f80 g737940 ( .a(n_42294), .o(n_42295) );
in01f80 g780019 ( .a(n_1266), .o(n_1270) );
ao12f80 g767615 ( .a(n_12479), .b(n_12713), .c(n_12506), .o(n_12805) );
in01f80 g775375 ( .a(n_5754), .o(n_5780) );
in01f80 newInst_3060 ( .a(newNet_3059), .o(newNet_3060) );
ao12f80 g745981 ( .a(n_35247), .b(n_35246), .c(n_35245), .o(n_35720) );
in01f80 FE_OCP_RBC2893_n_26152 ( .a(n_26152), .o(FE_OCP_RBN2893_n_26152) );
in01f80 g773918 ( .a(n_6941), .o(n_6916) );
in01f80 g780989 ( .a(n_357), .o(n_374) );
in01f80 g758486 ( .a(FE_OFN735_n_22641), .o(n_23115) );
in01f80 g777368 ( .a(n_3725), .o(n_3726) );
in01f80 g736907 ( .a(n_43634), .o(n_43635) );
oa22f80 g757229 ( .a(n_44218), .b(n_23206), .c(n_44219), .d(n_23207), .o(n_24502) );
na02f80 FE_RC_4169_0 ( .a(n_18333), .b(FE_RN_1817_0), .o(FE_RN_1818_0) );
na02f80 g736717 ( .a(n_43053), .b(n_43046), .o(n_43093) );
in01f80 g756484 ( .a(n_23967), .o(n_23968) );
no02f80 g771465 ( .a(n_8847), .b(n_7737), .o(n_8921) );
na02f80 g771360 ( .a(n_9253), .b(n_9318), .o(n_9408) );
in01f80 g765030 ( .a(n_15387), .o(n_15472) );
in01f80 FE_OCP_RBC2846_n_30678 ( .a(n_30678), .o(FE_OCP_RBN2846_n_30678) );
na02f80 g775419 ( .a(n_5824), .b(n_5823), .o(n_5825) );
no02f80 g766640 ( .a(n_13857), .b(n_13319), .o(n_13924) );
na02f80 FE_RC_2919_0 ( .a(FE_RN_1270_0), .b(n_24404), .o(n_24471) );
no02f80 g775709 ( .a(n_5539), .b(n_5072), .o(n_5545) );
na02f80 g741032 ( .a(n_38836), .b(n_38820), .o(n_38837) );
no02f80 g779382 ( .a(n_1513), .b(n_1437), .o(n_1524) );
in01f80 g737467 ( .a(n_42652), .o(n_42669) );
in01f80 g774818 ( .a(n_6308), .o(n_6309) );
in01f80 g761718 ( .a(n_19526), .o(n_19540) );
oa12f80 g772643 ( .a(n_8246), .b(n_8255), .c(n_8245), .o(n_10028) );
in01f80 g766447 ( .a(n_14099), .o(n_14120) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_24_ ( .ck(newNet_3410), .d(n_27793), .o(delay_add_ln22_unr17_stage7_stallmux_q_24_) );
no02f80 g778522 ( .a(n_2608), .b(n_2083), .o(n_2614) );
no02f80 g744845 ( .a(FE_OCP_RBN2614_n_35005), .b(FE_OCPN1796_n_30546), .o(n_35061) );
in01f80 g738480 ( .a(n_41410), .o(n_41411) );
na02f80 g753947 ( .a(n_26190), .b(n_23353), .o(n_26301) );
no02f80 g752300 ( .a(n_27936), .b(n_27889), .o(n_27962) );
na02f80 g745611 ( .a(n_34369), .b(n_34504), .o(n_34532) );
no02f80 g776027 ( .a(n_4915), .b(FE_OCPN846_n_4046), .o(n_4978) );
na02f80 g755699 ( .a(n_24488), .b(n_24457), .o(n_24552) );
in01f80 FE_OFC829_n_2405 ( .a(n_2405), .o(FE_OFN829_n_2405) );
in01f80 newInst_3386 ( .a(newNet_3385), .o(newNet_3386) );
in01f80 newInst_3173 ( .a(newNet_3172), .o(newNet_3173) );
na02f80 g755743 ( .a(n_24445), .b(n_23852), .o(n_24500) );
ao12f80 g779138 ( .a(n_1994), .b(n_1993), .c(n_1992), .o(n_2038) );
in01f80 g755501 ( .a(n_24687), .o(n_24688) );
oa12f80 g761052 ( .a(n_19310), .b(n_19309), .c(n_19308), .o(n_19407) );
in01f80 FE_OCPC3771_n_8669 ( .a(FE_OCPN3770_n_8669), .o(FE_OCPN3771_n_8669) );
in01f80 g757031 ( .a(n_23955), .o(n_23904) );
na02f80 g759469 ( .a(n_21029), .b(n_21028), .o(n_21055) );
in01f80 g746212 ( .a(n_33772), .o(n_33804) );
in01f80 g748919 ( .a(n_32450), .o(n_32406) );
in01f80 FE_OCPC871_n_2737 ( .a(FE_OCPN870_n_2737), .o(FE_OCPN871_n_2737) );
no02f80 g761314 ( .a(n_19828), .b(n_19792), .o(n_19829) );
oa12f80 g746338 ( .a(n_35044), .b(n_35043), .c(n_35042), .o(n_35631) );
no02f80 g740187 ( .a(FE_OCP_RBN3717_n_39913), .b(n_39599), .o(n_40135) );
no02f80 g774110 ( .a(n_6669), .b(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n_6691) );
in01f80 g740766 ( .a(n_39450), .o(n_39387) );
na02f80 g759106 ( .a(n_21348), .b(n_21222), .o(n_21421) );
na02f80 g752926 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .o(n_28156) );
na02f80 g761922 ( .a(n_18268), .b(n_18367), .o(n_18440) );
in01f80 newInst_1809 ( .a(newNet_1808), .o(newNet_1809) );
oa22f80 g768407 ( .a(n_12373), .b(n_12165), .c(n_12418), .d(n_12166), .o(n_12909) );
in01f80 g775937 ( .a(n_4776), .o(n_4849) );
oa22f80 g749171 ( .a(n_32116), .b(n_31627), .c(n_32154), .d(n_31628), .o(n_32228) );
na02f80 FE_RC_3981_0 ( .a(FE_RN_1725_0), .b(n_29697), .o(n_29730) );
na02f80 g783841 ( .a(n_45525), .b(FE_RN_846_0), .o(n_45527) );
na02f80 g756403 ( .a(n_23825), .b(n_23741), .o(n_23946) );
no02f80 g763182 ( .a(n_17341), .b(n_17342), .o(n_17507) );
na02f80 FE_RC_3540_0 ( .a(n_19025), .b(FE_RN_1532_0), .o(FE_RN_1533_0) );
ao22s80 g742586 ( .a(n_37460), .b(n_37061), .c(n_37459), .d(n_37062), .o(n_37965) );
in01f80 FE_OFC345_n_9247 ( .a(FE_OCP_RBN2677_n_9247), .o(FE_OFN345_n_9247) );
na02f80 g744639 ( .a(n_35211), .b(FE_OCP_RBN2684_n_35213), .o(n_35274) );
oa22f80 g779875 ( .a(n_44652), .b(n_1165), .c(n_44661), .d(n_1143), .o(n_1295) );
na03f80 FE_RC_3777_0 ( .a(n_34144), .b(n_34187), .c(n_34146), .o(n_34188) );
no02f80 g755732 ( .a(n_25142), .b(n_25091), .o(n_25171) );
no02f80 g743884 ( .a(n_35872), .b(n_35751), .o(n_35873) );
no02f80 g740055 ( .a(n_40042), .b(n_40041), .o(n_40076) );
na02f80 g775434 ( .a(n_5348), .b(n_5127), .o(n_5417) );
in01f80 FE_OCPC1432_n_29504 ( .a(FE_OCPN1431_n_29504), .o(FE_OCPN1432_n_29504) );
na02f80 g776005 ( .a(n_5164), .b(n_5176), .o(n_5321) );
no02f80 g744691 ( .a(n_35287), .b(FE_OCPN1794_n_30612), .o(n_35326) );
in01f80 g766509 ( .a(n_14117), .o(n_14181) );
no02f80 g763819 ( .a(n_17572), .b(n_17497), .o(n_18211) );
ao12f80 g771102 ( .a(n_9402), .b(n_9502), .c(n_9486), .o(n_9637) );
no02f80 g746721 ( .a(n_33145), .b(n_33110), .o(n_33111) );
oa12f80 g774979 ( .a(n_5965), .b(n_6041), .c(n_5923), .o(n_6100) );
in01f80 FE_OCP_RBC3686_n_16074 ( .a(n_16074), .o(FE_OCP_RBN3686_n_16074) );
in01f80 g750318 ( .a(n_29751), .o(n_29752) );
no02f80 g771869 ( .a(n_9207), .b(n_9322), .o(n_9429) );
na02f80 g771488 ( .a(n_9339), .b(n_9241), .o(n_9485) );
na02f80 g754117 ( .a(n_26091), .b(FE_OCPN1530_n_26090), .o(n_26092) );
no02f80 g751001 ( .a(n_30207), .b(n_30097), .o(n_30254) );
na02f80 g774745 ( .a(n_6414), .b(n_6265), .o(n_6438) );
in01f80 FE_RC_1189_0 ( .a(n_13017), .o(FE_RN_360_0) );
na02f80 g744767 ( .a(n_35150), .b(n_35174), .o(n_35269) );
in01f80 g755245 ( .a(n_25640), .o(n_25714) );
in01f80 newInst_1846 ( .a(newNet_61), .o(newNet_1846) );
na02f80 g781328 ( .a(n_7), .b(beta_21), .o(n_84) );
in01f80 g769334 ( .a(n_11525), .o(n_11606) );
no02f80 g763757 ( .a(n_16777), .b(n_16715), .o(n_16753) );
in01f80 g746426 ( .a(n_34294), .o(n_33385) );
oa12f80 g738836 ( .a(n_41289), .b(n_41288), .c(n_41287), .o(n_41654) );
na02f80 g747630 ( .a(n_32298), .b(n_32105), .o(n_32360) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_21_ ( .ck(newNet_2652), .d(n_22684), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_) );
na02f80 g773896 ( .a(n_7058), .b(n_7060), .o(n_7059) );
in01f80 g772987 ( .a(n_8091), .o(n_8055) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_0_ ( .ck(newNet_1550), .d(n_186), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_) );
oa22f80 g784566 ( .a(FE_OFN800_n_46285), .b(n_10783), .c(FE_OCP_RBN3709_n_46337), .d(n_10716), .o(n_46387) );
na02f80 g737736 ( .a(n_42285), .b(n_41984), .o(n_42451) );
na02f80 g740446 ( .a(n_39727), .b(n_39674), .o(n_39728) );
no02f80 g765151 ( .a(n_15457), .b(n_15379), .o(n_15527) );
in01f80 g777364 ( .a(n_4833), .o(n_4834) );
na02f80 g759913 ( .a(n_20608), .b(n_20538), .o(n_20713) );
na02f80 g769974 ( .a(n_11017), .b(FE_OCP_RBN2720_n_9494), .o(n_11107) );
no02f80 FE_RC_2053_0 ( .a(n_27121), .b(n_25963), .o(FE_RN_694_0) );
in01f80 FE_RC_3848_0 ( .a(FE_OCPN1741_n_19138), .o(FE_RN_1679_0) );
no02f80 g762883 ( .a(n_18013), .b(n_17463), .o(n_18084) );
no02f80 g755026 ( .a(n_25117), .b(n_25106), .o(n_25181) );
no02f80 g760416 ( .a(n_20065), .b(n_19942), .o(n_20100) );
no02f80 g750071 ( .a(n_29869), .b(n_29296), .o(n_30577) );
oa22f80 g741101 ( .a(FE_OCP_RBN3624_n_38870), .b(n_38543), .c(FE_OCPN957_n_39096), .d(n_38564), .o(n_39528) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_12_ ( .ck(newNet_463), .d(n_27844), .o(delay_xor_ln22_unr18_stage7_stallmux_q_12_) );
na02f80 FE_RC_3999_0 ( .a(n_29969), .b(n_30178), .o(FE_RN_1735_0) );
na02f80 g761147 ( .a(n_19075), .b(n_19045), .o(n_19114) );
no02f80 g780783 ( .a(n_519), .b(n_518), .o(n_520) );
na02f80 g769810 ( .a(n_11052), .b(FE_OCP_RBN3643_n_44490), .o(n_11123) );
no02f80 g745289 ( .a(n_35938), .b(n_35937), .o(n_35966) );
no02f80 g744910 ( .a(n_34935), .b(n_34957), .o(n_35063) );
na02f80 g742667 ( .a(n_37370), .b(n_37143), .o(n_37418) );
oa12f80 g780319 ( .a(n_945), .b(n_889), .c(n_870), .o(n_963) );
in01f80 newInst_1547 ( .a(newNet_1546), .o(newNet_1547) );
na02f80 g750068 ( .a(n_29896), .b(n_29327), .o(n_30196) );
na02f80 g763195 ( .a(n_17473), .b(n_17472), .o(n_17474) );
na02f80 g756573 ( .a(n_23561), .b(n_23560), .o(n_23584) );
no02f80 g765280 ( .a(n_15829), .b(n_15826), .o(n_16023) );
no02f80 g762247 ( .a(n_18496), .b(n_18694), .o(n_18663) );
ao12f80 g741975 ( .a(n_37833), .b(n_37917), .c(n_37866), .o(n_37991) );
in01f80 g750032 ( .a(n_30970), .o(n_30971) );
in01f80 FE_OCP_RBC1691_n_19052 ( .a(n_19052), .o(FE_OCP_RBN1691_n_19052) );
no02f80 g751974 ( .a(n_28836), .b(n_28879), .o(n_28943) );
na02f80 g756175 ( .a(n_24200), .b(n_23858), .o(n_24224) );
in01f80 FE_OFC753_n_44461 ( .a(FE_OCP_RBN2616_n_44561), .o(FE_OFN753_n_44461) );
in01f80 g770071 ( .a(n_10831), .o(n_10832) );
in01f80 g765110 ( .a(n_16133), .o(n_16134) );
ao12f80 g775608 ( .a(n_5201), .b(n_45484), .c(n_5177), .o(n_5389) );
in01f80 g752945 ( .a(n_27787), .o(n_27788) );
no02f80 g745427 ( .a(FE_OCP_RBN2993_n_35539), .b(n_35675), .o(n_35715) );
na02f80 g767915 ( .a(n_12843), .b(n_12783), .o(n_12873) );
no02f80 g780530 ( .a(n_659), .b(n_423), .o(n_707) );
na02f80 g762881 ( .a(n_17865), .b(n_17864), .o(n_17909) );
na02f80 g775309 ( .a(n_46998), .b(FE_OCP_RBN2842_n_4784), .o(n_6002) );
in01f80 g753328 ( .a(n_27071), .o(n_27072) );
oa22f80 g751874 ( .a(n_28066), .b(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .c(n_28070), .d(n_44735), .o(n_28381) );
oa12f80 g743879 ( .a(n_35711), .b(n_35710), .c(n_35709), .o(n_35791) );
in01f80 newInst_73 ( .a(newNet_72), .o(newNet_73) );
no02f80 g769175 ( .a(FE_OCP_RBN2111_n_11548), .b(n_11606), .o(n_11637) );
no02f80 g759404 ( .a(n_20735), .b(n_20583), .o(n_20776) );
oa22f80 g742869 ( .a(n_37113), .b(n_36919), .c(n_37187), .d(n_36920), .o(n_37770) );
na02f80 g741106 ( .a(n_39001), .b(n_38999), .o(n_39133) );
oa12f80 g770631 ( .a(n_9735), .b(n_10373), .c(n_9649), .o(n_10422) );
no02f80 g758121 ( .a(n_44268), .b(n_21242), .o(n_22342) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_23_ ( .ck(newNet_1986), .d(n_11778), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_) );
ao12f80 g772612 ( .a(n_7447), .b(n_8101), .c(n_7472), .o(n_8186) );
in01f80 g757717 ( .a(n_22613), .o(n_22675) );
na02f80 g742898 ( .a(n_36935), .b(n_36964), .o(n_37013) );
na02f80 g764416 ( .a(n_16095), .b(n_14618), .o(n_16205) );
na02f80 g738756 ( .a(n_41525), .b(n_41264), .o(n_41598) );
in01f80 FE_OCP_RBC2105_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(FE_OCP_RBN2004_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN2105_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
no02f80 g763938 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n_17530) );
in01f80 newInst_1348 ( .a(newNet_86), .o(newNet_1348) );
in01f80 g760819 ( .a(n_19558), .o(n_19559) );
na02f80 g760635 ( .a(n_19729), .b(n_19708), .o(n_19806) );
oa12f80 g750805 ( .a(n_30336), .b(n_30335), .c(n_30334), .o(n_31116) );
in01f80 g758147 ( .a(n_22046), .o(n_22344) );
oa22f80 FE_RC_1450_0 ( .a(n_22907), .b(n_22901), .c(n_22833), .d(n_22861), .o(n_22960) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_10_ ( .ck(newNet_3350), .d(n_31670), .o(delay_add_ln22_unr20_stage8_stallmux_q_10_) );
in01f80 newInst_1099 ( .a(newNet_525), .o(newNet_1099) );
in01f80 newInst_2525 ( .a(newNet_2524), .o(newNet_2525) );
na02f80 g736655 ( .a(n_43474), .b(n_43230), .o(n_43563) );
in01f80 g774498 ( .a(n_6561), .o(n_6562) );
oa12f80 g745279 ( .a(n_35561), .b(n_35605), .c(FE_OFN221_n_35655), .o(n_36222) );
na02f80 g736778 ( .a(n_43254), .b(n_43251), .o(n_43269) );
no02f80 g780805 ( .a(n_514), .b(n_536), .o(n_655) );
in01f80 g780510 ( .a(n_999), .o(n_1000) );
no02f80 g756037 ( .a(n_24902), .b(n_23837), .o(n_24954) );
in01f80 g738547 ( .a(n_41735), .o(n_41621) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_20_ ( .ck(newNet_2950), .d(n_6267), .o(delay_add_ln22_unr5_stage3_stallmux_q_20_) );
na03f80 g741062 ( .a(n_39068), .b(n_39131), .c(n_39130), .o(n_39278) );
in01f80 g749562 ( .a(n_30573), .o(n_30593) );
no02f80 g747310 ( .a(n_32818), .b(n_32666), .o(n_32729) );
oa12f80 g768096 ( .a(n_12398), .b(n_12569), .c(n_12353), .o(n_12615) );
in01f80 g773649 ( .a(n_47176), .o(n_7377) );
no02f80 g741177 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39230), .o(n_39242) );
oa22f80 g757819 ( .a(n_22392), .b(n_20231), .c(n_22355), .d(n_22580), .o(n_22449) );
na02f80 g737782 ( .a(n_42414), .b(n_42302), .o(n_42408) );
no02f80 g746031 ( .a(n_33959), .b(n_33958), .o(n_34032) );
no02f80 g779298 ( .a(FE_OCP_RBN3380_n_1732), .b(n_1503), .o(n_1813) );
in01f80 newInst_306 ( .a(newNet_225), .o(newNet_306) );
in01f80 g736393 ( .a(n_43775), .o(n_43814) );
in01f80 FE_RC_2654_0 ( .a(n_12590), .o(FE_RN_1108_0) );
in01f80 g740930 ( .a(n_39146), .o(n_39147) );
oa22f80 g739801 ( .a(n_40383), .b(n_40330), .c(n_40349), .d(n_40331), .o(n_40433) );
in01f80 g753294 ( .a(n_27028), .o(n_27044) );
ao22s80 g768517 ( .a(n_12286), .b(n_12334), .c(n_12285), .d(n_12291), .o(n_13366) );
na02f80 g775054 ( .a(n_6077), .b(n_5966), .o(n_6155) );
no02f80 g745024 ( .a(n_34768), .b(n_34396), .o(n_34794) );
in01f80 g756049 ( .a(n_25162), .o(n_25217) );
no02f80 g780912 ( .a(n_420), .b(n_439), .o(n_480) );
na02f80 g747736 ( .a(n_33571), .b(n_33684), .o(n_33699) );
no02f80 g777593 ( .a(n_3394), .b(n_3151), .o(n_3475) );
ms00f80 sin_out_reg_12_ ( .ck(newNet_84), .d(n_43802), .o(sin_out_12) );
no02f80 g784596 ( .a(FE_OCP_RBN2716_n_14982), .b(n_14190), .o(n_46419) );
na03f80 g780472 ( .a(n_951), .b(n_977), .c(n_976), .o(n_978) );
in01f80 newInst_3526 ( .a(newNet_3525), .o(newNet_3526) );
no02f80 g777294 ( .a(n_4675), .b(n_5165), .o(n_5188) );
in01f80 newInst_3550 ( .a(newNet_278), .o(newNet_3550) );
in01f80 g763725 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .o(n_16779) );
in01f80 newInst_59 ( .a(newNet_58), .o(newNet_59) );
ao22s80 g775069 ( .a(n_6017), .b(n_5907), .c(n_5996), .d(n_5910), .o(n_6108) );
no02f80 g765664 ( .a(n_15001), .b(n_13476), .o(n_15137) );
ao12f80 g757895 ( .a(n_22814), .b(n_22854), .c(n_22813), .o(n_23812) );
na02f80 g776646 ( .a(n_4436), .b(n_4435), .o(n_4492) );
no02f80 g754901 ( .a(n_25210), .b(n_24199), .o(n_25359) );
no02f80 g763079 ( .a(n_17903), .b(n_17902), .o(n_17904) );
no02f80 g757308 ( .a(n_23468), .b(n_23448), .o(n_23449) );
na02f80 g748009 ( .a(n_32982), .b(n_32556), .o(n_33040) );
in01f80 g768626 ( .a(n_12230), .o(n_12231) );
in01f80 g751592 ( .a(n_28647), .o(n_28599) );
na02f80 g758292 ( .a(n_22288), .b(n_20859), .o(n_22410) );
in01f80 newInst_778 ( .a(newNet_777), .o(newNet_778) );
in01f80 g753786 ( .a(n_26444), .o(n_26465) );
ao12f80 g763610 ( .a(n_17575), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .o(n_18382) );
in01f80 FE_OCP_RBC1838_n_19528 ( .a(n_19528), .o(FE_OCP_RBN1838_n_19528) );
na02f80 g741838 ( .a(n_38340), .b(n_38219), .o(n_38420) );
ao22s80 FE_RC_4133_0 ( .a(n_12888), .b(FE_OCP_RBN2206_n_12907), .c(n_12907), .d(FE_OCP_RBN2220_n_12888), .o(n_13096) );
na02f80 g754543 ( .a(n_26641), .b(n_26640), .o(n_26642) );
na02f80 g760386 ( .a(n_20129), .b(n_20148), .o(n_20228) );
na02f80 g758610 ( .a(n_21817), .b(n_20206), .o(n_21925) );
no02f80 g741624 ( .a(FE_OCP_RBN2398_n_38586), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38614) );
in01f80 newInst_3606 ( .a(newNet_2403), .o(newNet_3606) );
in01f80 g752721 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_), .o(n_28365) );
na02f80 g749242 ( .a(n_32094), .b(n_31457), .o(n_32116) );
in01f80 FE_OCPC1445_n_31473 ( .a(FE_OCP_DRV_N1608_n_31473), .o(FE_OCPN1445_n_31473) );
in01f80 newInst_2857 ( .a(newNet_2342), .o(newNet_2857) );
in01f80 newInst_2264 ( .a(newNet_2263), .o(newNet_2264) );
in01f80 g745331 ( .a(n_36164), .o(n_36165) );
ao12f80 g783822 ( .a(n_40619), .b(n_45507), .c(n_44610), .o(n_45508) );
na02f80 g739055 ( .a(n_41112), .b(n_41111), .o(n_41113) );
no02f80 g746242 ( .a(n_33642), .b(n_33594), .o(n_33621) );
in01f80 g772786 ( .a(n_8093), .o(n_8169) );
in01f80 g739174 ( .a(n_40942), .o(n_40960) );
in01f80 g747781 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38778) );
na02f80 FE_RC_2396_0 ( .a(n_42392), .b(FE_RN_941_0), .o(FE_RN_942_0) );
in01f80 g740894 ( .a(n_39310), .o(n_39217) );
oa22f80 g737177 ( .a(n_42974), .b(n_42693), .c(n_42973), .d(n_42694), .o(n_43001) );
no02f80 g775976 ( .a(n_4729), .b(n_4601), .o(n_4730) );
ao22s80 g767729 ( .a(n_13069), .b(n_12229), .c(n_13317), .d(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .o(n_13440) );
ao12f80 g771644 ( .a(n_8856), .b(n_8907), .c(n_8855), .o(n_9042) );
no02f80 g740540 ( .a(n_39709), .b(n_39713), .o(n_39748) );
na02f80 g737757 ( .a(n_42657), .b(n_42609), .o(n_42679) );
in01f80 FE_OCP_DRV_C1591_n_34327 ( .a(n_34327), .o(FE_OCP_DRV_N1591_n_34327) );
oa22f80 g748026 ( .a(n_31972), .b(n_32178), .c(n_31954), .d(n_32179), .o(n_32251) );
na02f80 FE_RC_1928_0 ( .a(FE_RN_610_0), .b(n_29273), .o(FE_RN_611_0) );
in01f80 g752675 ( .a(n_28138), .o(n_28158) );
in01f80 newInst_1256 ( .a(newNet_1255), .o(newNet_1256) );
in01f80 g772011 ( .a(n_9431), .o(n_9432) );
no02f80 g743109 ( .a(n_35713), .b(delay_sub_ln21_unr24_stage9_stallmux_q_7_), .o(n_37090) );
in01f80 g756311 ( .a(FE_OCPN3164_n_24117), .o(n_24116) );
in01f80 g755088 ( .a(n_25154), .o(n_25125) );
no02f80 g743043 ( .a(n_37147), .b(n_37146), .o(n_37386) );
no02f80 g754307 ( .a(n_25894), .b(n_25669), .o(n_26016) );
na02f80 g774814 ( .a(n_6311), .b(n_6172), .o(n_6344) );
oa22f80 g744624 ( .a(n_36574), .b(n_35992), .c(n_36596), .d(n_35993), .o(n_36661) );
na02f80 FE_RC_1559_0 ( .a(FE_RN_441_0), .b(FE_RN_442_0), .o(FE_RN_443_0) );
in01f80 g762688 ( .a(n_18052), .o(n_17893) );
na02f80 g739162 ( .a(n_40958), .b(n_40853), .o(n_40956) );
na02f80 g758299 ( .a(n_22288), .b(n_21324), .o(n_22405) );
na02f80 g767609 ( .a(n_13100), .b(n_12832), .o(n_13178) );
in01f80 newInst_3336 ( .a(newNet_3335), .o(newNet_3336) );
ao12f80 g751432 ( .a(FE_OCP_RBN2192_n_28597), .b(n_28647), .c(n_28646), .o(n_28648) );
na02f80 FE_RC_2582_0 ( .a(FE_RN_1065_0), .b(n_3365), .o(FE_RN_1066_0) );
na02f80 g740509 ( .a(n_39699), .b(n_38787), .o(n_39724) );
no02f80 g776447 ( .a(n_4643), .b(n_4642), .o(n_4799) );
oa22f80 g769017 ( .a(n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .c(FE_OCP_RBN3273_n_45224), .d(n_11593), .o(n_11761) );
na02f80 g754334 ( .a(FE_OCP_RBN1200_n_25763), .b(n_27416), .o(n_25827) );
in01f80 g741085 ( .a(n_39800), .o(n_39817) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_0_ ( .ck(newNet_472), .d(n_27652), .o(delay_xor_ln22_unr18_stage7_stallmux_q_0_) );
na02f80 g779244 ( .a(n_1853), .b(n_1842), .o(n_1843) );
no02f80 g763153 ( .a(n_17479), .b(n_17478), .o(n_17504) );
no02f80 g741212 ( .a(n_38818), .b(n_38817), .o(n_38831) );
na02f80 g749760 ( .a(n_29875), .b(n_29873), .o(n_29874) );
in01f80 g749097 ( .a(n_30960), .o(n_31029) );
in01f80 newInst_3359 ( .a(newNet_3358), .o(newNet_3359) );
in01f80 FE_OCP_RBC1380_n_21240 ( .a(n_21240), .o(FE_OCP_RBN1380_n_21240) );
no03m80 FE_RC_1535_0 ( .a(n_27999), .b(n_28096), .c(FE_RN_434_0), .o(n_28123) );
in01f80 g736437 ( .a(n_43731), .o(n_43732) );
in01f80 newInst_121 ( .a(newNet_120), .o(newNet_121) );
in01f80 g771924 ( .a(FE_OCP_RBN2499_n_8835), .o(n_10226) );
in01f80 g771339 ( .a(n_9114), .o(n_9197) );
in01f80 g770580 ( .a(n_10153), .o(n_10228) );
in01f80 FE_OCP_RBC3632_n_20568 ( .a(n_20568), .o(FE_OCP_RBN3632_n_20568) );
in01f80 newInst_654 ( .a(newNet_539), .o(newNet_654) );
no02f80 g765643 ( .a(n_15019), .b(FE_OCP_RBN2757_FE_RN_722_0), .o(n_15041) );
oa12f80 g767995 ( .a(n_12762), .b(n_12761), .c(n_12760), .o(n_12852) );
in01f80 g766900 ( .a(n_13657), .o(n_13658) );
na02f80 g763498 ( .a(n_16835), .b(n_16899), .o(n_16984) );
no02f80 g749062 ( .a(n_32230), .b(n_31542), .o(n_32295) );
ao12f80 g741862 ( .a(n_38296), .b(n_38243), .c(n_38309), .o(n_38438) );
no02f80 g765350 ( .a(n_15293), .b(n_15806), .o(n_15374) );
ao12f80 g752835 ( .a(n_28107), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n_28713) );
no02f80 g762998 ( .a(n_17562), .b(n_17517), .o(n_17679) );
in01f80 g779208 ( .a(n_1856), .o(n_1857) );
in01f80 g748149 ( .a(n_32136), .o(n_32137) );
na02f80 g750049 ( .a(n_29896), .b(n_30364), .o(n_30423) );
in01f80 FE_OCP_RBC2357_n_13818 ( .a(n_13818), .o(FE_OCP_RBN2357_n_13818) );
in01f80 FE_OCPC1247_n_43120 ( .a(FE_OCPN1245_n_43120), .o(FE_OCPN1247_n_43120) );
no02f80 g760138 ( .a(n_20404), .b(FE_OCP_RBN1696_n_19206), .o(n_20491) );
in01f80 FE_RC_671_0 ( .a(n_28290), .o(FE_RN_213_0) );
in01f80 newInst_3421 ( .a(newNet_1787), .o(newNet_3421) );
ao12f80 g752696 ( .a(n_27361), .b(n_27362), .c(n_27125), .o(n_27440) );
oa22f80 g752572 ( .a(n_27569), .b(n_27457), .c(n_27570), .d(n_27458), .o(n_27643) );
ao12f80 g737474 ( .a(n_42604), .b(n_42603), .c(n_42602), .o(n_43130) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_10_ ( .ck(newNet_2030), .d(n_10783), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_) );
na02f80 g770826 ( .a(n_10138), .b(n_10137), .o(n_10174) );
ao12f80 g751067 ( .a(n_30304), .b(n_30303), .c(n_29907), .o(n_30418) );
in01f80 g780123 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_24_), .o(n_1197) );
na02f80 g762270 ( .a(FE_OFN750_n_45003), .b(n_18660), .o(n_18816) );
na02f80 g760956 ( .a(n_19225), .b(n_18460), .o(n_19284) );
na02f80 g780211 ( .a(n_1041), .b(n_45809), .o(n_1116) );
na02f80 g745402 ( .a(n_35543), .b(n_35542), .o(n_35561) );
na02f80 g776314 ( .a(n_4552), .b(n_3951), .o(n_4626) );
no02f80 g780376 ( .a(n_858), .b(n_782), .o(n_995) );
na02f80 g770611 ( .a(n_10270), .b(FE_OCP_RBN3638_n_44490), .o(n_10398) );
ao12f80 g753408 ( .a(n_26769), .b(n_27589), .c(n_26832), .o(n_27611) );
oa22f80 FE_RC_887_0 ( .a(FE_OCP_RBN2365_n_24372), .b(n_24787), .c(n_24529), .d(n_24836), .o(n_24944) );
no02f80 g749445 ( .a(FE_OCP_RBN2755_n_30558), .b(n_30263), .o(n_30576) );
na02f80 g762614 ( .a(n_18022), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .o(n_18088) );
in01f80 FE_OCP_RBC3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
no02f80 g768281 ( .a(n_12553), .b(n_12551), .o(n_12552) );
na02f80 g764107 ( .a(n_16518), .b(n_16495), .o(n_16567) );
no02f80 g748239 ( .a(FE_OCP_RBN3083_n_31819), .b(n_31871), .o(n_31872) );
no02f80 g745396 ( .a(FE_OCP_RBN2987_n_35539), .b(n_36019), .o(n_36050) );
na02f80 g742588 ( .a(n_37469), .b(n_37468), .o(n_37470) );
na02f80 g753689 ( .a(n_26616), .b(n_26558), .o(n_26702) );
na02f80 g760684 ( .a(n_19635), .b(n_19101), .o(n_19672) );
no02f80 g752058 ( .a(n_28121), .b(n_28120), .o(n_28122) );
no02f80 FE_RC_2309_0 ( .a(FE_RN_875_0), .b(n_25904), .o(n_25948) );
in01f80 g758110 ( .a(n_22131), .o(n_22130) );
in01f80 FE_OCP_RBC2689_n_38870 ( .a(FE_OCP_RBN2688_n_38870), .o(FE_OCP_RBN2689_n_38870) );
na02f80 g778094 ( .a(n_2866), .b(n_2865), .o(n_2867) );
no02f80 g759551 ( .a(n_20767), .b(n_20332), .o(n_20768) );
na02f80 g763285 ( .a(n_17227), .b(n_17226), .o(n_17228) );
no02f80 g769699 ( .a(n_11226), .b(n_11179), .o(n_11294) );
in01f80 g766878 ( .a(n_14491), .o(n_14422) );
no02f80 g760312 ( .a(n_20081), .b(n_20022), .o(n_20193) );
no02f80 g760128 ( .a(n_20537), .b(FE_OCPN1782_FE_OCP_RBN1701_n_19353), .o(n_20531) );
in01f80 newInst_3640 ( .a(newNet_3639), .o(newNet_3640) );
no02f80 g767681 ( .a(n_13083), .b(n_13173), .o(n_13180) );
na02f80 g749248 ( .a(n_30653), .b(n_30559), .o(n_30713) );
na02f80 g755241 ( .a(n_25686), .b(n_25685), .o(n_25687) );
ao22s80 FE_RC_551_0 ( .a(FE_OCPN1410_n_27014), .b(n_30507), .c(n_30466), .d(n_30492), .o(n_30575) );
na02f80 g755831 ( .a(n_24998), .b(n_25005), .o(n_25058) );
no02f80 g737697 ( .a(n_42216), .b(n_41915), .o(n_42474) );
in01f80 g781195 ( .a(n_174), .o(n_171) );
na02f80 g776767 ( .a(n_3831), .b(n_2947), .o(n_3993) );
na02f80 g749936 ( .a(n_29864), .b(n_29890), .o(n_29927) );
na02f80 g757765 ( .a(n_22592), .b(n_22442), .o(n_22623) );
no02f80 g755529 ( .a(n_24510), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24539) );
no02f80 g742926 ( .a(n_37159), .b(n_37048), .o(n_37207) );
na02f80 g741477 ( .a(n_38790), .b(n_38773), .o(n_38808) );
in01f80 newInst_1620 ( .a(newNet_1619), .o(newNet_1620) );
na02f80 g749543 ( .a(n_30436), .b(n_30114), .o(n_30498) );
in01f80 g760551 ( .a(n_19944), .o(n_19963) );
no02f80 g768547 ( .a(FE_OCP_RBN2163_n_12312), .b(n_11945), .o(n_12345) );
in01f80 g779036 ( .a(n_2154), .o(n_2155) );
na02f80 g746788 ( .a(n_33078), .b(n_33077), .o(n_33082) );
in01f80 g776044 ( .a(n_5226), .o(n_5227) );
in01f80 FE_RC_4166_0 ( .a(n_18333), .o(FE_RN_1815_0) );
in01f80 newInst_993 ( .a(newNet_992), .o(newNet_993) );
no02f80 FE_RC_497_0 ( .a(FE_RN_147_0), .b(FE_RN_148_0), .o(FE_RN_149_0) );
no02f80 g755983 ( .a(n_24264), .b(n_23789), .o(n_24290) );
ao12f80 g766044 ( .a(n_14994), .b(n_14993), .c(n_14992), .o(n_15823) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_26_ ( .ck(newNet_2086), .d(FE_OCP_RBN3123_n_6557), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_) );
in01f80 g754647 ( .a(n_27131), .o(n_27315) );
na02f80 g779727 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(n_1794) );
no02f80 g761352 ( .a(n_19028), .b(n_19027), .o(n_19029) );
oa12f80 g755913 ( .a(n_25197), .b(n_25160), .c(n_25132), .o(n_25802) );
na02f80 g767092 ( .a(n_13432), .b(n_12848), .o(n_13513) );
in01f80 g761807 ( .a(n_18642), .o(n_20635) );
na02f80 g739772 ( .a(n_40468), .b(n_40295), .o(n_40509) );
no02f80 g758903 ( .a(FE_OCP_RBN3220_n_21358), .b(n_21226), .o(n_21431) );
oa12f80 g751926 ( .a(n_28858), .b(n_28897), .c(n_28834), .o(n_29409) );
oa12f80 g778637 ( .a(n_2590), .b(n_3297), .c(n_2577), .o(n_3409) );
oa22f80 g769312 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .c(n_11542), .d(FE_OCPN1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12094) );
in01f80 FE_OFC737_n_22641 ( .a(FE_OFN734_n_22641), .o(FE_OFN737_n_22641) );
in01f80 g767836 ( .a(n_12795), .o(n_14685) );
no02f80 g758096 ( .a(n_21973), .b(FE_OCP_RBN1844_n_20910), .o(n_22048) );
na02f80 g775456 ( .a(n_5723), .b(n_4376), .o(n_5886) );
na02f80 g764588 ( .a(n_16154), .b(n_16109), .o(n_16110) );
no02f80 g771595 ( .a(n_10341), .b(n_10340), .o(n_10385) );
ao22s80 FE_RC_3709_0 ( .a(n_43612), .b(n_43882), .c(n_43611), .d(n_43883), .o(n_43908) );
oa22f80 g784343 ( .a(FE_OFN774_n_46137), .b(n_6318), .c(n_46195), .d(n_46994), .o(n_46149) );
na02f80 g761542 ( .a(n_19545), .b(n_19544), .o(n_19546) );
in01f80 g753109 ( .a(n_27546), .o(n_27547) );
in01f80 FE_OCP_RBC2938_n_26456 ( .a(n_26456), .o(FE_OCP_RBN2938_n_26456) );
in01f80 g767443 ( .a(n_13139), .o(n_13175) );
na02f80 g771895 ( .a(n_8698), .b(n_8678), .o(n_8784) );
in01f80 g760665 ( .a(n_19748), .o(n_19749) );
na02f80 g751188 ( .a(n_29782), .b(n_28929), .o(n_29853) );
na02f80 g743937 ( .a(n_36901), .b(n_46209), .o(n_36942) );
no02f80 FE_RC_2574_0 ( .a(n_2935), .b(n_2900), .o(FE_RN_1058_0) );
na02f80 g762327 ( .a(n_18126), .b(n_18146), .o(n_18198) );
na03f80 FE_RC_1657_0 ( .a(n_36917), .b(n_36932), .c(n_36931), .o(n_37033) );
ao12f80 g745770 ( .a(n_34145), .b(n_44102), .c(n_34127), .o(n_34657) );
in01f80 g743676 ( .a(n_36394), .o(n_36395) );
no02f80 g757602 ( .a(n_22795), .b(n_44061), .o(n_22796) );
no02f80 g737685 ( .a(n_42367), .b(n_42366), .o(n_42443) );
in01f80 g741129 ( .a(n_39360), .o(n_39361) );
in01f80 newInst_40 ( .a(newNet_10), .o(newNet_40) );
no02f80 g760470 ( .a(n_20062), .b(n_19583), .o(n_20063) );
in01f80 g755311 ( .a(n_25036), .o(n_25037) );
no02f80 g737463 ( .a(n_42599), .b(n_42630), .o(n_42653) );
na02f80 g747257 ( .a(n_32811), .b(n_32810), .o(n_32812) );
in01f80 FE_OCP_RBC2744_n_15319 ( .a(n_15319), .o(FE_OCP_RBN2744_n_15319) );
na02f80 g756931 ( .a(n_23806), .b(n_23803), .o(n_23950) );
no02f80 g778137 ( .a(n_2899), .b(n_2898), .o(n_2922) );
in01f80 FE_OCPC1477_n_28775 ( .a(n_28775), .o(FE_OCPN1477_n_28775) );
no02f80 g778367 ( .a(n_2686), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_), .o(n_2798) );
in01f80 g770159 ( .a(n_10892), .o(n_10893) );
in01f80 g745682 ( .a(n_34286), .o(n_34369) );
in01f80 newInst_783 ( .a(newNet_782), .o(newNet_783) );
na02f80 g759940 ( .a(n_21374), .b(n_21370), .o(n_21624) );
na02f80 g753244 ( .a(n_27113), .b(n_27243), .o(n_27214) );
no02f80 g771997 ( .a(FE_OCP_RBN3574_n_44563), .b(n_9151), .o(n_9322) );
ao22s80 g763716 ( .a(n_17259), .b(n_17427), .c(n_17258), .d(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_18418) );
na02f80 g760307 ( .a(n_20228), .b(n_18944), .o(n_20285) );
na02f80 g758577 ( .a(n_21905), .b(n_21815), .o(n_21906) );
in01f80 g743641 ( .a(n_36514), .o(n_36481) );
no02f80 g764455 ( .a(n_16124), .b(n_45331), .o(n_16193) );
in01f80 g744634 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_36578) );
oa22f80 g784530 ( .a(n_12144), .b(FE_OFN802_n_46285), .c(n_12112), .d(FE_OFN771_n_46337), .o(n_46351) );
no02f80 g771399 ( .a(n_9641), .b(n_9640), .o(n_9721) );
na02f80 g741869 ( .a(n_38286), .b(n_38083), .o(n_38340) );
in01f80 newInst_2753 ( .a(newNet_2752), .o(newNet_2753) );
in01f80 newInst_1495 ( .a(newNet_1494), .o(newNet_1495) );
ao12f80 g773020 ( .a(n_7762), .b(n_7761), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n_9324) );
ao22s80 g778646 ( .a(n_2455), .b(n_2047), .c(n_2434), .d(n_2046), .o(n_2550) );
no02f80 g742120 ( .a(n_38078), .b(n_38157), .o(n_38486) );
na02f80 g736675 ( .a(n_43282), .b(n_43231), .o(n_43332) );
oa12f80 g772035 ( .a(n_8652), .b(n_8692), .c(n_8651), .o(n_8766) );
in01f80 FE_RC_2590_0 ( .a(FE_RN_1072_0), .o(n_12230) );
ao12f80 g746185 ( .a(n_33690), .b(n_33711), .c(n_33689), .o(n_33775) );
in01f80 FE_OCP_RBC1694_n_19052 ( .a(FE_OCP_RBN1693_n_19052), .o(FE_OCP_RBN1694_n_19052) );
na02f80 g774278 ( .a(n_6717), .b(n_6737), .o(n_6718) );
ao12f80 g745984 ( .a(n_34635), .b(n_35218), .c(n_34697), .o(n_35321) );
in01f80 g753183 ( .a(n_27150), .o(n_27233) );
in01f80 g743449 ( .a(n_36751), .o(n_36701) );
in01f80 FE_OCP_RBC3396_n_28651 ( .a(n_28651), .o(FE_OCP_RBN3396_n_28651) );
in01f80 g761200 ( .a(n_19060), .o(n_19061) );
in01f80 FE_OCPC962_n_28506 ( .a(FE_OCPN961_n_28506), .o(FE_OCPN962_n_28506) );
in01f80 FE_OCP_RBC2693_n_15083 ( .a(n_15083), .o(FE_OCP_RBN2693_n_15083) );
in01f80 g756493 ( .a(n_23788), .o(n_23789) );
na02f80 g752130 ( .a(n_28012), .b(n_27872), .o(n_28071) );
no02f80 g737498 ( .a(n_42541), .b(n_42589), .o(n_42635) );
in01f80 newInst_2157 ( .a(newNet_2156), .o(newNet_2157) );
na02f80 g751881 ( .a(n_28956), .b(n_29006), .o(n_29007) );
na02f80 g739380 ( .a(n_40810), .b(n_40809), .o(n_41127) );
in01f80 fopt783810 ( .a(FE_OCP_RBN2341_n_29470), .o(n_45489) );
na02f80 g765621 ( .a(n_15103), .b(n_14238), .o(n_15172) );
na02f80 g766275 ( .a(n_14436), .b(n_14398), .o(n_14461) );
na02f80 g737674 ( .a(n_42392), .b(n_41982), .o(n_42700) );
in01f80 FE_OCP_RBC3125_n_27578 ( .a(n_27578), .o(FE_OCP_RBN3125_n_27578) );
in01f80 FE_OCPC1233_n_2414 ( .a(n_2414), .o(FE_OCPN1233_n_2414) );
oa12f80 g773448 ( .a(n_7207), .b(n_7534), .c(n_7167), .o(n_7542) );
oa12f80 g748788 ( .a(n_31263), .b(n_31262), .c(n_31261), .o(n_31326) );
ao22s80 g769627 ( .a(n_11340), .b(n_11332), .c(n_11317), .d(n_11331), .o(n_11409) );
na02f80 g757087 ( .a(n_23232), .b(n_23249), .o(n_23332) );
oa12f80 g762300 ( .a(n_18058), .b(n_18080), .c(n_18057), .o(n_18111) );
oa12f80 g760051 ( .a(n_20914), .b(n_20275), .c(n_20293), .o(n_20378) );
no02f80 g766064 ( .a(FE_OCP_RBN3591_n_14704), .b(n_14758), .o(n_14759) );
ao12f80 g761221 ( .a(n_19787), .b(n_19712), .c(n_19986), .o(n_20037) );
in01f80 FE_OCP_RBC2685_n_38870 ( .a(n_38870), .o(FE_OCP_RBN2685_n_38870) );
no02f80 g761330 ( .a(n_19952), .b(n_19845), .o(n_20012) );
ao12f80 g774836 ( .a(n_5260), .b(n_6266), .c(n_5329), .o(n_6316) );
in01f80 FE_OCP_RBC1206_n_16814 ( .a(n_16814), .o(FE_OCP_RBN1206_n_16814) );
in01f80 g775594 ( .a(n_47270), .o(n_5765) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_15_ ( .ck(newNet_360), .d(n_1292), .o(delay_xor_ln22_unr3_stage2_stallmux_q_15_) );
in01f80 g758273 ( .a(n_22411), .o(n_22436) );
in01f80 g768262 ( .a(n_12695), .o(n_12696) );
na02f80 g740959 ( .a(n_39252), .b(n_39273), .o(n_39333) );
in01f80 fopt782839 ( .a(n_27620), .o(n_44265) );
in01f80 g741164 ( .a(n_38886), .o(n_38887) );
in01f80 newInst_1892 ( .a(newNet_1891), .o(newNet_1892) );
in01f80 FE_OCP_RBC2417_n_24720 ( .a(n_24720), .o(FE_OCP_RBN2417_n_24720) );
no02f80 g761310 ( .a(n_18872), .b(n_18514), .o(n_18925) );
in01f80 g779783 ( .a(n_1422), .o(n_1463) );
in01f80 g739941 ( .a(n_40369), .o(n_40370) );
ms00f80 sin_out_reg_17_ ( .ck(newNet_68), .d(n_43890), .o(sin_out_17) );
na02f80 g742767 ( .a(n_37389), .b(n_37253), .o(n_37439) );
no04s80 FE_RC_733_0 ( .a(FE_OCPN908_n_23227), .b(n_23226), .c(n_23126), .d(n_23038), .o(n_23228) );
in01f80 FE_OCP_RBC2115_n_45224 ( .a(FE_OCP_RBN3266_n_45224), .o(FE_OCP_RBN2115_n_45224) );
in01f80 newInst_26 ( .a(newNet_2), .o(newNet_26) );
in01f80 g776514 ( .a(n_4103), .o(n_4104) );
na02f80 g740564 ( .a(n_39705), .b(n_38795), .o(n_39730) );
no02f80 g740404 ( .a(n_39942), .b(n_39602), .o(n_40308) );
in01f80 g747570 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .o(n_32464) );
in01f80 fopt783532 ( .a(n_45145), .o(n_45144) );
na02f80 g752903 ( .a(n_27050), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27882) );
oa22f80 g772213 ( .a(n_8523), .b(n_7640), .c(n_8524), .d(n_7639), .o(n_8637) );
na02f80 g762436 ( .a(n_18043), .b(n_17918), .o(n_18073) );
na02f80 g746121 ( .a(n_33677), .b(n_33178), .o(n_33737) );
in01f80 g775899 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_6_), .o(n_5312) );
in01f80 newInst_549 ( .a(newNet_234), .o(newNet_549) );
oa12f80 g756878 ( .a(n_24061), .b(n_24188), .c(n_24023), .o(n_24675) );
in01f80 g770644 ( .a(FE_OCP_RBN2798_n_10106), .o(n_10278) );
no02f80 FE_RC_3060_0 ( .a(FE_RN_1342_0), .b(n_26920), .o(n_46422) );
na02f80 g739891 ( .a(n_40297), .b(n_39996), .o(n_40402) );
in01f80 FE_OCPC1423_delay_sub_ln23_0_unr21_stage8_stallmux_q ( .a(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(FE_OCPN1423_delay_sub_ln23_0_unr21_stage8_stallmux_q) );
na02f80 g753825 ( .a(n_26405), .b(n_23486), .o(n_26467) );
in01f80 g747456 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .o(n_32388) );
na02f80 g764560 ( .a(n_16001), .b(n_16048), .o(n_16049) );
in01f80 g751124 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30546) );
no02f80 g776883 ( .a(n_3965), .b(n_3901), .o(n_4212) );
no02f80 g761486 ( .a(n_19649), .b(n_18935), .o(n_19993) );
in01f80 g750620 ( .a(n_29401), .o(n_29418) );
no02f80 g765779 ( .a(n_15288), .b(n_14490), .o(n_15481) );
in01f80 newInst_2126 ( .a(newNet_2125), .o(newNet_2126) );
ao12f80 g772765 ( .a(n_8098), .b(n_8097), .c(n_8096), .o(n_9223) );
no02f80 g745078 ( .a(n_34688), .b(n_34239), .o(n_34729) );
in01f80 FE_OCPC1860_n_35415 ( .a(FE_OCPN1859_n_35415), .o(FE_OCPN1860_n_35415) );
oa12f80 g765248 ( .a(n_15227), .b(n_15226), .c(n_15225), .o(n_15303) );
oa12f80 g742360 ( .a(n_37777), .b(n_37817), .c(n_37757), .o(n_37853) );
in01f80 newInst_2580 ( .a(newNet_2579), .o(newNet_2580) );
oa22f80 g755940 ( .a(n_25160), .b(n_24236), .c(n_25188), .d(n_25092), .o(n_25437) );
na02f80 g759970 ( .a(n_20581), .b(n_20456), .o(n_20634) );
no02f80 g744078 ( .a(n_44223), .b(n_35005), .o(n_36144) );
in01f80 FE_OCP_DRV_C1567_n_19751 ( .a(n_19751), .o(FE_OCP_DRV_N1567_n_19751) );
oa12f80 g760473 ( .a(n_20517), .b(n_20516), .c(n_20515), .o(n_21373) );
in01f80 newInst_3305 ( .a(newNet_1285), .o(newNet_3305) );
in01f80 g749959 ( .a(n_29834), .o(n_29835) );
ao22s80 g736481 ( .a(n_43711), .b(n_43552), .c(FE_OCP_RBN3109_n_43711), .d(n_43551), .o(n_43760) );
in01f80 g771017 ( .a(n_10027), .o(n_10083) );
in01f80 FE_OCP_RBC3474_n_7886 ( .a(FE_OCP_RBN3470_n_7886), .o(FE_OCP_RBN3474_n_7886) );
ao12f80 g764923 ( .a(n_15391), .b(n_15320), .c(FE_OCP_RBN2715_n_14982), .o(n_15438) );
na02f80 g761264 ( .a(n_19902), .b(n_19903), .o(n_19958) );
in01f80 g754460 ( .a(n_26869), .o(n_26870) );
oa12f80 g747586 ( .a(n_32068), .b(n_45755), .c(n_47272), .o(n_32349) );
in01f80 g753142 ( .a(n_27490), .o(n_27491) );
na02f80 g752116 ( .a(n_28097), .b(n_28119), .o(n_28221) );
no02f80 g764692 ( .a(n_15812), .b(n_15524), .o(n_15813) );
no02f80 g745387 ( .a(n_36049), .b(n_35926), .o(n_36080) );
na02f80 g765550 ( .a(n_15103), .b(n_14152), .o(n_15181) );
in01f80 g764486 ( .a(n_16158), .o(n_16159) );
ao12f80 g755494 ( .a(n_24982), .b(n_25468), .c(n_25407), .o(n_25526) );
na02f80 g776051 ( .a(n_5110), .b(n_5109), .o(n_5216) );
in01f80 newInst_3520 ( .a(newNet_1925), .o(newNet_3520) );
in01f80 g775205 ( .a(n_5963), .o(n_5986) );
ao12f80 g757274 ( .a(n_23077), .b(n_44068), .c(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .o(n_23107) );
na02f80 g750976 ( .a(n_28934), .b(FE_OCP_RBN3395_n_28651), .o(n_28948) );
in01f80 g774216 ( .a(n_6689), .o(n_6690) );
in01f80 g742989 ( .a(n_36968), .o(n_37131) );
in01f80 g763608 ( .a(n_16808), .o(n_16880) );
no02f80 g757390 ( .a(n_44084), .b(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .o(n_23307) );
in01f80 newInst_1470 ( .a(newNet_1469), .o(newNet_1470) );
na02f80 g779536 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n_1382) );
no02f80 g770713 ( .a(n_10236), .b(n_10152), .o(n_10379) );
no02f80 g769772 ( .a(n_46424), .b(FE_OCP_RBN3036_n_47269), .o(n_11167) );
na02f80 g751413 ( .a(n_28527), .b(n_28520), .o(n_28610) );
in01f80 g773762 ( .a(n_7234), .o(n_7235) );
no02f80 g741528 ( .a(n_38732), .b(n_38731), .o(n_38754) );
in01f80 FE_RC_1425_0 ( .a(FE_RN_416_0), .o(n_22556) );
na02f80 g774767 ( .a(n_6412), .b(n_6326), .o(n_6471) );
na02f80 g763247 ( .a(n_16917), .b(n_16833), .o(n_16954) );
no02f80 FE_RC_2465_0 ( .a(FE_RN_988_0), .b(FE_RN_990_0), .o(n_14435) );
in01f80 FE_OCP_RBC3505_n_13860 ( .a(FE_OCP_RBN2388_n_13860), .o(FE_OCP_RBN3505_n_13860) );
na02f80 g745756 ( .a(n_34338), .b(FE_OCP_RBN2451_n_34278), .o(n_34362) );
no02f80 g753114 ( .a(n_27152), .b(n_27183), .o(n_27224) );
na02f80 g776976 ( .a(n_4034), .b(n_3957), .o(n_4209) );
na02f80 g739587 ( .a(FE_OCP_RBN3338_n_44610), .b(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n_40609) );
no02f80 g743163 ( .a(n_36946), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_), .o(n_37029) );
na02f80 g741329 ( .a(FE_OCP_RBN3582_n_44944), .b(n_38641), .o(n_39118) );
in01f80 g745408 ( .a(n_35634), .o(n_35724) );
no02f80 g759451 ( .a(n_20732), .b(n_20774), .o(n_20829) );
in01f80 newInst_3196 ( .a(newNet_213), .o(newNet_3196) );
in01f80 newInst_2776 ( .a(newNet_1200), .o(newNet_2776) );
na02f80 g772722 ( .a(n_8266), .b(n_7743), .o(n_8268) );
na02f80 g740786 ( .a(n_39463), .b(n_39322), .o(n_39512) );
ao22s80 FE_RC_773_0 ( .a(n_10322), .b(n_10511), .c(n_10323), .d(n_10512), .o(n_10644) );
in01f80 newInst_2618 ( .a(newNet_2242), .o(newNet_2618) );
no02f80 g757265 ( .a(n_23451), .b(n_23026), .o(n_23530) );
no02f80 g777325 ( .a(n_3690), .b(n_5242), .o(n_3797) );
in01f80 g755252 ( .a(n_24945), .o(n_24946) );
na02f80 g776738 ( .a(n_4156), .b(n_4263), .o(n_4264) );
na02f80 g761860 ( .a(n_18472), .b(n_18470), .o(n_18473) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_0_ ( .ck(newNet_1883), .d(FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(cordic_combinational_sub_ln23_0_unr16_z_0_) );
na02f80 g743522 ( .a(n_36489), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36510) );
na02f80 g758921 ( .a(n_21332), .b(n_21192), .o(n_21363) );
na02f80 g738388 ( .a(n_41416), .b(n_41391), .o(n_41455) );
in01f80 g763606 ( .a(n_16833), .o(n_16834) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_27_ ( .ck(newNet_800), .d(n_1299), .o(delay_xor_ln21_unr3_stage2_stallmux_q_27_) );
in01f80 newInst_2336 ( .a(newNet_2335), .o(newNet_2336) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_30_ ( .ck(newNet_3494), .d(n_22901), .o(delay_add_ln22_unr14_stage6_stallmux_q_30_) );
in01f80 g761056 ( .a(FE_OCPN969_n_19342), .o(n_19372) );
na02f80 g740853 ( .a(n_39378), .b(n_39398), .o(n_39881) );
no02f80 g745511 ( .a(n_34354), .b(n_34353), .o(n_34355) );
na02f80 g776174 ( .a(n_4555), .b(FE_OCP_RBN2723_n_4219), .o(n_4717) );
na02f80 g739145 ( .a(n_40943), .b(n_40794), .o(n_40962) );
na02f80 g760240 ( .a(FE_OCP_RBN3613_n_20249), .b(FE_OCP_RBN3834_n_19241), .o(n_20432) );
in01f80 g739604 ( .a(n_40654), .o(n_40649) );
na02f80 g737513 ( .a(n_42455), .b(n_42496), .o(n_42535) );
na02f80 g758007 ( .a(n_22263), .b(n_22083), .o(n_22303) );
in01f80 newInst_888 ( .a(newNet_887), .o(newNet_888) );
ao12f80 g770196 ( .a(n_10726), .b(n_10745), .c(n_10725), .o(n_10799) );
na02f80 g753708 ( .a(n_26580), .b(n_26478), .o(n_26581) );
no02f80 g745739 ( .a(n_34266), .b(n_34283), .o(n_34284) );
in01f80 g777746 ( .a(n_3303), .o(n_3279) );
na02f80 g745615 ( .a(n_34286), .b(n_33594), .o(n_34486) );
oa22f80 g757917 ( .a(n_22106), .b(n_22032), .c(n_22132), .d(n_22033), .o(n_22275) );
in01f80 FE_OCP_RBC3716_n_39913 ( .a(FE_OCP_RBN3715_n_39913), .o(FE_OCP_RBN3716_n_39913) );
na02f80 g772873 ( .a(n_7981), .b(n_7971), .o(n_8115) );
na02f80 g738142 ( .a(n_42079), .b(n_42078), .o(n_42080) );
oa12f80 g780712 ( .a(n_482), .b(n_626), .c(n_451), .o(n_631) );
in01f80 g776853 ( .a(n_4202), .o(n_4203) );
na02f80 g779016 ( .a(n_2075), .b(n_1506), .o(n_2132) );
in01f80 g758858 ( .a(n_21783), .o(n_21784) );
no02f80 g749260 ( .a(n_30814), .b(FE_OCPN1490_n_30823), .o(n_30846) );
na02f80 g764576 ( .a(n_16191), .b(n_14524), .o(n_16079) );
na02f80 g766016 ( .a(n_15030), .b(n_15029), .o(n_15031) );
oa22f80 g750025 ( .a(FE_OCPN1786_n_30134), .b(n_29553), .c(FE_OCP_RBN2571_n_29922), .d(FE_OCP_RBN3492_n_29553), .o(n_30401) );
ao12f80 g765220 ( .a(n_15840), .b(n_16245), .c(n_15748), .o(n_16256) );
na02f80 g773608 ( .a(n_7403), .b(n_7369), .o(n_7414) );
na02f80 g780574 ( .a(n_923), .b(n_610), .o(n_1015) );
no02f80 g748715 ( .a(n_31165), .b(n_31164), .o(n_31268) );
in01f80 g743209 ( .a(n_37661), .o(n_37739) );
oa12f80 g750453 ( .a(n_30521), .b(n_30552), .c(n_30520), .o(n_31253) );
in01f80 fopt783917 ( .a(n_36447), .o(n_45617) );
no02f80 g774061 ( .a(n_6797), .b(n_6740), .o(n_6973) );
in01f80 g743099 ( .a(n_37100), .o(n_37049) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_10_ ( .ck(newNet_370), .d(n_1325), .o(delay_xor_ln22_unr3_stage2_stallmux_q_10_) );
in01f80 g768950 ( .a(n_11873), .o(n_11841) );
na02f80 g779077 ( .a(n_2076), .b(n_1765), .o(n_2105) );
no02f80 g766125 ( .a(n_14519), .b(n_13272), .o(n_14558) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_29_ ( .ck(newNet_1586), .d(n_27656), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_) );
no02f80 g776348 ( .a(n_4517), .b(n_4422), .o(n_4592) );
no02f80 g739573 ( .a(n_40655), .b(n_40649), .o(n_40650) );
oa12f80 g773798 ( .a(n_6754), .b(n_7180), .c(n_6706), .o(n_7181) );
no02f80 g771196 ( .a(n_9552), .b(n_9352), .o(n_9458) );
na02f80 g775573 ( .a(n_5729), .b(n_5783), .o(n_5849) );
in01f80 g761678 ( .a(n_18861), .o(n_19027) );
in01f80 g770546 ( .a(n_10467), .o(n_10468) );
na02f80 g753492 ( .a(n_26874), .b(n_26873), .o(n_26982) );
na02f80 g744456 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_36775) );
no02f80 FE_RC_2739_0 ( .a(FE_RN_1160_0), .b(n_9450), .o(FE_RN_1161_0) );
ao12f80 g746281 ( .a(n_33206), .b(n_33476), .c(n_33105), .o(n_33549) );
ao12f80 g757770 ( .a(FE_OCP_RBN1710_n_22150), .b(n_22511), .c(n_22507), .o(n_22558) );
in01f80 g757259 ( .a(n_23197), .o(n_23134) );
no02f80 g777994 ( .a(n_3128), .b(n_3127), .o(n_3154) );
no02f80 g751706 ( .a(n_28366), .b(n_28365), .o(n_28387) );
ms00f80 cos_out_reg_20_ ( .ck(newNet_3724), .d(n_43860), .o(cos_out_20) );
in01f80 newInst_3091 ( .a(newNet_1401), .o(newNet_3091) );
in01f80 g750153 ( .a(n_30921), .o(n_30922) );
in01f80 FE_OCP_RBC3585_n_25295 ( .a(n_25295), .o(FE_OCP_RBN3585_n_25295) );
oa12f80 g771634 ( .a(n_8858), .b(n_8891), .c(n_8813), .o(n_9017) );
no02f80 g769188 ( .a(n_11838), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n_11866) );
no02f80 g753219 ( .a(n_27120), .b(n_25997), .o(n_27309) );
in01f80 g743808 ( .a(n_36046), .o(n_36324) );
ao22s80 FE_RC_612_0 ( .a(n_40969), .b(n_41213), .c(n_41214), .d(n_40970), .o(n_41285) );
in01f80 g746106 ( .a(n_33964), .o(n_34590) );
no02f80 g755869 ( .a(n_25284), .b(n_25340), .o(n_25341) );
in01f80 g769989 ( .a(n_10919), .o(n_10974) );
no02f80 g766118 ( .a(n_14571), .b(FE_OCP_RBN3534_n_13765), .o(n_14604) );
in01f80 g758837 ( .a(n_21511), .o(n_21512) );
no02f80 g757213 ( .a(n_23533), .b(n_23532), .o(n_23534) );
in01f80 FE_OCPC1460_n_37232 ( .a(FE_OCPN1459_n_37232), .o(FE_OCPN1460_n_37232) );
no02f80 g784787 ( .a(FE_OCP_RBN3085_n_31819), .b(n_31943), .o(n_47273) );
oa12f80 g767731 ( .a(n_12822), .b(n_12863), .c(n_12821), .o(n_13795) );
na02f80 g770358 ( .a(n_10689), .b(n_10657), .o(n_10658) );
no02f80 g745127 ( .a(n_34683), .b(n_34682), .o(n_34684) );
no02f80 g775808 ( .a(n_5354), .b(n_5317), .o(n_5461) );
no02f80 g771778 ( .a(n_9021), .b(FE_OCP_RBN3548_n_44575), .o(n_9105) );
in01f80 fopt783477 ( .a(n_45073), .o(n_45080) );
no02f80 g736942 ( .a(FE_OCPN912_n_43022), .b(n_43135), .o(n_43256) );
na02f80 g769559 ( .a(n_11350), .b(n_11303), .o(n_11393) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_15_ ( .ck(newNet_2212), .d(n_938), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_) );
in01f80 FE_OCP_RBC2813_n_25817 ( .a(n_25817), .o(FE_OCP_RBN2813_n_25817) );
no03m80 g751308 ( .a(n_44045), .b(n_29708), .c(n_28922), .o(n_29742) );
na02f80 g758252 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .o(n_22650) );
oa12f80 g770492 ( .a(n_10022), .b(n_10101), .c(n_10020), .o(n_10243) );
na02f80 g751744 ( .a(n_29029), .b(n_28988), .o(n_29079) );
in01f80 g738050 ( .a(n_42147), .o(n_42154) );
in01f80 FE_OCP_RBC1165_n_13726 ( .a(FE_OCP_RBN1164_n_13726), .o(FE_OCP_RBN1165_n_13726) );
in01f80 g755972 ( .a(FE_OFN788_n_25834), .o(n_29561) );
in01f80 g759215 ( .a(n_21014), .o(n_21015) );
oa22f80 g752662 ( .a(n_27441), .b(n_27191), .c(n_27440), .d(n_27190), .o(n_27534) );
in01f80 g754200 ( .a(n_26146), .o(n_26165) );
oa12f80 g739125 ( .a(n_40787), .b(n_40964), .c(n_40919), .o(n_41002) );
in01f80 g781353 ( .a(beta_30), .o(n_110) );
in01f80 g771975 ( .a(n_10037), .o(n_10038) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_10_ ( .ck(newNet_1771), .d(n_22115), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_) );
na02f80 g736572 ( .a(n_43682), .b(n_43473), .o(n_43683) );
no02f80 FE_RC_2218_0 ( .a(FE_RN_801_0), .b(n_32443), .o(FE_RN_802_0) );
na02f80 g763064 ( .a(n_17549), .b(n_17619), .o(n_17637) );
ao12f80 g762932 ( .a(n_17765), .b(FE_OCP_RBN2141_FE_OCPN861_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .o(n_17792) );
na02f80 g751713 ( .a(n_28385), .b(n_28033), .o(n_28386) );
na02f80 g771401 ( .a(n_9524), .b(n_9439), .o(n_9610) );
in01f80 FE_OCP_RBC3639_n_44490 ( .a(n_44490), .o(FE_OCP_RBN3639_n_44490) );
ao22s80 g757758 ( .a(FE_OCP_RBN3107_n_22590), .b(FE_OCP_RBN3101_n_22504), .c(n_22590), .d(n_22504), .o(n_22739) );
no02f80 g761087 ( .a(n_20016), .b(n_19960), .o(n_20039) );
na02f80 g741717 ( .a(n_38481), .b(n_38480), .o(n_38482) );
na02f80 g768878 ( .a(n_11907), .b(n_11692), .o(n_11908) );
no02f80 FE_RC_1814_0 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_6_), .b(n_17667), .o(FE_RN_539_0) );
no02f80 g774300 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .o(n_6964) );
na02f80 g772260 ( .a(n_8729), .b(n_8730), .o(n_8812) );
na02f80 FE_RC_565_0 ( .a(FE_RN_171_0), .b(FE_RN_172_0), .o(FE_RN_173_0) );
in01f80 g774579 ( .a(n_6556), .o(n_6676) );
ms00f80 delay_sub_ln23_0_unr1_stage2_stallmux_q_reg_1_ ( .ck(newNet_1660), .d(n_600), .o(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_) );
oa12f80 g765867 ( .a(n_15000), .b(n_14999), .c(n_14998), .o(n_15065) );
in01f80 g758060 ( .a(n_22880), .o(n_22881) );
na02f80 g777879 ( .a(n_3112), .b(n_2736), .o(n_3212) );
na02f80 FE_RC_4138_0 ( .a(FE_OCP_RBN3802_n_44721), .b(n_44365), .o(n_16900) );
no02f80 FE_RC_2705_0 ( .a(FE_OCP_RBN3466_n_7886), .b(n_8385), .o(FE_RN_1137_0) );
na02f80 g737007 ( .a(n_43230), .b(n_43001), .o(n_43500) );
in01f80 g775559 ( .a(n_5622), .o(n_5755) );
no02f80 g747481 ( .a(FE_OCP_RBN3333_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .o(n_32731) );
no03m80 FE_RC_3889_0 ( .a(n_28095), .b(n_28096), .c(n_28092), .o(n_28117) );
in01f80 g745838 ( .a(n_34238), .o(n_34256) );
in01f80 FE_OCP_RBC3389_n_33108 ( .a(FE_OCP_RBN3388_n_33108), .o(FE_OCP_RBN3389_n_33108) );
in01f80 g771037 ( .a(n_9668), .o(n_9669) );
no02f80 g758072 ( .a(n_22468), .b(FE_OCP_RBN1710_n_22150), .o(n_22469) );
na02f80 g775201 ( .a(n_5896), .b(n_5620), .o(n_5953) );
no02f80 g778706 ( .a(n_2365), .b(n_2364), .o(n_2383) );
no02f80 g737770 ( .a(n_42221), .b(n_42220), .o(n_42237) );
in01f80 newInst_2980 ( .a(newNet_2979), .o(newNet_2980) );
no02f80 g776162 ( .a(n_4652), .b(n_3082), .o(n_4848) );
na02f80 g747349 ( .a(n_33577), .b(n_33579), .o(n_33627) );
na02f80 g769922 ( .a(n_10974), .b(FE_OCP_RBN3643_n_44490), .o(n_11122) );
na02f80 g766347 ( .a(n_14360), .b(n_14361), .o(n_14460) );
oa12f80 g765178 ( .a(n_16345), .b(n_16344), .c(FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_16409) );
na02f80 g767974 ( .a(n_12775), .b(n_12994), .o(n_13425) );
na02f80 g755301 ( .a(n_24900), .b(n_24729), .o(n_24921) );
in01f80 g745175 ( .a(n_35554), .o(n_34893) );
na02f80 g781242 ( .a(n_158), .b(n_103), .o(n_141) );
na02f80 g744783 ( .a(n_35145), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35150) );
no02f80 g750592 ( .a(n_29423), .b(n_29404), .o(n_29527) );
no02f80 FE_RC_2480_0 ( .a(FE_RN_1000_0), .b(n_40468), .o(n_40495) );
na02f80 g778774 ( .a(n_2222), .b(n_2221), .o(n_2223) );
in01f80 g772056 ( .a(n_8747), .o(n_8694) );
na03f80 FE_RC_3292_0 ( .a(n_22634), .b(n_22769), .c(n_22714), .o(n_22822) );
no02f80 g746979 ( .a(FE_OCP_RBN2167_n_32892), .b(n_32991), .o(n_32992) );
no02f80 g746533 ( .a(n_35070), .b(n_34637), .o(n_35279) );
in01f80 newInst_928 ( .a(newNet_927), .o(newNet_928) );
na02f80 g776375 ( .a(n_4720), .b(n_4719), .o(n_4787) );
in01f80 g745300 ( .a(n_36219), .o(n_36220) );
in01f80 fopt783668 ( .a(n_45319), .o(n_45318) );
no02f80 g765860 ( .a(n_14827), .b(n_14861), .o(n_14921) );
na02f80 g759271 ( .a(n_20866), .b(n_20831), .o(n_20949) );
in01f80 g739920 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n_40341) );
no02f80 FE_RC_2923_0 ( .a(n_25757), .b(n_25789), .o(FE_RN_1272_0) );
na02f80 g775511 ( .a(n_5624), .b(n_5616), .o(n_5617) );
no02f80 g738832 ( .a(n_41295), .b(n_40987), .o(n_41327) );
na02f80 g762373 ( .a(n_45118), .b(n_18529), .o(n_18575) );
oa12f80 g755383 ( .a(n_25574), .b(n_25573), .c(n_25572), .o(n_26348) );
in01f80 FE_OCP_RBC3446_n_37945 ( .a(FE_OCP_RBN3443_n_37945), .o(FE_OCP_RBN3446_n_37945) );
no02f80 g745635 ( .a(n_34287), .b(n_34244), .o(n_34342) );
in01f80 g767502 ( .a(n_13009), .o(n_13059) );
in01f80 g754831 ( .a(n_25952), .o(n_25953) );
in01f80 newInst_3255 ( .a(newNet_1279), .o(newNet_3255) );
in01f80 g774778 ( .a(n_6456), .o(n_6457) );
no02f80 g770133 ( .a(n_10676), .b(FE_OCP_RBN3637_n_44490), .o(n_10704) );
oa12f80 g780089 ( .a(n_1172), .b(n_1184), .c(n_1171), .o(n_1187) );
na02f80 g780813 ( .a(n_504), .b(n_420), .o(n_513) );
na02f80 g771534 ( .a(FE_OCP_RBN2612_n_9075), .b(FE_OCP_RBN3556_n_44575), .o(n_9153) );
in01f80 FE_OCP_RBC2655_n_9198 ( .a(n_9198), .o(FE_OCP_RBN2655_n_9198) );
na02f80 g753772 ( .a(n_26463), .b(n_26518), .o(n_26594) );
ao22s80 FE_RC_3909_0 ( .a(n_16324), .b(n_16291), .c(n_16287), .d(n_16325), .o(n_16474) );
na02f80 g779576 ( .a(n_1362), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1467) );
ao22s80 FE_RC_2857_0 ( .a(n_13418), .b(n_14072), .c(n_13514), .d(FE_OCP_RBN2434_n_14072), .o(n_14177) );
in01f80 g746971 ( .a(n_32959), .o(n_32996) );
in01f80 g756278 ( .a(n_24121), .o(n_24137) );
na02f80 g770041 ( .a(n_10933), .b(n_10930), .o(n_10988) );
in01f80 g736368 ( .a(n_43788), .o(n_43833) );
in01f80 g773524 ( .a(n_8406), .o(n_7464) );
no02f80 g762079 ( .a(FE_OCP_RBN2203_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_22_), .o(n_18356) );
in01f80 g737641 ( .a(n_42799), .o(n_42800) );
no02f80 g750408 ( .a(n_30551), .b(n_30098), .o(n_30663) );
in01f80 g738035 ( .a(n_42156), .o(n_42157) );
in01f80 newInst_1225 ( .a(newNet_1148), .o(newNet_1225) );
in01f80 FE_RC_499_0 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_9_), .o(FE_RN_150_0) );
in01f80 g740710 ( .a(n_46949), .o(n_39965) );
in01f80 newInst_1901 ( .a(newNet_1900), .o(newNet_1901) );
in01f80 newInst_199 ( .a(newNet_198), .o(newNet_199) );
in01f80 FE_OCP_RBC3488_n_3390 ( .a(n_3390), .o(FE_OCP_RBN3488_n_3390) );
in01f80 FE_OCP_RBC3570_n_9188 ( .a(n_9188), .o(FE_OCP_RBN3570_n_9188) );
na02f80 g776720 ( .a(n_4249), .b(n_4365), .o(n_4416) );
in01f80 FE_OCP_RBC2241_n_44881 ( .a(FE_OCP_RBN2239_n_44881), .o(FE_OCP_RBN2241_n_44881) );
na02f80 g739251 ( .a(n_40776), .b(n_40858), .o(n_40883) );
na02f80 g749799 ( .a(n_31536), .b(n_31144), .o(n_31640) );
no02f80 g762186 ( .a(n_18167), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .o(n_18193) );
in01f80 g739295 ( .a(n_41038), .o(n_41039) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_4_ ( .ck(newNet_2245), .d(n_39958), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_) );
na02f80 g770500 ( .a(n_10394), .b(n_44490), .o(n_10473) );
oa22f80 g763709 ( .a(n_16757), .b(n_17336), .c(n_16725), .d(n_17753), .o(n_16804) );
na02f80 g778101 ( .a(n_2950), .b(FE_OCP_RBN3479_n_3006), .o(n_2979) );
no02f80 g742743 ( .a(n_37409), .b(n_36984), .o(n_37407) );
na02f80 g736974 ( .a(n_43242), .b(n_43300), .o(n_43455) );
ao12f80 g761159 ( .a(n_19989), .b(n_19907), .c(n_19845), .o(n_19990) );
in01f80 g777244 ( .a(n_3881), .o(n_3882) );
in01f80 g771719 ( .a(n_8842), .o(n_8828) );
in01f80 g772538 ( .a(n_8376), .o(n_8386) );
in01f80 FE_OCPC1520_n_31403 ( .a(FE_OCPN1519_n_31403), .o(FE_OCPN1520_n_31403) );
no02f80 g771285 ( .a(n_9787), .b(n_9699), .o(n_9923) );
in01f80 g773482 ( .a(n_7538), .o(n_7539) );
no02f80 g765885 ( .a(n_14814), .b(n_14215), .o(n_14855) );
ao12f80 g777051 ( .a(n_2798), .b(n_3484), .c(n_2663), .o(n_3561) );
na02f80 g751571 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_21_), .o(n_28545) );
in01f80 newInst_1971 ( .a(newNet_1892), .o(newNet_1971) );
ao12f80 g773012 ( .a(n_8113), .b(n_8032), .c(n_7886), .o(n_8143) );
na02f80 g765485 ( .a(n_15018), .b(n_14989), .o(n_15050) );
in01f80 fopt782983 ( .a(n_44453), .o(n_44454) );
oa12f80 g747774 ( .a(n_33293), .b(n_33571), .c(n_33279), .o(n_33841) );
no02f80 g738964 ( .a(n_41154), .b(n_40912), .o(n_41191) );
in01f80 FE_RC_3836_0 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .o(FE_RN_1672_0) );
in01f80 g759067 ( .a(n_21529), .o(n_21530) );
in01f80 newInst_1934 ( .a(newNet_1210), .o(newNet_1934) );
na02f80 g754817 ( .a(n_25949), .b(n_25290), .o(n_26106) );
na02f80 FE_RC_2753_0 ( .a(FE_RN_1168_0), .b(FE_RN_1170_0), .o(n_43874) );
no02f80 g745446 ( .a(n_35511), .b(n_34964), .o(n_35524) );
in01f80 newInst_842 ( .a(newNet_60), .o(newNet_842) );
na02f80 g776331 ( .a(n_4827), .b(n_4780), .o(n_4781) );
no02f80 g770426 ( .a(FE_OCP_RBN2925_n_10525), .b(n_10562), .o(n_10585) );
na02f80 FE_RC_2458_0 ( .a(FE_RN_983_0), .b(FE_RN_985_0), .o(n_13765) );
in01f80 g760181 ( .a(n_20658), .o(n_20659) );
na02f80 g759349 ( .a(n_20890), .b(n_20825), .o(n_20919) );
na02f80 g779797 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .o(n_1682) );
no02f80 g770925 ( .a(n_9753), .b(n_9759), .o(n_9944) );
na02f80 FE_RC_600_0 ( .a(n_25855), .b(FE_RN_188_0), .o(n_46962) );
in01f80 newInst_1443 ( .a(newNet_1442), .o(newNet_1443) );
na02f80 g737389 ( .a(n_46942), .b(n_42792), .o(n_42794) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_12_ ( .ck(newNet_2417), .d(n_36340), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_) );
ms00f80 cos_out_reg_14_ ( .ck(newNet_3745), .d(n_43818), .o(cos_out_14) );
in01f80 newInst_985 ( .a(newNet_984), .o(newNet_985) );
in01f80 g771651 ( .a(n_9102), .o(n_9103) );
oa22f80 FE_RC_3251_0 ( .a(n_21726), .b(n_21945), .c(n_21944), .d(n_21701), .o(n_22037) );
no02f80 g772680 ( .a(FE_OCP_RBN2428_n_8300), .b(n_8342), .o(n_8343) );
oa12f80 g752485 ( .a(n_27418), .b(n_27691), .c(n_27667), .o(n_27692) );
in01f80 g742759 ( .a(n_38235), .o(n_37452) );
na02f80 g766940 ( .a(n_14212), .b(n_14206), .o(n_14838) );
no02f80 g775926 ( .a(n_5275), .b(n_5353), .o(n_5616) );
in01f80 g737921 ( .a(n_42328), .o(n_42300) );
ao12f80 g757174 ( .a(n_23534), .b(n_23533), .c(n_23532), .o(n_24087) );
in01f80 g762116 ( .a(n_18883), .o(n_18930) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_5_ ( .ck(newNet_947), .d(n_22742), .o(delay_xor_ln21_unr15_stage6_stallmux_q_5_) );
oa22f80 g779225 ( .a(n_1889), .b(n_1650), .c(n_1872), .d(n_1649), .o(n_1938) );
na02f80 g743389 ( .a(n_36717), .b(n_36688), .o(n_36733) );
in01f80 newInst_156 ( .a(newNet_155), .o(newNet_156) );
in01f80 g744068 ( .a(n_47267), .o(n_36007) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_13_ ( .ck(newNet_192), .d(n_46363), .o(delay_xor_ln22_unr9_stage4_stallmux_q_13_) );
na02f80 g737057 ( .a(n_43046), .b(n_42956), .o(n_43126) );
oa12f80 g778360 ( .a(n_2478), .b(n_2508), .c(n_2477), .o(n_3902) );
na02f80 g737390 ( .a(n_42782), .b(n_42466), .o(n_42783) );
in01f80 g755188 ( .a(n_25098), .o(n_25099) );
in01f80 newInst_1200 ( .a(newNet_1199), .o(newNet_1200) );
ao12f80 g751337 ( .a(n_29464), .b(n_29463), .c(n_29462), .o(n_29938) );
no02f80 g740921 ( .a(n_39258), .b(n_39103), .o(n_39259) );
in01f80 g758603 ( .a(n_22527), .o(n_22528) );
no02f80 g760590 ( .a(n_19859), .b(n_19815), .o(n_19884) );
no02f80 g777792 ( .a(n_3288), .b(n_2437), .o(n_3324) );
na02f80 g766765 ( .a(n_13803), .b(n_13827), .o(n_13804) );
oa12f80 g740694 ( .a(n_39210), .b(n_39450), .c(n_39155), .o(n_39479) );
ao12f80 g773932 ( .a(n_6971), .b(n_6970), .c(n_6984), .o(n_7874) );
na02f80 g758307 ( .a(n_22288), .b(n_21226), .o(n_22463) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_4_ ( .ck(newNet_699), .d(n_46146), .o(delay_xor_ln21_unr6_stage3_stallmux_q_4_) );
oa22f80 g744996 ( .a(n_36314), .b(n_36159), .c(n_36313), .d(n_36160), .o(n_36384) );
in01f80 g747290 ( .a(n_34645), .o(n_33685) );
in01f80 g778230 ( .a(n_2826), .o(n_2827) );
in01f80 g759055 ( .a(n_21630), .o(n_21631) );
na02f80 g773747 ( .a(n_7220), .b(n_7081), .o(n_7284) );
oa12f80 g771095 ( .a(n_9492), .b(n_9553), .c(n_9552), .o(n_9628) );
in01f80 newInst_142 ( .a(newNet_117), .o(newNet_142) );
na02f80 g745520 ( .a(n_34351), .b(n_34350), .o(n_34352) );
ao12f80 g759481 ( .a(FE_OCP_RBN1359_FE_RN_677_0), .b(FE_OCP_RBN1217_n_20595), .c(n_20374), .o(n_20653) );
na02f80 g761786 ( .a(n_19160), .b(n_19159), .o(n_19161) );
no02f80 g748344 ( .a(n_31731), .b(n_31762), .o(n_31831) );
in01f80 g753524 ( .a(n_26822), .o(n_26823) );
na02f80 g747198 ( .a(n_33818), .b(n_33557), .o(n_33888) );
in01f80 newInst_3412 ( .a(newNet_3411), .o(newNet_3412) );
na02f80 g746600 ( .a(FE_OCP_RBN2598_n_34388), .b(n_34611), .o(n_34697) );
na02f80 g745444 ( .a(n_34436), .b(n_34450), .o(n_34489) );
in01f80 g738473 ( .a(n_41808), .o(n_41809) );
na02f80 g760462 ( .a(n_20078), .b(n_20073), .o(n_20074) );
na02f80 g765145 ( .a(n_16175), .b(n_15874), .o(n_16258) );
in01f80 g766497 ( .a(n_14146), .o(n_14147) );
in01f80 FE_OCP_RBC3575_n_4528 ( .a(n_4528), .o(FE_OCP_RBN3575_n_4528) );
na02f80 g740427 ( .a(FE_OCP_RBN3029_n_39942), .b(n_39558), .o(n_40166) );
oa12f80 g737857 ( .a(n_42577), .b(FE_OCPN1231_n_42201), .c(n_42276), .o(n_42620) );
no02f80 g754537 ( .a(n_26550), .b(n_26551), .o(n_26552) );
in01f80 g747762 ( .a(n_32277), .o(n_32278) );
in01f80 g762761 ( .a(n_17834), .o(n_17803) );
in01f80 g748382 ( .a(n_31475), .o(n_31610) );
oa22f80 g737215 ( .a(n_42940), .b(n_42677), .c(n_42975), .d(n_42678), .o(n_42990) );
oa12f80 g757884 ( .a(n_21954), .b(n_22088), .c(n_21941), .o(n_22205) );
in01f80 FE_OCP_RBC2710_n_35075 ( .a(n_35075), .o(FE_OCP_RBN2710_n_35075) );
no02f80 g742145 ( .a(n_37900), .b(n_37546), .o(n_38063) );
in01f80 g771481 ( .a(n_9208), .o(n_9288) );
oa12f80 g753698 ( .a(n_26461), .b(n_26525), .c(n_26392), .o(n_26623) );
na02f80 g747475 ( .a(n_32351), .b(n_44962), .o(n_32433) );
in01f80 newInst_2608 ( .a(newNet_2607), .o(newNet_2608) );
in01f80 g757284 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .o(n_23004) );
no02f80 g747957 ( .a(n_33116), .b(n_33115), .o(n_33117) );
na02f80 g738443 ( .a(n_41745), .b(n_41691), .o(n_41766) );
in01f80 newInst_1505 ( .a(newNet_1504), .o(newNet_1505) );
no02f80 g778186 ( .a(n_2843), .b(n_2680), .o(n_2885) );
na02f80 g764750 ( .a(n_16029), .b(n_16027), .o(n_16028) );
ao12f80 g752686 ( .a(n_27183), .b(n_27245), .c(n_27153), .o(n_27404) );
oa12f80 g745033 ( .a(n_34380), .b(n_34873), .c(n_34852), .o(n_34874) );
na02f80 g773732 ( .a(n_7225), .b(n_45844), .o(n_7227) );
na02f80 g773583 ( .a(n_7409), .b(n_7408), .o(n_7410) );
in01f80 g771969 ( .a(n_9876), .o(n_9827) );
oa12f80 g759564 ( .a(FE_OCP_RBN3677_n_21051), .b(n_21881), .c(n_21454), .o(n_21455) );
na02f80 g750702 ( .a(n_29279), .b(n_28827), .o(n_29276) );
in01f80 FE_OCP_RBC2051_delay_xor_ln22_unr15_stage6_stallmux_q_2_ ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .o(FE_OCP_RBN2051_delay_xor_ln22_unr15_stage6_stallmux_q_2_) );
na02f80 g765923 ( .a(n_14748), .b(n_14801), .o(n_14856) );
in01f80 g756066 ( .a(n_24336), .o(n_24491) );
na02f80 g748328 ( .a(n_31765), .b(n_30300), .o(n_31766) );
na02f80 g755420 ( .a(n_24867), .b(n_24853), .o(n_24963) );
na02f80 g763515 ( .a(FE_OCP_RBN3082_n_16977), .b(n_16011), .o(n_17167) );
no02f80 g752243 ( .a(n_28538), .b(n_28195), .o(n_28586) );
no02f80 g757846 ( .a(n_22983), .b(n_22765), .o(n_23027) );
in01f80 fopt783563 ( .a(n_45145), .o(n_45180) );
in01f80 newInst_1080 ( .a(newNet_900), .o(newNet_1080) );
in01f80 g749266 ( .a(n_32152), .o(n_32153) );
na02f80 g759172 ( .a(n_21046), .b(n_45091), .o(n_21192) );
no02f80 g745540 ( .a(n_34704), .b(n_34993), .o(n_34624) );
no02f80 g761905 ( .a(n_18302), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .o(n_18321) );
ao12f80 g754747 ( .a(n_25337), .b(n_25336), .c(n_25335), .o(n_26966) );
no02f80 g739421 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n_40825) );
oa12f80 g775365 ( .a(n_5875), .b(n_5874), .c(n_5873), .o(n_5929) );
oa22f80 g758777 ( .a(n_21580), .b(n_21612), .c(n_21579), .d(n_21679), .o(n_21706) );
in01f80 g745857 ( .a(n_35390), .o(n_35406) );
in01f80 FE_RC_3674_0 ( .a(FE_OCPN1411_n_21007), .o(FE_RN_1614_0) );
na02f80 g756411 ( .a(n_23928), .b(n_23972), .o(n_24014) );
in01f80 FE_OCPC1790_n_18119 ( .a(FE_OCPN1789_n_18119), .o(FE_OCPN1790_n_18119) );
in01f80 newInst_3365 ( .a(newNet_3364), .o(newNet_3365) );
in01f80 newInst_1602 ( .a(newNet_1601), .o(newNet_1602) );
no02f80 g740511 ( .a(n_39746), .b(n_39745), .o(n_39758) );
na02f80 g766653 ( .a(FE_OCP_RBN3477_n_13756), .b(FE_OCP_RBN2243_n_13017), .o(n_13817) );
in01f80 g749813 ( .a(n_31619), .o(n_31620) );
ao12f80 g743229 ( .a(n_38045), .b(n_38044), .c(n_46242), .o(n_38128) );
in01f80 g743035 ( .a(n_37180), .o(n_37181) );
in01f80 FE_RC_971_0 ( .a(n_26181), .o(FE_RN_280_0) );
in01f80 FE_OCPC899_n_44593 ( .a(FE_OCP_RBN3554_n_44575), .o(FE_OCPN899_n_44593) );
no02f80 g772965 ( .a(n_7927), .b(n_7818), .o(n_8009) );
no02f80 g755804 ( .a(n_24429), .b(n_22089), .o(n_24519) );
in01f80 g739302 ( .a(n_40971), .o(n_40972) );
in01f80 g752784 ( .a(n_27905), .o(n_27906) );
in01f80 g740264 ( .a(n_40173), .o(n_40174) );
na02f80 g763680 ( .a(n_17367), .b(n_17098), .o(n_17369) );
na02f80 g749332 ( .a(n_30586), .b(n_30566), .o(n_30747) );
in01f80 g743223 ( .a(n_36846), .o(n_36889) );
na02f80 g780328 ( .a(n_942), .b(n_850), .o(n_1046) );
na02f80 g767799 ( .a(n_12863), .b(n_12821), .o(n_12822) );
ao22s80 FE_RC_825_0 ( .a(n_8543), .b(n_8567), .c(n_8542), .d(n_8566), .o(n_8687) );
in01f80 g763335 ( .a(n_17130), .o(n_17131) );
oa12f80 g758707 ( .a(n_21698), .b(n_22284), .c(n_21722), .o(n_22396) );
no02f80 g767902 ( .a(n_13889), .b(n_11944), .o(n_12768) );
in01f80 g773717 ( .a(n_7281), .o(n_7282) );
na02f80 g743290 ( .a(n_36756), .b(n_36724), .o(n_36769) );
oa22f80 g742483 ( .a(n_37595), .b(n_36686), .c(n_37620), .d(n_37625), .o(n_38685) );
no02f80 g751755 ( .a(n_28309), .b(n_28015), .o(n_28334) );
no02f80 g736614 ( .a(n_43646), .b(n_43406), .o(n_43641) );
no02f80 g742049 ( .a(n_37900), .b(n_37948), .o(n_38057) );
na02f80 g752812 ( .a(n_27879), .b(n_27926), .o(n_28244) );
in01f80 fopt784718 ( .a(n_47200), .o(n_47199) );
na02f80 g773463 ( .a(n_7560), .b(n_7146), .o(n_7561) );
oa12f80 g749415 ( .a(n_30217), .b(FE_OCP_RBN2755_n_30558), .c(n_30577), .o(n_30605) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_25_ ( .ck(newNet_3407), .d(n_27800), .o(delay_add_ln22_unr17_stage7_stallmux_q_25_) );
no02f80 g756598 ( .a(n_23606), .b(n_23658), .o(n_23740) );
no02f80 g774504 ( .a(n_6524), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_), .o(n_6593) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_24_ ( .ck(newNet_1221), .d(n_6085), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_) );
in01f80 g756382 ( .a(n_23887), .o(n_23888) );
in01f80 FE_OCP_RBC3582_n_44944 ( .a(FE_OCP_RBN2545_n_44944), .o(FE_OCP_RBN3582_n_44944) );
no02f80 FE_RC_1399_0 ( .a(n_15856), .b(n_15942), .o(FE_RN_408_0) );
oa12f80 g740998 ( .a(n_38970), .b(n_38969), .c(n_38968), .o(n_39084) );
no03m80 FE_RC_339_0 ( .a(n_12071), .b(n_11796), .c(n_12108), .o(n_12234) );
in01f80 FE_RC_2653_0 ( .a(n_12581), .o(FE_RN_1107_0) );
na02f80 g771992 ( .a(FE_OCPN903_n_44581), .b(n_9223), .o(n_9380) );
no02f80 g766596 ( .a(n_14016), .b(n_13909), .o(n_14087) );
na02f80 g772024 ( .a(n_8783), .b(n_8055), .o(n_8887) );
in01f80 g765877 ( .a(n_14919), .o(n_14920) );
in01f80 FE_OCP_RBC2726_n_4219 ( .a(FE_OCP_RBN2723_n_4219), .o(FE_OCP_RBN2726_n_4219) );
in01f80 g744002 ( .a(n_36301), .o(n_36302) );
oa12f80 g759826 ( .a(n_21252), .b(n_21714), .c(n_21169), .o(n_21887) );
in01f80 FE_RC_1831_0 ( .a(n_13992), .o(FE_RN_550_0) );
na02f80 g743592 ( .a(n_36484), .b(n_36307), .o(n_36529) );
in01f80 g752613 ( .a(n_27614), .o(n_27615) );
oa22f80 g774530 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln23_unr6_stage3_stallmux_q), .c(FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(FE_OCP_RBN1988_delay_xor_ln23_unr6_stage3_stallmux_q), .o(n_6528) );
ao12f80 g742935 ( .a(n_37001), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n_37325) );
na02f80 g770365 ( .a(FE_OCP_RBN3691_n_10567), .b(n_10609), .o(n_10639) );
no02f80 g747375 ( .a(n_32389), .b(n_44962), .o(n_32438) );
no02f80 g751064 ( .a(n_30091), .b(n_30088), .o(n_30951) );
na02f80 g778510 ( .a(n_2342), .b(n_1933), .o(n_2356) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_31_ ( .ck(newNet_3114), .d(n_40592), .o(delay_add_ln22_unr27_stage10_stallmux_q_31_) );
ao22s80 FE_RC_3455_0 ( .a(n_20310), .b(FE_OCP_RBN1841_n_20505), .c(n_20505), .d(n_20312), .o(n_20640) );
no02f80 g758588 ( .a(n_22037), .b(n_22036), .o(n_22063) );
oa12f80 g760499 ( .a(n_19941), .b(n_20007), .c(n_19880), .o(n_20026) );
in01f80 g777933 ( .a(n_3169), .o(n_3170) );
in01f80 newInst_2349 ( .a(newNet_2348), .o(newNet_2349) );
no02f80 g764458 ( .a(n_16084), .b(n_16191), .o(n_16192) );
oa12f80 g752700 ( .a(n_27243), .b(n_27244), .c(n_27151), .o(n_27313) );
ao12f80 g737453 ( .a(n_42545), .b(n_42639), .c(n_42582), .o(n_42671) );
na02f80 g777088 ( .a(n_3690), .b(n_3733), .o(n_3886) );
in01f80 FE_OCP_RBC2437_n_8402 ( .a(n_8402), .o(FE_OCP_RBN2437_n_8402) );
no02f80 FE_RC_1318_0 ( .a(FE_RN_387_0), .b(FE_RN_388_0), .o(FE_RN_389_0) );
na02f80 g778625 ( .a(n_2391), .b(n_2452), .o(n_3044) );
in01f80 g758399 ( .a(n_23486), .o(n_23590) );
in01f80 g764705 ( .a(n_15942), .o(n_15984) );
in01f80 g758385 ( .a(FE_OCPN1494_n_23398), .o(n_23414) );
in01f80 newInst_423 ( .a(newNet_422), .o(newNet_423) );
in01f80 FE_OCP_RBC1716_n_20734 ( .a(FE_OCP_RBN1715_n_20734), .o(FE_OCP_RBN1716_n_20734) );
in01f80 g775267 ( .a(n_5818), .o(n_5800) );
in01f80 g776705 ( .a(n_4245), .o(n_4246) );
in01f80 FE_OCP_RBC3466_n_7886 ( .a(FE_OCP_RBN3459_n_7886), .o(FE_OCP_RBN3466_n_7886) );
na02f80 g757385 ( .a(n_22995), .b(n_22994), .o(n_22996) );
in01f80 g756768 ( .a(n_23496), .o(n_23497) );
na02f80 g765011 ( .a(n_15529), .b(n_15580), .o(n_15676) );
ao22s80 FE_RC_3269_0 ( .a(n_11388), .b(n_11413), .c(n_11389), .d(FE_OCP_RBN3095_n_11413), .o(n_11527) );
oa12f80 g761708 ( .a(n_19402), .b(n_19401), .c(n_18739), .o(n_19489) );
in01f80 g750832 ( .a(n_29143), .o(n_29161) );
in01f80 newInst_1274 ( .a(newNet_1230), .o(newNet_1274) );
in01f80 g775156 ( .a(n_6039), .o(n_6040) );
in01f80 newInst_1381 ( .a(newNet_1380), .o(newNet_1381) );
na02f80 g742042 ( .a(n_38136), .b(n_38163), .o(n_38214) );
in01f80 newInst_1051 ( .a(newNet_1050), .o(newNet_1051) );
na02f80 g768460 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_21_), .o(n_12390) );
no02f80 g738314 ( .a(n_41648), .b(n_41820), .o(n_41822) );
in01f80 g764224 ( .a(n_16552), .o(n_16576) );
in01f80 g748067 ( .a(n_32026), .o(n_32027) );
in01f80 g745420 ( .a(n_35630), .o(n_35722) );
no02f80 g753462 ( .a(n_26806), .b(n_26827), .o(n_26967) );
na02f80 g765292 ( .a(n_15919), .b(n_16018), .o(n_16060) );
no02f80 g740047 ( .a(n_39982), .b(n_39905), .o(n_39906) );
in01f80 g742298 ( .a(n_37973), .o(n_38007) );
ao12f80 g764762 ( .a(n_15270), .b(n_45137), .c(n_15272), .o(n_15660) );
in01f80 g744243 ( .a(n_36868), .o(n_36869) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_14_ ( .ck(newNet_2782), .d(n_16699), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_) );
in01f80 newInst_3595 ( .a(newNet_3594), .o(newNet_3595) );
ms00f80 delay_sub_ln23_unr9_stage4_stallmux_q_reg_2_ ( .ck(newNet_1046), .d(FE_OFN800_n_46285), .o(delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
na02f80 g775622 ( .a(n_5267), .b(n_5358), .o(n_5377) );
na02f80 g751771 ( .a(n_28931), .b(n_28993), .o(n_28962) );
na02f80 g771523 ( .a(n_9078), .b(n_9189), .o(n_9245) );
in01f80 g740964 ( .a(n_39165), .o(n_39194) );
no02f80 g767566 ( .a(n_13239), .b(n_12924), .o(n_13382) );
na02f80 g751941 ( .a(n_28125), .b(n_28124), .o(n_28187) );
in01f80 newInst_3142 ( .a(newNet_3141), .o(newNet_3142) );
ao12f80 g774059 ( .a(n_6803), .b(n_6835), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n_6897) );
no02f80 g751980 ( .a(n_28897), .b(n_28327), .o(n_29170) );
in01f80 g765325 ( .a(FE_OCP_RBN2738_n_15300), .o(n_15336) );
oa12f80 g745207 ( .a(n_34136), .b(n_34415), .c(n_34414), .o(n_34494) );
no02f80 FE_RC_4226_0 ( .a(FE_RN_1854_0), .b(FE_RN_1734_0), .o(FE_RN_1855_0) );
in01f80 g738738 ( .a(n_41529), .o(n_41850) );
oa12f80 g775886 ( .a(n_5158), .b(n_5157), .c(n_5156), .o(n_5323) );
ao12f80 g768777 ( .a(n_11677), .b(n_11958), .c(n_11459), .o(n_11959) );
no02f80 g752693 ( .a(n_27998), .b(n_27933), .o(n_28082) );
ao12f80 g741853 ( .a(n_38327), .b(n_38287), .c(n_38304), .o(n_38444) );
na02f80 g769245 ( .a(n_11582), .b(n_11464), .o(n_11674) );
na02f80 g755036 ( .a(n_25118), .b(n_25107), .o(n_25108) );
in01f80 g737407 ( .a(n_43106), .o(n_42805) );
na02f80 g759012 ( .a(n_22053), .b(n_22052), .o(n_22054) );
oa12f80 g744227 ( .a(n_35489), .b(n_35488), .c(n_35495), .o(n_35507) );
na02f80 g776195 ( .a(n_4954), .b(n_4953), .o(n_5052) );
in01f80 g773690 ( .a(n_7611), .o(n_8226) );
no02f80 g744518 ( .a(n_35384), .b(n_35232), .o(n_35411) );
no02f80 g765345 ( .a(n_15127), .b(n_15180), .o(n_15298) );
in01f80 g765366 ( .a(n_16304), .o(n_16305) );
oa12f80 g760443 ( .a(n_20560), .b(n_20559), .c(n_20558), .o(n_21481) );
in01f80 g748085 ( .a(n_32024), .o(n_32025) );
in01f80 newInst_2518 ( .a(newNet_2517), .o(newNet_2518) );
ao12f80 g767482 ( .a(n_12844), .b(n_13393), .c(n_12963), .o(n_13474) );
no02f80 g749781 ( .a(n_31368), .b(n_31324), .o(n_31388) );
na02f80 g736935 ( .a(n_43242), .b(n_42805), .o(n_43461) );
na02f80 g768299 ( .a(n_12532), .b(n_12517), .o(n_12565) );
no03m80 FE_RC_4224_0 ( .a(n_29960), .b(n_29958), .c(n_29915), .o(FE_RN_1853_0) );
in01f80 g750532 ( .a(n_29479), .o(n_29530) );
in01f80 g744452 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_), .o(n_35473) );
in01f80 g736646 ( .a(n_43479), .o(n_43480) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_8_ ( .ck(newNet_3361), .d(n_26969), .o(delay_add_ln22_unr17_stage7_stallmux_q_8_) );
in01f80 g763573 ( .a(n_16868), .o(n_16869) );
oa12f80 g763046 ( .a(n_17636), .b(n_17635), .c(n_17634), .o(n_19010) );
oa22f80 g744527 ( .a(n_36644), .b(n_36211), .c(n_36645), .d(n_36212), .o(n_36700) );
no02f80 g768746 ( .a(n_12129), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .o(n_12182) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_20_ ( .ck(newNet_3051), .d(FE_RN_1424_0), .o(delay_add_ln22_unr2_stage2_stallmux_q_20_) );
in01f80 g760152 ( .a(n_20778), .o(n_20664) );
na02f80 g741056 ( .a(n_38985), .b(n_38917), .o(n_39055) );
no02f80 g780579 ( .a(n_666), .b(n_563), .o(n_705) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_26_ ( .ck(newNet_3299), .d(FE_OCP_RBN3129_n_32266), .o(delay_add_ln22_unr20_stage8_stallmux_q_26_) );
no02f80 FE_RC_2486_0 ( .a(FE_RN_1004_0), .b(n_10422), .o(FE_RN_1005_0) );
in01f80 g736885 ( .a(n_43595), .o(n_43596) );
in01f80 FE_RC_564_0 ( .a(FE_RN_173_0), .o(n_31742) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_30_ ( .ck(newNet_3601), .d(n_17812), .o(delay_add_ln22_unr11_stage5_stallmux_q_30_) );
na02f80 g738743 ( .a(n_41564), .b(n_41366), .o(n_41715) );
no02f80 g737442 ( .a(n_42687), .b(n_42681), .o(n_42704) );
no02f80 g739100 ( .a(n_41048), .b(n_40845), .o(n_41049) );
no02f80 g775253 ( .a(n_5867), .b(n_5809), .o(n_5938) );
no02f80 g765518 ( .a(n_15565), .b(n_15786), .o(n_15667) );
ao22s80 FE_RC_878_0 ( .a(n_10320), .b(n_10317), .c(n_10318), .d(n_10321), .o(n_10480) );
no02f80 g752967 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(n_28326) );
oa12f80 g750984 ( .a(n_28887), .b(n_28933), .c(n_28842), .o(n_28971) );
na02f80 g743382 ( .a(n_36592), .b(n_36750), .o(n_36593) );
ao12f80 g760630 ( .a(n_20083), .b(n_20277), .c(n_20113), .o(n_20329) );
no02f80 g757061 ( .a(n_23616), .b(n_22886), .o(n_23617) );
ao12f80 g745081 ( .a(n_34825), .b(n_34824), .c(n_34823), .o(n_35611) );
oa12f80 g770659 ( .a(n_10164), .b(n_10353), .c(n_10083), .o(n_10431) );
in01f80 FE_OCP_RBC2659_n_4101 ( .a(n_4101), .o(FE_OCP_RBN2659_n_4101) );
no02f80 g746747 ( .a(n_33185), .b(n_33155), .o(n_33218) );
in01f80 g740180 ( .a(n_39977), .o(n_40072) );
ao22s80 FE_RC_845_0 ( .a(n_9550), .b(n_9583), .c(n_9551), .d(n_9626), .o(n_9819) );
no02f80 g742137 ( .a(n_38272), .b(n_38248), .o(n_38385) );
na02f80 g750066 ( .a(n_29869), .b(n_29161), .o(n_30077) );
no02f80 g741452 ( .a(n_38803), .b(n_38813), .o(n_38844) );
in01f80 g752716 ( .a(n_27244), .o(n_27241) );
no02f80 g746918 ( .a(FE_OCP_RBN3385_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n_33149) );
in01f80 g742648 ( .a(n_37459), .o(n_37460) );
ao12f80 g736418 ( .a(n_43443), .b(n_43721), .c(n_43514), .o(n_43747) );
oa12f80 g769616 ( .a(n_10250), .b(n_11333), .c(n_10341), .o(n_11384) );
ao12f80 g738287 ( .a(n_41840), .b(n_41839), .c(n_41838), .o(n_42212) );
na02f80 g744890 ( .a(n_35077), .b(n_30587), .o(n_35136) );
no02f80 g748706 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_), .o(n_32559) );
na02f80 g761165 ( .a(n_19046), .b(n_19058), .o(n_19112) );
in01f80 g759628 ( .a(n_20790), .o(n_20791) );
no02f80 g747711 ( .a(n_32264), .b(n_31993), .o(n_32265) );
in01f80 newInst_1032 ( .a(newNet_1031), .o(newNet_1032) );
in01f80 newInst_2477 ( .a(newNet_2476), .o(newNet_2477) );
no02f80 g769074 ( .a(n_11602), .b(n_11686), .o(n_11687) );
no02f80 FE_RC_3383_0 ( .a(n_13004), .b(FE_OCP_RBN2206_n_12907), .o(FE_RN_1466_0) );
no02f80 g756020 ( .a(n_25032), .b(n_24767), .o(n_25193) );
oa12f80 g784684 ( .a(n_3683), .b(n_3575), .c(n_3460), .o(n_47014) );
na02f80 g751372 ( .a(n_29362), .b(n_28946), .o(n_29457) );
no02f80 g751731 ( .a(n_44143), .b(n_28065), .o(n_28385) );
no02f80 g762874 ( .a(n_17656), .b(n_17655), .o(n_17827) );
na02f80 g777910 ( .a(n_3055), .b(n_3159), .o(n_3174) );
in01f80 g772374 ( .a(n_8574), .o(n_8575) );
na02f80 g779157 ( .a(n_2007), .b(n_2006), .o(n_2221) );
in01f80 g769852 ( .a(FE_OCP_RBN2998_n_11004), .o(n_11031) );
na02f80 g742838 ( .a(n_37253), .b(n_37161), .o(n_37254) );
na02f80 g753210 ( .a(n_27207), .b(n_26114), .o(n_27387) );
in01f80 g763502 ( .a(n_16837), .o(n_16874) );
in01f80 FE_OCP_RBC3124_n_6557 ( .a(n_6557), .o(FE_OCP_RBN3124_n_6557) );
ao12f80 g762658 ( .a(n_18052), .b(FE_OCP_RBN2142_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .o(n_17970) );
na02f80 FE_RC_3476_0 ( .a(n_35780), .b(n_35732), .o(FE_RN_1494_0) );
no02f80 g770688 ( .a(n_9896), .b(n_9862), .o(n_9935) );
in01f80 g737347 ( .a(n_42842), .o(n_42852) );
in01f80 g759255 ( .a(n_21203), .o(n_21216) );
no02f80 g749754 ( .a(n_30177), .b(n_30175), .o(n_30223) );
in01f80 g740199 ( .a(n_39907), .o(n_39862) );
in01f80 g753767 ( .a(n_26497), .o(n_26498) );
in01f80 newInst_2799 ( .a(newNet_2798), .o(newNet_2799) );
in01f80 g749651 ( .a(n_32076), .o(n_30326) );
in01f80 g772890 ( .a(n_7821), .o(n_7822) );
in01f80 g753251 ( .a(n_27143), .o(n_27173) );
no02f80 g770629 ( .a(n_10379), .b(FE_OCP_RBN3558_n_8687), .o(n_10380) );
in01f80 g740317 ( .a(n_39816), .o(n_39812) );
na02f80 g737944 ( .a(n_42270), .b(n_42152), .o(n_42351) );
in01f80 g771240 ( .a(n_9565), .o(n_9566) );
in01f80 newInst_1984 ( .a(newNet_1983), .o(newNet_1984) );
oa22f80 g755078 ( .a(n_25551), .b(n_24621), .c(n_25373), .d(n_24650), .o(n_25747) );
no02f80 g749029 ( .a(n_31026), .b(n_31025), .o(n_31027) );
na02f80 g765038 ( .a(n_15348), .b(n_15425), .o(n_15464) );
no02f80 g741010 ( .a(n_38932), .b(n_38966), .o(n_39016) );
in01f80 newInst_2146 ( .a(newNet_2145), .o(newNet_2146) );
in01f80 g738638 ( .a(n_41540), .o(n_41660) );
in01f80 newInst_1953 ( .a(newNet_1952), .o(newNet_1953) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_12_ ( .ck(newNet_2217), .d(n_1099), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_18_ ( .ck(newNet_1016), .d(n_17879), .o(delay_xor_ln21_unr12_stage5_stallmux_q_18_) );
no02f80 g751041 ( .a(n_29881), .b(n_29878), .o(n_29882) );
in01f80 g772981 ( .a(n_7861), .o(n_7862) );
in01f80 g745578 ( .a(n_34344), .o(n_34319) );
ao12f80 g736285 ( .a(n_43471), .b(n_43885), .c(n_43384), .o(n_43892) );
in01f80 g770013 ( .a(n_10962), .o(n_11007) );
no02f80 g750051 ( .a(n_29896), .b(n_30364), .o(n_30383) );
na02f80 g758764 ( .a(n_21871), .b(n_21808), .o(n_21893) );
in01f80 FE_RC_667_0 ( .a(n_36918), .o(FE_RN_211_0) );
no02f80 g745190 ( .a(n_34656), .b(n_34630), .o(n_34631) );
na02f80 g737010 ( .a(n_43230), .b(n_43010), .o(n_43499) );
in01f80 g766314 ( .a(n_14403), .o(n_14404) );
oa22f80 g745343 ( .a(n_35956), .b(n_35809), .c(FE_OCP_RBN2995_n_35539), .d(n_34671), .o(n_36225) );
na03f80 g742720 ( .a(n_37366), .b(n_37353), .c(n_37219), .o(n_37399) );
in01f80 g742656 ( .a(n_37499), .o(n_37520) );
no02f80 g741898 ( .a(n_38358), .b(n_38353), .o(n_38354) );
in01f80 FE_OCP_RBC1721_n_21004 ( .a(n_21004), .o(FE_OCP_RBN1721_n_21004) );
no02f80 g744038 ( .a(n_44223), .b(n_34540), .o(n_35751) );
oa22f80 g784365 ( .a(FE_OFN86_n_46137), .b(n_5937), .c(FE_OFN805_n_46196), .d(n_5972), .o(n_46171) );
in01f80 FE_RC_1101_0 ( .a(n_40494), .o(FE_RN_327_0) );
in01f80 g740907 ( .a(n_39460), .o(n_39840) );
in01f80 fopt783091 ( .a(n_44570), .o(n_44568) );
no02f80 g745946 ( .a(n_33969), .b(n_33968), .o(n_33985) );
no02f80 g762284 ( .a(n_18613), .b(n_18524), .o(n_19019) );
in01f80 newInst_3006 ( .a(newNet_3005), .o(newNet_3006) );
no02f80 g773427 ( .a(n_7584), .b(n_6680), .o(n_7585) );
no02f80 g737573 ( .a(n_42410), .b(n_42334), .o(n_42427) );
in01f80 FE_OCP_RBC1705_n_21658 ( .a(n_21658), .o(FE_OCP_RBN1705_n_21658) );
ao12f80 g779423 ( .a(n_1508), .b(n_1506), .c(n_1507), .o(n_1561) );
no02f80 g767281 ( .a(n_13436), .b(n_13429), .o(n_13512) );
oa22f80 FE_RC_4262_0 ( .a(n_32551), .b(n_32583), .c(n_32552), .d(n_32641), .o(n_32671) );
in01f80 FE_OCPC1521_n_26054 ( .a(n_26054), .o(FE_OCPN1521_n_26054) );
no02f80 g775443 ( .a(n_5685), .b(n_5596), .o(n_5785) );
in01f80 newInst_3023 ( .a(newNet_3022), .o(newNet_3023) );
no02f80 FE_RC_1784_0 ( .a(n_27923), .b(FE_RN_521_0), .o(FE_RN_522_0) );
na02f80 g755264 ( .a(n_25529), .b(n_25120), .o(n_25660) );
in01f80 FE_OCPUNCOC3143_n_19138 ( .a(n_19138), .o(FE_OCPUNCON3143_n_19138) );
in01f80 newInst_3019 ( .a(newNet_2919), .o(newNet_3019) );
na02f80 g775421 ( .a(n_5690), .b(n_5547), .o(n_5876) );
in01f80 FE_OCPC1480_n_23872 ( .a(FE_OCPN1479_n_23872), .o(FE_OCPN1480_n_23872) );
na02f80 g749023 ( .a(n_31049), .b(n_30930), .o(n_31096) );
in01f80 newInst_3236 ( .a(newNet_2466), .o(newNet_3236) );
oa12f80 g751812 ( .a(n_29126), .b(n_29123), .c(n_28897), .o(n_29804) );
oa12f80 g776935 ( .a(n_3511), .b(n_3572), .c(n_3459), .o(n_3724) );
ao12f80 g781176 ( .a(n_67), .b(n_174), .c(beta_31), .o(n_175) );
in01f80 newInst_3284 ( .a(newNet_570), .o(newNet_3284) );
in01f80 newInst_221 ( .a(newNet_58), .o(newNet_221) );
oa12f80 g771890 ( .a(n_8635), .b(n_45503), .c(n_8634), .o(n_8703) );
in01f80 FE_OCP_RBC3068_n_43230 ( .a(FE_OCP_RBN3067_n_43230), .o(FE_OCP_RBN3068_n_43230) );
in01f80 newInst_2228 ( .a(newNet_2227), .o(newNet_2228) );
no02f80 g775165 ( .a(n_5994), .b(n_5091), .o(n_5995) );
in01f80 g759962 ( .a(n_21295), .o(n_21296) );
in01f80 FE_RC_3209_0 ( .a(n_954), .o(FE_RN_1427_0) );
in01f80 g772457 ( .a(n_8517), .o(n_8573) );
na02f80 g762086 ( .a(n_18222), .b(n_18216), .o(n_18223) );
in01f80 FE_OCPC1000_n_45660 ( .a(FE_OCP_RBN2121_n_45224), .o(FE_OCPN1000_n_45660) );
ao12f80 g737334 ( .a(n_42450), .b(n_42854), .c(n_42464), .o(n_42881) );
no02f80 g750019 ( .a(n_30195), .b(n_30108), .o(n_30218) );
in01f80 g741236 ( .a(n_38915), .o(n_38916) );
no02f80 g765167 ( .a(n_15123), .b(n_15159), .o(n_15275) );
in01f80 g739244 ( .a(n_40921), .o(n_40922) );
in01f80 newInst_3392 ( .a(newNet_3391), .o(newNet_3392) );
na02f80 g753225 ( .a(n_27204), .b(FE_OCP_RBN3682_n_26171), .o(n_27340) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_13_ ( .ck(newNet_3336), .d(n_31998), .o(delay_add_ln22_unr20_stage8_stallmux_q_13_) );
in01f80 g767628 ( .a(n_13134), .o(n_13135) );
ao12f80 g741919 ( .a(n_38072), .b(n_38074), .c(n_38071), .o(n_38146) );
oa22f80 g779397 ( .a(n_1496), .b(n_1461), .c(n_1495), .d(n_1460), .o(n_1571) );
no02f80 g775656 ( .a(n_5130), .b(FE_OCP_RBN2727_n_4219), .o(n_5173) );
no02f80 g773993 ( .a(n_6800), .b(n_6841), .o(n_6914) );
in01f80 g772978 ( .a(n_7863), .o(n_7864) );
no02f80 g747746 ( .a(n_33990), .b(n_33970), .o(n_34332) );
na02f80 g736995 ( .a(n_43230), .b(n_43265), .o(n_43502) );
ao12f80 g742952 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37042), .c(n_36429), .o(n_37163) );
in01f80 FE_OCP_RBC2518_n_8762 ( .a(n_8762), .o(FE_OCP_RBN2518_n_8762) );
oa22f80 g780225 ( .a(n_1003), .b(n_1203), .c(n_969), .d(FE_OFN794_n_45813), .o(n_1102) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_12_ ( .ck(newNet_2879), .d(n_10959), .o(delay_add_ln22_unr8_stage4_stallmux_q_12_) );
in01f80 g775112 ( .a(n_5976), .o(n_5977) );
in01f80 g745539 ( .a(n_34624), .o(n_34625) );
na02f80 g769337 ( .a(n_9652), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11590) );
no02f80 g752282 ( .a(n_27913), .b(n_44735), .o(n_28032) );
na02f80 g736593 ( .a(n_43626), .b(n_43404), .o(n_43657) );
no02f80 g764681 ( .a(n_15946), .b(n_15905), .o(n_15987) );
in01f80 fopt783328 ( .a(n_44875), .o(n_44881) );
na02f80 g742233 ( .a(n_44867), .b(n_37493), .o(n_37928) );
oa12f80 g767493 ( .a(n_12640), .b(n_12948), .c(n_12622), .o(n_13097) );
no02f80 g759673 ( .a(n_20682), .b(n_20760), .o(n_20721) );
no02f80 FE_RC_2541_0 ( .a(FE_OCP_RBN2548_n_44944), .b(FE_RN_1037_0), .o(FE_RN_1038_0) );
in01f80 newInst_3530 ( .a(newNet_3529), .o(newNet_3530) );
oa12f80 g777947 ( .a(n_3046), .b(n_3045), .c(n_3044), .o(n_4537) );
in01f80 FE_RC_2686_0 ( .a(n_9012), .o(FE_RN_1124_0) );
in01f80 newInst_1312 ( .a(newNet_1311), .o(newNet_1312) );
na02f80 g778954 ( .a(n_2198), .b(delay_add_ln22_unr2_stage2_stallmux_q_19_), .o(n_2243) );
na02f80 g747831 ( .a(n_33392), .b(n_33354), .o(n_33601) );
in01f80 FE_RC_2489_0 ( .a(n_24067), .o(FE_RN_1007_0) );
oa12f80 g778408 ( .a(n_2395), .b(n_2419), .c(n_2394), .o(n_2495) );
ao12f80 g746858 ( .a(n_33159), .b(FE_OCP_RBN3390_n_33108), .c(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(n_33467) );
no02f80 g747698 ( .a(n_33318), .b(n_33315), .o(n_33394) );
no02f80 g777223 ( .a(n_3665), .b(n_3699), .o(n_3832) );
in01f80 g769350 ( .a(n_11709), .o(n_11710) );
no02f80 g740395 ( .a(FE_OCP_RBN3021_n_39942), .b(n_39910), .o(n_39912) );
in01f80 g759138 ( .a(n_21163), .o(n_22251) );
oa12f80 g738607 ( .a(n_41535), .b(n_41713), .c(n_41526), .o(n_41943) );
na02f80 g755598 ( .a(n_25310), .b(n_25345), .o(n_25408) );
na02f80 g744291 ( .a(FE_OCP_RBN2902_n_44174), .b(n_35023), .o(n_35814) );
na02f80 g777096 ( .a(n_3832), .b(n_3794), .o(n_4035) );
na02f80 FE_RC_1992_0 ( .a(n_20002), .b(FE_RN_650_0), .o(n_20062) );
in01f80 newInst_2171 ( .a(newNet_2170), .o(newNet_2171) );
na02f80 g767060 ( .a(n_14758), .b(n_14256), .o(n_14385) );
in01f80 g770170 ( .a(n_10803), .o(n_10804) );
na02f80 g744049 ( .a(n_44221), .b(n_34677), .o(n_35747) );
oa22f80 g743777 ( .a(n_36322), .b(n_36289), .c(n_36323), .d(n_36290), .o(n_36389) );
in01f80 newInst_3155 ( .a(newNet_1977), .o(newNet_3155) );
ao12f80 g746630 ( .a(n_34333), .b(n_34359), .c(n_34332), .o(n_34889) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_14_ ( .ck(newNet_3333), .d(n_31958), .o(delay_add_ln22_unr20_stage8_stallmux_q_14_) );
na02f80 g773124 ( .a(n_7654), .b(n_45825), .o(n_7703) );
oa12f80 g763759 ( .a(n_17202), .b(n_17096), .c(n_17427), .o(n_17372) );
in01f80 newInst_2358 ( .a(newNet_2168), .o(newNet_2358) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_12_ ( .ck(newNet_1033), .d(n_17777), .o(delay_xor_ln21_unr12_stage5_stallmux_q_12_) );
no02f80 g764244 ( .a(n_16296), .b(n_16336), .o(n_16443) );
no02f80 g759124 ( .a(n_21346), .b(n_45024), .o(n_21388) );
in01f80 g767718 ( .a(n_12745), .o(n_12746) );
oa12f80 g736308 ( .a(n_305), .b(n_43866), .c(FE_OFN2_n_43918), .o(n_43905) );
na02f80 g742087 ( .a(FE_OCP_RBN3445_n_37945), .b(n_38235), .o(n_38316) );
na02f80 g763407 ( .a(n_16975), .b(n_16038), .o(n_17215) );
na02f80 g776019 ( .a(n_5061), .b(n_5018), .o(n_5098) );
no03m80 FE_RC_463_0 ( .a(FE_RN_134_0), .b(n_23131), .c(n_23460), .o(n_23504) );
oa22f80 FE_RC_4117_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .b(FE_OCP_RBN3282_n_44365), .c(n_44365), .d(FE_OCP_RBN3801_delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(n_16801) );
no02f80 g754011 ( .a(n_26129), .b(n_26128), .o(n_26130) );
oa22f80 g756836 ( .a(n_23420), .b(n_23304), .c(n_23386), .d(n_23303), .o(n_24838) );
na02f80 FE_RC_3847_0 ( .a(n_23369), .b(FE_RN_1678_0), .o(n_23615) );
no02f80 g760482 ( .a(n_20021), .b(FE_OCP_RBN1156_n_18375), .o(n_20092) );
no02f80 g748655 ( .a(n_31269), .b(n_31268), .o(n_31270) );
no02f80 g756643 ( .a(n_23555), .b(n_23554), .o(n_23577) );
no02f80 g765080 ( .a(n_15238), .b(n_15239), .o(n_15349) );
no02f80 g760828 ( .a(n_19585), .b(FE_OCPN1790_n_18119), .o(n_19685) );
na02f80 g748820 ( .a(n_32497), .b(n_32447), .o(n_32656) );
na02f80 g768567 ( .a(n_12161), .b(n_12236), .o(n_12336) );
in01f80 g755783 ( .a(n_24398), .o(n_24399) );
oa22f80 g753360 ( .a(n_26882), .b(n_26776), .c(n_26852), .d(n_26777), .o(n_26969) );
na02f80 g745748 ( .a(n_34184), .b(n_34160), .o(n_34185) );
oa12f80 g767406 ( .a(n_13546), .b(n_13545), .c(n_13544), .o(n_14038) );
no02f80 g758222 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_), .o(n_22839) );
no02f80 g761393 ( .a(n_18922), .b(n_18946), .o(n_19025) );
no02f80 FE_RC_2810_0 ( .a(n_9578), .b(n_9672), .o(FE_RN_1202_0) );
in01f80 g780431 ( .a(n_921), .o(n_920) );
na02f80 g746244 ( .a(FE_OCP_RBN1354_n_33584), .b(n_33594), .o(n_33662) );
na02f80 g767457 ( .a(n_13230), .b(n_13231), .o(n_13367) );
in01f80 g736343 ( .a(n_43829), .o(n_43830) );
ao12f80 g766617 ( .a(n_14309), .b(n_14308), .c(n_14307), .o(n_16138) );
na02f80 g744125 ( .a(n_36184), .b(n_36243), .o(n_36262) );
na02f80 g745864 ( .a(n_44102), .b(n_33614), .o(n_34219) );
in01f80 g743112 ( .a(n_37108), .o(n_37045) );
in01f80 g761633 ( .a(n_18893), .o(n_18892) );
no02f80 g777966 ( .a(n_3069), .b(n_3068), .o(n_3070) );
oa12f80 g743394 ( .a(n_37788), .b(n_37787), .c(n_46248), .o(n_37826) );
no02f80 g779588 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .o(n_1861) );
na02f80 g739356 ( .a(n_45153), .b(n_40514), .o(n_40829) );
no02f80 g738913 ( .a(n_41215), .b(n_41048), .o(n_41252) );
na02f80 g743991 ( .a(n_36264), .b(n_35697), .o(n_36332) );
in01f80 newInst_2008 ( .a(newNet_2007), .o(newNet_2008) );
no02f80 g738167 ( .a(n_42006), .b(n_41912), .o(n_42025) );
na02f80 g736606 ( .a(n_43623), .b(n_43625), .o(n_43637) );
na02f80 g773881 ( .a(n_7086), .b(n_7085), .o(n_7333) );
ao12f80 g774388 ( .a(n_6836), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .o(n_7313) );
in01f80 g743512 ( .a(n_37711), .o(n_37712) );
in01f80 FE_OCP_RBC2438_n_8402 ( .a(FE_OCP_RBN2437_n_8402), .o(FE_OCP_RBN2438_n_8402) );
in01f80 g743531 ( .a(n_36520), .o(n_36505) );
na02f80 g736695 ( .a(n_43433), .b(n_43363), .o(n_43434) );
in01f80 g770618 ( .a(n_10454), .o(n_10455) );
na02f80 g772252 ( .a(n_8753), .b(n_8752), .o(n_8770) );
na02f80 g757660 ( .a(n_22582), .b(n_22634), .o(n_22672) );
na02f80 g766563 ( .a(n_13867), .b(n_12930), .o(n_13955) );
na02f80 g778716 ( .a(FE_OCP_RBN2294_n_2438), .b(n_2472), .o(n_2491) );
in01f80 g780882 ( .a(n_497), .o(n_508) );
in01f80 fopt783089 ( .a(n_44568), .o(n_44566) );
no02f80 g742264 ( .a(n_37824), .b(n_37812), .o(n_37861) );
na02f80 g741987 ( .a(n_37895), .b(n_37906), .o(n_37954) );
na02f80 g747614 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_32347) );
no02f80 g742253 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37352), .o(n_38310) );
no02f80 g760412 ( .a(n_20080), .b(n_20100), .o(n_20164) );
in01f80 g774561 ( .a(FE_OCPN895_n_6521), .o(n_6624) );
in01f80 g754286 ( .a(n_25915), .o(n_27170) );
in01f80 FE_OCPC1392_n_7925 ( .a(FE_OCPN1391_n_7925), .o(FE_OCPN1392_n_7925) );
ao12f80 g774379 ( .a(n_6749), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .o(n_6920) );
na02f80 g772912 ( .a(n_7845), .b(n_7847), .o(n_8066) );
no02f80 g766934 ( .a(n_13972), .b(n_14109), .o(n_14620) );
na02f80 FE_RC_3480_0 ( .a(n_40074), .b(n_40037), .o(FE_RN_1496_0) );
in01f80 newInst_2537 ( .a(newNet_2536), .o(newNet_2537) );
in01f80 g759853 ( .a(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_22207) );
na02f80 g772573 ( .a(n_8221), .b(FE_OCP_RBN2301_n_7817), .o(n_8248) );
in01f80 g737504 ( .a(n_43083), .o(n_42596) );
in01f80 FE_RC_4027_0 ( .a(n_14452), .o(FE_RN_1749_0) );
na02f80 g777163 ( .a(n_5368), .b(n_5298), .o(n_5385) );
na02f80 g764384 ( .a(n_16416), .b(n_16386), .o(n_16451) );
na02f80 g746891 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_18_), .o(n_33107) );
no02f80 g744937 ( .a(n_34905), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34935) );
in01f80 g737713 ( .a(n_42445), .o(n_42418) );
ao12f80 g737517 ( .a(n_42533), .b(n_42532), .c(n_42531), .o(n_43121) );
in01f80 newInst_832 ( .a(newNet_831), .o(newNet_832) );
in01f80 g746933 ( .a(n_32914), .o(n_32944) );
na02f80 FE_RC_309_0 ( .a(FE_RN_92_0), .b(n_21576), .o(n_46966) );
ao12f80 g756439 ( .a(n_23572), .b(n_23876), .c(n_22936), .o(n_24011) );
in01f80 g750773 ( .a(n_29364), .o(n_29365) );
no02f80 g766308 ( .a(n_14194), .b(n_13257), .o(n_14242) );
in01f80 newInst_184 ( .a(newNet_121), .o(newNet_184) );
na02f80 g766215 ( .a(n_14468), .b(n_13469), .o(n_14471) );
in01f80 FE_OCP_RBC3110_n_43711 ( .a(n_43711), .o(FE_OCP_RBN3110_n_43711) );
ao12f80 g770113 ( .a(n_10360), .b(FE_OCP_RBN2899_n_44853), .c(n_10699), .o(n_10731) );
in01f80 g749178 ( .a(n_32203), .o(n_32204) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_0_ ( .ck(newNet_3266), .d(n_35309), .o(delay_add_ln22_unr23_stage9_stallmux_q_0_) );
in01f80 newInst_3661 ( .a(newNet_3605), .o(newNet_3661) );
na02f80 g771625 ( .a(n_9237), .b(n_9036), .o(n_9276) );
ao12f80 g768474 ( .a(n_12298), .b(n_12302), .c(n_11707), .o(n_12418) );
in01f80 g749493 ( .a(n_30467), .o(n_30468) );
ao12f80 g745783 ( .a(n_34111), .b(n_34094), .c(n_34076), .o(n_34191) );
na02f80 g744698 ( .a(n_36513), .b(n_36026), .o(n_36574) );
na02f80 g766204 ( .a(n_14447), .b(FE_OCP_RBN2481_n_14270), .o(n_14448) );
in01f80 g746361 ( .a(n_33539), .o(n_33540) );
ao22s80 g736687 ( .a(n_43065), .b(n_43072), .c(n_43064), .d(n_43050), .o(n_43151) );
in01f80 FE_OCP_DRV_C1536_n_12633 ( .a(FE_OCP_DRV_N1535_n_12633), .o(FE_OCP_DRV_N1536_n_12633) );
in01f80 g770776 ( .a(n_10030), .o(n_10068) );
no02f80 g764607 ( .a(n_16035), .b(n_16072), .o(n_16216) );
in01f80 newInst_1588 ( .a(newNet_752), .o(newNet_1588) );
no02f80 g748886 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n_32414) );
na02f80 g781094 ( .a(n_258), .b(n_249), .o(n_250) );
no02f80 g776922 ( .a(n_3995), .b(n_4046), .o(n_4176) );
na02f80 g772958 ( .a(n_7814), .b(n_8568), .o(n_7846) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_27_ ( .ck(newNet_2372), .d(FE_OFN615_n_36594), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_) );
no02f80 g773563 ( .a(n_7450), .b(n_7449), .o(n_7451) );
no02f80 g773501 ( .a(n_7489), .b(n_7294), .o(n_7526) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_17_ ( .ck(newNet_3633), .d(n_16916), .o(delay_add_ln22_unr11_stage5_stallmux_q_17_) );
in01f80 g780230 ( .a(n_1138), .o(n_1152) );
na02f80 g770269 ( .a(n_10752), .b(n_10751), .o(n_10753) );
in01f80 g755508 ( .a(FE_OCPN1048_n_24819), .o(n_24865) );
in01f80 g780523 ( .a(n_825), .o(n_826) );
no02f80 g749148 ( .a(n_30858), .b(n_30809), .o(n_30875) );
in01f80 g743541 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .o(n_36991) );
in01f80 newInst_2541 ( .a(newNet_2540), .o(newNet_2541) );
in01f80 g754251 ( .a(FE_OCP_RBN2815_n_25986), .o(n_26011) );
in01f80 g779699 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n_1373) );
ao12f80 g773781 ( .a(n_7120), .b(n_7137), .c(n_7119), .o(n_7212) );
in01f80 g773053 ( .a(n_8021), .o(n_8069) );
na02f80 g736824 ( .a(n_43128), .b(n_42856), .o(n_43141) );
oa12f80 g745646 ( .a(n_34102), .b(n_34101), .c(n_34121), .o(n_34151) );
no02f80 g764965 ( .a(n_15498), .b(n_15496), .o(n_15612) );
na02f80 g751884 ( .a(n_29001), .b(n_29285), .o(n_29073) );
no02f80 g738874 ( .a(n_41261), .b(n_41260), .o(n_41262) );
in01f80 FE_RC_1533_0 ( .a(n_28095), .o(FE_RN_433_0) );
in01f80 g780364 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .o(n_1392) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_12_ ( .ck(newNet_1344), .d(n_1166), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_) );
oa12f80 g775022 ( .a(n_6188), .b(n_6128), .c(n_6106), .o(n_6201) );
oa12f80 g779262 ( .a(n_1763), .b(n_1762), .c(n_1789), .o(n_2466) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_18_ ( .ck(newNet_731), .d(n_46178), .o(delay_xor_ln21_unr6_stage3_stallmux_q_18_) );
no02f80 FE_RC_2307_0 ( .a(FE_RN_869_0), .b(FE_RN_874_0), .o(n_25904) );
in01f80 g762356 ( .a(n_18578), .o(n_18533) );
in01f80 g753973 ( .a(n_27035), .o(n_27051) );
ao12f80 g745871 ( .a(n_34016), .b(n_34015), .c(n_34017), .o(n_35482) );
no02f80 g762401 ( .a(n_18421), .b(n_18418), .o(n_18444) );
na02f80 g745284 ( .a(n_34514), .b(n_34459), .o(n_34513) );
na02f80 g769239 ( .a(n_11480), .b(n_11399), .o(n_11550) );
na02f80 g774297 ( .a(FE_OCP_RBN3252_delay_xor_ln22_unr6_stage3_stallmux_q_0_), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6642) );
na02f80 g773446 ( .a(n_7561), .b(n_7147), .o(n_7659) );
in01f80 newInst_816 ( .a(newNet_643), .o(newNet_816) );
in01f80 newInst_582 ( .a(newNet_581), .o(newNet_582) );
na02f80 g769861 ( .a(n_11154), .b(n_10239), .o(n_11176) );
no02f80 FE_RC_4102_0 ( .a(FE_RN_1795_0), .b(n_32000), .o(n_32088) );
in01f80 g765685 ( .a(n_15874), .o(n_16245) );
in01f80 g755157 ( .a(n_25100), .o(n_25101) );
in01f80 newInst_2841 ( .a(newNet_2840), .o(newNet_2841) );
na02f80 g773496 ( .a(n_7446), .b(n_6413), .o(n_7501) );
in01f80 FE_OCPC884_n_42216 ( .a(n_42216), .o(FE_OCPN884_n_42216) );
na02f80 g739207 ( .a(n_40890), .b(n_40889), .o(n_41229) );
in01f80 g738938 ( .a(n_41631), .o(n_41275) );
in01f80 newInst_2893 ( .a(newNet_2892), .o(newNet_2893) );
in01f80 FE_OCP_RBC2167_n_32892 ( .a(n_32892), .o(FE_OCP_RBN2167_n_32892) );
na02f80 g761019 ( .a(n_20039), .b(n_19985), .o(n_20055) );
in01f80 newInst_2716 ( .a(newNet_2527), .o(newNet_2716) );
oa22f80 FE_RC_746_0 ( .a(FE_OCP_RBN2393_n_8288), .b(FE_OCP_RBN3455_FE_OCPN1240_n_7721), .c(FE_OCPN890_n_7802), .d(n_8288), .o(n_8410) );
oa22f80 FE_RC_1178_0 ( .a(n_22966), .b(n_22945), .c(n_22965), .d(n_22900), .o(n_23069) );
no02f80 g741806 ( .a(n_38397), .b(n_38396), .o(n_38398) );
in01f80 newInst_1642 ( .a(newNet_1641), .o(newNet_1642) );
no02f80 g741339 ( .a(n_44944), .b(n_38470), .o(n_38928) );
in01f80 FE_OCP_RBC2324_n_13616 ( .a(n_13616), .o(FE_OCP_RBN2324_n_13616) );
oa22f80 g754605 ( .a(FE_OCP_RBN2957_n_26231), .b(n_26512), .c(FE_OCP_RBN2960_n_26231), .d(n_25745), .o(n_26884) );
no02f80 g753939 ( .a(n_26196), .b(FE_OCPN1748_n_23354), .o(n_26359) );
na02f80 g757002 ( .a(n_23619), .b(n_23618), .o(n_23620) );
na02f80 g754735 ( .a(n_25461), .b(n_25460), .o(n_25462) );
in01f80 g738517 ( .a(n_41667), .o(n_41730) );
in01f80 g773722 ( .a(n_7801), .o(n_7296) );
in01f80 newInst_309 ( .a(newNet_308), .o(newNet_309) );
in01f80 FE_RC_3796_0 ( .a(n_19615), .o(FE_RN_1658_0) );
no02f80 g764356 ( .a(n_16418), .b(n_16318), .o(n_16419) );
in01f80 g744142 ( .a(n_35859), .o(n_35860) );
no02f80 g740346 ( .a(n_40247), .b(n_40168), .o(n_40271) );
in01f80 g775669 ( .a(n_5598), .o(n_5599) );
in01f80 FE_OCP_DRV_C1596_n_21458 ( .a(FE_OCP_DRV_N1595_n_21458), .o(FE_OCP_DRV_N1596_n_21458) );
in01f80 newInst_228 ( .a(newNet_227), .o(newNet_228) );
in01f80 g736897 ( .a(n_43583), .o(n_43584) );
na02f80 g777268 ( .a(n_3546), .b(n_2913), .o(n_3653) );
in01f80 newInst_3360 ( .a(newNet_3359), .o(newNet_3360) );
na02f80 g771755 ( .a(n_10158), .b(n_10121), .o(n_10248) );
no02f80 g772653 ( .a(n_8318), .b(n_7886), .o(n_8320) );
in01f80 g743121 ( .a(n_37042), .o(n_37146) );
in01f80 g765308 ( .a(n_16017), .o(n_16098) );
na02f80 g753511 ( .a(n_26778), .b(n_26422), .o(n_26805) );
no02f80 g741667 ( .a(n_38552), .b(n_38567), .o(n_38596) );
no02f80 g753981 ( .a(n_26249), .b(n_26248), .o(n_26362) );
in01f80 FE_OCP_RBC3852_n_20848 ( .a(n_20848), .o(FE_OCP_RBN3852_n_20848) );
no02f80 g772249 ( .a(n_8753), .b(n_8752), .o(n_8794) );
in01f80 g762669 ( .a(FE_OCP_DRV_N1556_n_19384), .o(n_19508) );
in01f80 FE_RC_3394_0 ( .a(n_16466), .o(FE_RN_1469_0) );
in01f80 g779596 ( .a(n_2011), .o(n_2012) );
na02f80 g773219 ( .a(n_7802), .b(n_7982), .o(n_7960) );
na02f80 g744031 ( .a(n_44223), .b(FE_OCP_DRV_N1598_n_35644), .o(n_36304) );
in01f80 g765927 ( .a(n_14818), .o(n_14819) );
na02f80 g740504 ( .a(n_39683), .b(n_39690), .o(n_39701) );
in01f80 FE_OCP_RBC2428_n_8300 ( .a(n_8300), .o(FE_OCP_RBN2428_n_8300) );
no02f80 g772352 ( .a(n_8606), .b(n_8605), .o(n_8607) );
na02f80 g743343 ( .a(n_36730), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36786) );
no02f80 g737750 ( .a(n_42200), .b(n_42207), .o(n_42240) );
ao12f80 g780334 ( .a(n_861), .b(n_937), .c(n_860), .o(n_962) );
in01f80 FE_OCP_RBC3090_FE_OCPN1052_n_31674 ( .a(FE_OCPN1052_n_31674), .o(FE_OCP_RBN3090_FE_OCPN1052_n_31674) );
in01f80 g768678 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_), .o(n_12188) );
no02f80 g767768 ( .a(n_13317), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .o(n_13369) );
in01f80 g754563 ( .a(n_26681), .o(n_26682) );
in01f80 newInst_3668 ( .a(newNet_3667), .o(newNet_3668) );
no02f80 g778591 ( .a(n_2534), .b(n_2533), .o(n_2844) );
in01f80 g776663 ( .a(n_4218), .o(n_4243) );
no02f80 g764635 ( .a(n_16449), .b(n_15883), .o(n_16547) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_31_ ( .ck(newNet_1806), .d(n_16888), .o(n_17093) );
na02f80 g746753 ( .a(n_32977), .b(n_33021), .o(n_33037) );
na02f80 g758229 ( .a(FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .o(n_22699) );
no02f80 g754555 ( .a(n_26486), .b(n_26512), .o(n_26513) );
in01f80 newInst_1240 ( .a(newNet_1239), .o(newNet_1240) );
in01f80 g779712 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .o(n_1368) );
oa12f80 g745436 ( .a(n_34274), .b(n_34298), .c(n_34273), .o(n_35469) );
na02f80 g768066 ( .a(n_12709), .b(n_12699), .o(n_12718) );
na02f80 g749825 ( .a(n_30976), .b(n_30975), .o(n_30977) );
in01f80 g774242 ( .a(n_6652), .o(n_6653) );
in01f80 g778962 ( .a(n_2160), .o(n_2189) );
in01f80 g777659 ( .a(n_3539), .o(n_3540) );
ao12f80 g754876 ( .a(n_25046), .b(n_25187), .c(n_25105), .o(n_25282) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_24_ ( .ck(newNet_3304), .d(FE_OCP_RBN3122_n_32239), .o(delay_add_ln22_unr20_stage8_stallmux_q_24_) );
no02f80 g750925 ( .a(n_30105), .b(n_30288), .o(n_30305) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_8_ ( .ck(newNet_689), .d(n_46171), .o(delay_xor_ln21_unr6_stage3_stallmux_q_8_) );
in01f80 FE_OCP_RBC2186_n_37686 ( .a(n_37686), .o(FE_OCP_RBN2186_n_37686) );
na02f80 g780884 ( .a(n_377), .b(n_398), .o(n_426) );
in01f80 g758240 ( .a(n_22783), .o(n_22760) );
in01f80 g736936 ( .a(n_43213), .o(n_43272) );
na02f80 g771403 ( .a(n_9166), .b(n_8927), .o(n_9215) );
in01f80 g754525 ( .a(n_26714), .o(n_26686) );
in01f80 g774123 ( .a(n_6719), .o(n_6701) );
in01f80 newInst_378 ( .a(newNet_377), .o(newNet_378) );
oa22f80 g777021 ( .a(n_5447), .b(n_3700), .c(n_3620), .d(n_3788), .o(n_3995) );
no02f80 g738273 ( .a(n_41777), .b(n_41595), .o(n_41873) );
in01f80 newInst_2534 ( .a(newNet_2533), .o(newNet_2534) );
no02f80 g755068 ( .a(n_25353), .b(n_25291), .o(n_25378) );
oa12f80 g764887 ( .a(n_16136), .b(n_16026), .c(n_16135), .o(n_16356) );
no02f80 g754017 ( .a(n_26121), .b(n_26037), .o(n_26155) );
na02f80 g736596 ( .a(n_43334), .b(n_43084), .o(n_43417) );
no02f80 g771623 ( .a(n_9328), .b(n_9286), .o(n_9368) );
in01f80 g767384 ( .a(n_13336), .o(n_13343) );
na02f80 g744264 ( .a(FE_OCPN1510_n_44174), .b(n_35569), .o(n_36188) );
in01f80 g739423 ( .a(n_40806), .o(n_40807) );
in01f80 g757757 ( .a(n_22739), .o(n_22789) );
in01f80 newInst_1284 ( .a(newNet_1200), .o(newNet_1284) );
na02f80 g779123 ( .a(n_1979), .b(FE_RN_518_0), .o(n_2239) );
in01f80 g745203 ( .a(n_34440), .o(n_34601) );
in01f80 FE_OCPC1522_n_26054 ( .a(FE_OCPN1521_n_26054), .o(FE_OCPN1522_n_26054) );
oa22f80 g753658 ( .a(n_27198), .b(n_26681), .c(n_27199), .d(n_26682), .o(n_27318) );
in01f80 FE_RC_465_0 ( .a(n_28381), .o(FE_RN_135_0) );
na02f80 g750463 ( .a(n_29546), .b(FE_OFN788_n_25834), .o(n_29549) );
in01f80 newInst_3402 ( .a(newNet_1628), .o(newNet_3402) );
no02f80 g771096 ( .a(n_9554), .b(FE_OCP_RBN2588_n_9492), .o(n_9638) );
in01f80 FE_OCP_RBC3519_n_8498 ( .a(FE_OCP_RBN3517_n_8498), .o(FE_OCP_RBN3519_n_8498) );
no02f80 g748717 ( .a(n_31163), .b(n_31162), .o(n_31204) );
no02f80 g755094 ( .a(n_25099), .b(n_23793), .o(n_25147) );
in01f80 g756798 ( .a(n_23411), .o(n_23396) );
in01f80 g758988 ( .a(n_21326), .o(n_21327) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_20_ ( .ck(newNet_1617), .d(n_27318), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_) );
in01f80 FE_RC_375_0 ( .a(n_12456), .o(FE_RN_111_0) );
oa12f80 g763775 ( .a(n_17101), .b(n_17304), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .o(n_17365) );
no02f80 g759381 ( .a(n_20801), .b(n_20776), .o(n_20889) );
oa22f80 g758020 ( .a(n_22015), .b(n_21962), .c(n_22014), .d(n_21963), .o(n_22107) );
no02f80 g738382 ( .a(n_41664), .b(n_41665), .o(n_41941) );
in01f80 FE_RC_3577_0 ( .a(n_14169), .o(FE_RN_1556_0) );
in01f80 newInst_2244 ( .a(newNet_696), .o(newNet_2244) );
in01f80 newInst_1275 ( .a(newNet_1274), .o(newNet_1275) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_25_ ( .ck(newNet_1216), .d(n_6183), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_) );
na02f80 g746555 ( .a(n_34550), .b(n_34585), .o(n_34551) );
in01f80 g740735 ( .a(n_39553), .o(n_40007) );
na02f80 g780868 ( .a(n_354), .b(beta_3), .o(n_367) );
in01f80 g740510 ( .a(n_39758), .o(n_39759) );
ao12f80 g738610 ( .a(n_41486), .b(n_41716), .c(n_41062), .o(n_41835) );
in01f80 g746917 ( .a(n_33149), .o(n_33150) );
in01f80 newInst_1866 ( .a(newNet_1605), .o(newNet_1866) );
no02f80 g766955 ( .a(n_13897), .b(n_14039), .o(n_14392) );
no02f80 g766863 ( .a(n_13574), .b(n_13595), .o(n_13693) );
oa12f80 g737262 ( .a(n_42295), .b(n_42918), .c(n_42344), .o(n_42927) );
ao12f80 g759793 ( .a(n_21142), .b(n_21141), .c(n_21140), .o(n_21798) );
no02f80 g747956 ( .a(n_33119), .b(n_33118), .o(n_33120) );
no02f80 g773577 ( .a(n_7372), .b(delay_add_ln22_unr5_stage3_stallmux_q_20_), .o(n_7384) );
no02f80 g780082 ( .a(n_1192), .b(n_790), .o(n_1213) );
no02f80 g741880 ( .a(n_38205), .b(n_38040), .o(n_38206) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_11_ ( .ck(newNet_983), .d(n_22893), .o(delay_xor_ln21_unr15_stage6_stallmux_q_11_) );
na02f80 g763419 ( .a(n_16976), .b(n_17032), .o(n_17132) );
na02f80 g744211 ( .a(n_36090), .b(n_35780), .o(n_36238) );
no02f80 g780421 ( .a(n_821), .b(FE_OFN759_n_45813), .o(n_860) );
in01f80 g777189 ( .a(n_5342), .o(n_5343) );
in01f80 FE_RC_4150_0 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(FE_RN_1805_0) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_26_ ( .ck(newNet_2171), .d(n_981), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_) );
oa12f80 g757826 ( .a(n_22982), .b(n_22983), .c(n_22981), .o(n_23698) );
na02f80 g776915 ( .a(n_3948), .b(n_3920), .o(n_3949) );
in01f80 g740208 ( .a(n_39975), .o(n_39998) );
oa22f80 FE_RC_3893_0 ( .a(n_19170), .b(n_19241), .c(n_18010), .d(FE_OCP_RBN3833_n_19241), .o(n_19377) );
na02f80 g776306 ( .a(n_4473), .b(n_3297), .o(n_4665) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_3_ ( .ck(newNet_624), .d(n_46379), .o(delay_xor_ln21_unr9_stage4_stallmux_q_3_) );
no02f80 g779121 ( .a(n_1999), .b(n_1759), .o(n_2024) );
na02f80 g767686 ( .a(n_13193), .b(n_13121), .o(n_13257) );
ao12f80 g767713 ( .a(n_13319), .b(n_13084), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n_13363) );
in01f80 newInst_2977 ( .a(newNet_2976), .o(newNet_2977) );
in01f80 newInst_2547 ( .a(newNet_375), .o(newNet_2547) );
oa22f80 FE_RC_1149_0 ( .a(n_1476), .b(n_1716), .c(n_1477), .d(n_1672), .o(n_1753) );
na02f80 g750181 ( .a(n_29753), .b(n_28656), .o(n_29814) );
no02f80 g753446 ( .a(n_26987), .b(n_26537), .o(n_27006) );
in01f80 FE_OCPC1531_n_21790 ( .a(n_21790), .o(FE_OCPN1531_n_21790) );
na02f80 g759719 ( .a(n_21671), .b(n_21670), .o(n_21672) );
na02f80 g776119 ( .a(n_4855), .b(n_4742), .o(n_4920) );
no02f80 g752606 ( .a(n_27573), .b(n_27300), .o(n_27598) );
in01f80 g767308 ( .a(n_13538), .o(n_13608) );
no02f80 g761370 ( .a(n_19024), .b(n_19022), .o(n_19186) );
in01f80 g780246 ( .a(n_1089), .o(n_1067) );
in01f80 g740266 ( .a(n_40171), .o(n_40172) );
oa12f80 g779242 ( .a(n_1769), .b(n_1795), .c(n_1768), .o(n_1835) );
in01f80 g761741 ( .a(n_18852), .o(n_18853) );
no02f80 g773069 ( .a(n_7920), .b(n_7996), .o(n_8014) );
na02f80 g781073 ( .a(sin_out_1), .b(FE_OFN5_n_43918), .o(n_299) );
in01f80 g767254 ( .a(n_13562), .o(n_13563) );
no02f80 g754574 ( .a(FE_OCP_RBN2959_n_26231), .b(n_26734), .o(n_26769) );
in01f80 g747600 ( .a(n_32427), .o(n_32512) );
na02f80 g737771 ( .a(n_42496), .b(n_42403), .o(n_42531) );
na02f80 g772938 ( .a(n_7884), .b(n_7883), .o(n_7931) );
in01f80 FE_OCP_RBC1147_n_13098 ( .a(FE_OCP_RBN1145_n_13098), .o(FE_OCP_RBN1147_n_13098) );
no02f80 g758899 ( .a(n_21433), .b(n_21432), .o(n_21546) );
no02f80 g779156 ( .a(n_1921), .b(n_1919), .o(n_1920) );
ao22s80 g778972 ( .a(FE_OCP_RBN3434_n_2224), .b(n_1996), .c(n_2224), .d(n_1997), .o(n_2284) );
ms00f80 sin_out_reg_3_ ( .ck(newNet_26), .d(n_43680), .o(sin_out_3) );
na02f80 g770752 ( .a(n_9971), .b(n_9963), .o(n_10058) );
in01f80 newInst_3157 ( .a(newNet_3156), .o(newNet_3157) );
in01f80 g742558 ( .a(n_37638), .o(n_37639) );
in01f80 g753745 ( .a(n_27132), .o(n_27133) );
na02f80 g736902 ( .a(n_43189), .b(n_43482), .o(n_43579) );
in01f80 g758219 ( .a(n_23006), .o(n_23051) );
oa12f80 g739761 ( .a(n_40368), .b(n_40468), .c(n_40132), .o(n_40526) );
in01f80 g770945 ( .a(n_9893), .o(n_9894) );
na02f80 g737780 ( .a(n_42327), .b(n_42304), .o(n_42305) );
na02f80 g771292 ( .a(n_9513), .b(n_8185), .o(n_9659) );
in01f80 FE_RC_1102_0 ( .a(n_40756), .o(FE_RN_328_0) );
in01f80 newInst_926 ( .a(newNet_925), .o(newNet_926) );
na02f80 g765486 ( .a(n_14985), .b(n_14210), .o(n_15022) );
ao12f80 g747986 ( .a(n_31560), .b(n_31813), .c(n_31613), .o(n_31883) );
na02f80 g772566 ( .a(n_8248), .b(n_8277), .o(n_8385) );
in01f80 FE_OCP_RBC2282_n_29111 ( .a(n_29111), .o(FE_OCP_RBN2282_n_29111) );
na02f80 g755084 ( .a(n_25582), .b(n_25612), .o(n_25691) );
oa12f80 g772712 ( .a(n_8181), .b(n_8180), .c(n_8197), .o(n_8239) );
no02f80 g751990 ( .a(n_28793), .b(n_28810), .o(n_29200) );
in01f80 newInst_1376 ( .a(newNet_1375), .o(newNet_1376) );
no02f80 g750739 ( .a(n_44139), .b(n_29160), .o(n_29342) );
na02f80 g743125 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .o(n_37161) );
na02f80 g761319 ( .a(n_19710), .b(n_19731), .o(n_19732) );
na02f80 g777703 ( .a(n_3354), .b(n_3353), .o(n_3355) );
na02f80 g759013 ( .a(n_22009), .b(n_22008), .o(n_22010) );
na02f80 g753602 ( .a(n_26669), .b(n_26563), .o(n_26694) );
ao12f80 g737622 ( .a(n_42370), .b(n_42305), .c(n_42202), .o(n_42371) );
in01f80 FE_OCP_RBC2805_n_30534 ( .a(n_30534), .o(FE_OCP_RBN2805_n_30534) );
na02f80 g755578 ( .a(n_24505), .b(n_24620), .o(n_24537) );
oa22f80 g739828 ( .a(n_40414), .b(n_40360), .c(n_40415), .d(n_40359), .o(n_40459) );
in01f80 g746710 ( .a(n_33290), .o(n_33328) );
in01f80 g751214 ( .a(n_28852), .o(n_28807) );
in01f80 g747945 ( .a(n_33683), .o(n_33170) );
no02f80 g784778 ( .a(n_35861), .b(n_44223), .o(n_47264) );
ao12f80 g763707 ( .a(n_46426), .b(n_16643), .c(n_47268), .o(n_16712) );
na03f80 g756526 ( .a(n_23808), .b(n_24077), .c(n_24110), .o(n_24238) );
in01f80 g748633 ( .a(n_31332), .o(n_31333) );
in01f80 FE_OCP_RBC3448_n_37945 ( .a(FE_OCP_RBN3445_n_37945), .o(FE_OCP_RBN3448_n_37945) );
in01f80 newInst_1243 ( .a(newNet_1238), .o(newNet_1243) );
na02f80 g745466 ( .a(n_34561), .b(n_34369), .o(n_34653) );
no02f80 g757501 ( .a(n_22827), .b(delay_add_ln22_unr14_stage6_stallmux_q_1_), .o(n_22940) );
ao12f80 g737636 ( .a(n_42396), .b(n_42392), .c(n_42423), .o(n_42762) );
na02f80 g763245 ( .a(n_17736), .b(n_17711), .o(n_17712) );
in01f80 FE_OCPC1514_FE_OFN738_n_22641 ( .a(FE_OCPN1513_FE_OFN738_n_22641), .o(FE_OCPN1514_FE_OFN738_n_22641) );
in01f80 g758580 ( .a(n_22094), .o(n_22095) );
in01f80 newInst_3677 ( .a(newNet_3676), .o(newNet_3677) );
in01f80 g769600 ( .a(n_11392), .o(n_11372) );
in01f80 newInst_19 ( .a(newNet_18), .o(newNet_19) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_15_ ( .ck(newNet_3332), .d(n_31999), .o(delay_add_ln22_unr20_stage8_stallmux_q_15_) );
na02f80 g767843 ( .a(n_12852), .b(n_11663), .o(n_13015) );
na02f80 g745413 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35602), .o(n_35604) );
in01f80 newInst_2914 ( .a(newNet_2667), .o(newNet_2914) );
no02f80 g757210 ( .a(n_44068), .b(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .o(n_23114) );
in01f80 newInst_488 ( .a(newNet_487), .o(newNet_488) );
in01f80 g753024 ( .a(n_27923), .o(n_27899) );
in01f80 g773497 ( .a(n_7490), .o(n_7491) );
oa12f80 g751394 ( .a(FE_OCPN1038_n_28318), .b(n_28478), .c(FE_OCPN1036_n_28288), .o(n_28536) );
na02f80 g750089 ( .a(n_29841), .b(n_29866), .o(n_29894) );
in01f80 g747651 ( .a(n_32394), .o(n_32463) );
na02f80 g776405 ( .a(n_4641), .b(n_4677), .o(n_4809) );
na02f80 g738472 ( .a(n_41393), .b(n_41392), .o(n_41414) );
no02f80 g748107 ( .a(n_32807), .b(n_32806), .o(n_32808) );
in01f80 FE_OFC810_n_1941 ( .a(FE_OFN827_n_1941), .o(FE_OFN810_n_1941) );
in01f80 g781235 ( .a(n_131), .o(n_132) );
in01f80 g769789 ( .a(n_11236), .o(n_11237) );
no02f80 g767437 ( .a(n_13505), .b(n_13504), .o(n_13506) );
in01f80 FE_OCP_RBC2599_n_34388 ( .a(FE_OCP_RBN2598_n_34388), .o(FE_OCP_RBN2599_n_34388) );
na02f80 g772328 ( .a(n_8660), .b(n_8682), .o(n_8719) );
ao12f80 g780852 ( .a(n_369), .b(n_354), .c(n_368), .o(n_370) );
in01f80 g772467 ( .a(n_8460), .o(n_8466) );
no03m80 FE_RC_1125_0 ( .a(FE_RN_341_0), .b(n_23390), .c(n_23211), .o(n_23313) );
oa12f80 g773748 ( .a(n_7231), .b(n_7230), .c(n_7229), .o(n_7700) );
in01f80 g759036 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_), .o(n_23135) );
in01f80 newInst_2886 ( .a(newNet_2885), .o(newNet_2886) );
na02f80 g768967 ( .a(n_11852), .b(n_11798), .o(n_11825) );
oa12f80 g742890 ( .a(n_46256), .b(n_37126), .c(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n_37127) );
ao22s80 g754606 ( .a(FE_OCP_RBN3704_n_26231), .b(n_25371), .c(FE_OCP_RBN2960_n_26231), .d(n_25342), .o(n_26933) );
na02f80 g753714 ( .a(n_26444), .b(n_26409), .o(n_26540) );
oa12f80 g777983 ( .a(n_2870), .b(n_3063), .c(n_3034), .o(n_3081) );
no02f80 g769605 ( .a(n_11383), .b(n_11394), .o(n_11415) );
ao12f80 g775157 ( .a(n_46427), .b(n_6008), .c(n_6007), .o(n_6039) );
in01f80 newInst_716 ( .a(newNet_715), .o(newNet_716) );
in01f80 g763964 ( .a(n_16799), .o(n_16853) );
no02f80 g737723 ( .a(n_42235), .b(n_42234), .o(n_42236) );
oa12f80 g778072 ( .a(n_2202), .b(n_2942), .c(n_2181), .o(n_3000) );
na02f80 g768369 ( .a(n_12540), .b(n_12564), .o(n_12577) );
no03m80 g765015 ( .a(n_16210), .b(n_16104), .c(n_15970), .o(n_16263) );
in01f80 FE_OCP_RBC2453_n_38537 ( .a(n_38537), .o(FE_OCP_RBN2453_n_38537) );
ao12f80 g762063 ( .a(n_18180), .b(n_18196), .c(n_18179), .o(n_19855) );
ao12f80 g780110 ( .a(n_732), .b(n_1029), .c(n_753), .o(n_1119) );
no02f80 g768656 ( .a(n_12195), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .o(n_12228) );
na02f80 g739575 ( .a(FE_OCP_RBN3336_n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .o(n_40622) );
in01f80 g759814 ( .a(n_21821), .o(n_21822) );
in01f80 g743850 ( .a(n_36071), .o(n_36103) );
na02f80 g738954 ( .a(n_41220), .b(n_40960), .o(n_41277) );
na02f80 FE_RC_1940_0 ( .a(FE_RN_618_0), .b(n_29063), .o(n_29118) );
in01f80 newInst_1108 ( .a(newNet_1107), .o(newNet_1108) );
in01f80 g749577 ( .a(n_31709), .o(n_31780) );
no02f80 g776433 ( .a(n_4266), .b(FE_OCPN846_n_4046), .o(n_4428) );
na02f80 g775390 ( .a(n_5437), .b(n_5056), .o(n_5528) );
in01f80 FE_OCP_RBC2181_n_1916 ( .a(n_1916), .o(FE_OCP_RBN2181_n_1916) );
in01f80 g737168 ( .a(n_43030), .o(n_43103) );
in01f80 g749293 ( .a(n_30630), .o(n_30657) );
in01f80 g777413 ( .a(n_3564), .o(n_3639) );
ao12f80 g756406 ( .a(n_23496), .b(n_23742), .c(n_23541), .o(n_23826) );
in01f80 g757586 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_3_), .o(n_22797) );
na02f80 g757924 ( .a(n_23056), .b(FE_OFN735_n_22641), .o(n_23083) );
in01f80 g781325 ( .a(n_78), .o(n_79) );
na02f80 g759592 ( .a(n_20642), .b(n_20553), .o(n_20729) );
oa12f80 g774603 ( .a(n_6222), .b(n_6373), .c(n_6244), .o(n_6388) );
in01f80 g755604 ( .a(n_24528), .o(n_25531) );
in01f80 g750678 ( .a(n_30703), .o(n_30832) );
in01f80 newInst_2867 ( .a(newNet_2866), .o(newNet_2867) );
in01f80 g775888 ( .a(n_5049), .o(n_5076) );
na02f80 g770010 ( .a(n_10876), .b(n_10908), .o(n_11005) );
ao22s80 FE_RC_3992_0 ( .a(FE_RN_1731_0), .b(FE_OCP_RBN2421_n_24505), .c(n_25104), .d(n_25016), .o(n_25127) );
in01f80 newInst_241 ( .a(newNet_240), .o(newNet_241) );
no02f80 FE_RC_4197_0 ( .a(FE_RN_1839_0), .b(n_19139), .o(n_19237) );
na02f80 g741049 ( .a(n_39359), .b(n_39425), .o(n_39457) );
ao12f80 g777956 ( .a(n_3070), .b(n_3069), .c(n_3068), .o(n_4662) );
na02f80 g739121 ( .a(n_41055), .b(n_41054), .o(n_41056) );
no02f80 g764256 ( .a(n_16431), .b(n_16430), .o(n_16514) );
oa12f80 g738935 ( .a(n_41242), .b(n_41241), .c(n_41240), .o(n_41320) );
no02f80 g750073 ( .a(n_29896), .b(n_29477), .o(n_30194) );
in01f80 g756177 ( .a(n_24246), .o(n_24223) );
in01f80 g780152 ( .a(n_1190), .o(n_1183) );
in01f80 FE_OCPC987_n_28402 ( .a(FE_OCPN986_n_28402), .o(FE_OCPN987_n_28402) );
no02f80 g736631 ( .a(n_43565), .b(n_43407), .o(n_43625) );
na02f80 g750306 ( .a(n_29764), .b(n_29729), .o(n_29793) );
na02f80 g743018 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_28_), .o(n_36996) );
na02f80 g754462 ( .a(n_25567), .b(FE_OCP_RBN3585_n_25295), .o(n_25633) );
na02f80 g737943 ( .a(n_42201), .b(n_42138), .o(n_42343) );
no02f80 g766734 ( .a(n_13726), .b(n_13662), .o(n_13728) );
in01f80 g768575 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_19_), .o(n_12327) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_29_ ( .ck(newNet_1202), .d(n_6384), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_) );
in01f80 newInst_1223 ( .a(newNet_1222), .o(newNet_1223) );
in01f80 g755615 ( .a(n_24621), .o(n_24650) );
no02f80 g777611 ( .a(n_3401), .b(n_2695), .o(n_3412) );
no02f80 g738037 ( .a(n_42139), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42140) );
no02f80 FE_RC_4026_0 ( .a(FE_RN_1748_0), .b(n_44211), .o(n_35575) );
ao12f80 g772892 ( .a(n_7338), .b(n_7731), .c(n_7355), .o(n_7798) );
na02f80 g752569 ( .a(n_27608), .b(n_27471), .o(n_27691) );
in01f80 newInst_1113 ( .a(newNet_1112), .o(newNet_1113) );
in01f80 newInst_454 ( .a(newNet_453), .o(newNet_454) );
in01f80 g783831 ( .a(n_45517), .o(n_45518) );
ao22s80 g773660 ( .a(n_7282), .b(n_6892), .c(n_7281), .d(n_6893), .o(n_7723) );
oa12f80 g736539 ( .a(n_43153), .b(n_43629), .c(n_43538), .o(n_43654) );
in01f80 newInst_473 ( .a(newNet_442), .o(newNet_473) );
na02f80 g776418 ( .a(n_4358), .b(n_4457), .o(n_4543) );
no02f80 g775737 ( .a(n_5335), .b(n_3922), .o(n_5440) );
no02f80 g739289 ( .a(n_40901), .b(n_40904), .o(n_41208) );
na02f80 FE_RC_4016_0 ( .a(n_14215), .b(FE_OCP_RBN3648_n_15281), .o(FE_RN_1744_0) );
no02f80 g770552 ( .a(FE_OCP_RBN2877_n_10354), .b(FE_OCP_RBN3680_n_10338), .o(n_10436) );
ao22s80 g747347 ( .a(n_32615), .b(n_44962), .c(FE_OCP_RBN3331_n_44962), .d(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .o(n_32663) );
ao12f80 g749897 ( .a(FE_OCP_RBN3011_n_31117), .b(n_31216), .c(n_31210), .o(n_31249) );
oa12f80 g776406 ( .a(n_4562), .b(n_4608), .c(n_4561), .o(n_4631) );
no02f80 g741254 ( .a(FE_OCP_RBN2685_n_38870), .b(n_38612), .o(n_39155) );
in01f80 newInst_1909 ( .a(newNet_1166), .o(newNet_1909) );
in01f80 newInst_248 ( .a(newNet_4), .o(newNet_248) );
in01f80 g746723 ( .a(n_33270), .o(n_33609) );
na02f80 g741896 ( .a(n_38335), .b(n_38334), .o(n_38336) );
ao22s80 FE_RC_4114_0 ( .a(n_28997), .b(n_28625), .c(n_28624), .d(n_28998), .o(n_29091) );
in01f80 g761051 ( .a(n_19407), .o(n_19408) );
in01f80 g742050 ( .a(n_37946), .o(n_37947) );
na02f80 FE_RC_2311_0 ( .a(n_34613), .b(FE_RN_876_0), .o(FE_RN_877_0) );
oa12f80 g736342 ( .a(n_43566), .b(n_43814), .c(n_43437), .o(n_43831) );
na02f80 g747742 ( .a(n_33601), .b(n_33600), .o(n_33602) );
in01f80 g747508 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_3_), .o(n_32591) );
no02f80 g742021 ( .a(n_37909), .b(n_44872), .o(n_37978) );
no02f80 g748893 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n_32444) );
na02f80 g747105 ( .a(n_32789), .b(n_32821), .o(n_32831) );
in01f80 g760438 ( .a(n_21251), .o(n_20699) );
in01f80 FE_OCPC1015_n_32820 ( .a(FE_OCPN1014_n_32820), .o(FE_OCPN1015_n_32820) );
na02f80 g756050 ( .a(n_25026), .b(n_25130), .o(n_25162) );
na02f80 g760982 ( .a(n_19217), .b(n_19153), .o(n_19277) );
in01f80 g780812 ( .a(n_513), .o(n_514) );
na02f80 g778310 ( .a(n_2796), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .o(n_2895) );
no02f80 g751053 ( .a(n_29995), .b(n_29600), .o(n_29996) );
no02f80 g742309 ( .a(n_37794), .b(n_37838), .o(n_37812) );
in01f80 FE_OCP_RBC3501_n_8187 ( .a(FE_OCP_RBN3500_n_8187), .o(FE_OCP_RBN3501_n_8187) );
ao12f80 g744561 ( .a(n_36681), .b(n_36622), .c(n_36178), .o(n_36682) );
oa12f80 g751853 ( .a(n_28793), .b(n_28943), .c(n_28942), .o(n_28945) );
no02f80 FE_RC_1919_0 ( .a(n_19184), .b(FE_RN_605_0), .o(n_19225) );
in01f80 g779638 ( .a(n_1497), .o(n_1498) );
ao12f80 g746063 ( .a(n_33832), .b(n_33831), .c(n_33830), .o(n_33904) );
na02f80 g777974 ( .a(n_3072), .b(n_3071), .o(n_3073) );
in01f80 g773425 ( .a(n_7554), .o(n_7582) );
in01f80 g764097 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17015) );
oa12f80 g755737 ( .a(n_23883), .b(n_24274), .c(FE_OCPN1470_n_23818), .o(n_24323) );
na02f80 g749127 ( .a(FE_OCP_RBN2889_n_46957), .b(n_27131), .o(n_30881) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_14_ ( .ck(newNet_1643), .d(n_27092), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_) );
ao12f80 g756285 ( .a(n_23991), .b(n_24609), .c(n_24006), .o(n_24707) );
na02f80 g739606 ( .a(FE_OCP_RBN3336_n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .o(n_40641) );
ao12f80 g774239 ( .a(n_6651), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .o(n_6932) );
no02f80 g773911 ( .a(n_6980), .b(n_6979), .o(n_6981) );
ao12f80 g749698 ( .a(n_31455), .b(n_31417), .c(n_31311), .o(n_31578) );
na02f80 g766059 ( .a(n_14737), .b(FE_OCP_RBN3584_n_14681), .o(n_14781) );
na02f80 g762836 ( .a(n_17597), .b(n_17135), .o(n_17629) );
in01f80 g742581 ( .a(n_37637), .o(n_37983) );
na02f80 g756269 ( .a(n_24080), .b(n_23682), .o(n_24122) );
oa12f80 g737851 ( .a(n_42416), .b(n_42547), .c(n_42323), .o(n_42693) );
na02f80 g745280 ( .a(n_35680), .b(FE_OCP_RBN2993_n_35539), .o(n_35769) );
na02f80 g753128 ( .a(n_27461), .b(n_27337), .o(n_27500) );
in01f80 newInst_940 ( .a(newNet_939), .o(newNet_940) );
na02f80 g741208 ( .a(FE_OCP_RBN2685_n_38870), .b(n_38633), .o(n_39150) );
in01f80 newInst_269 ( .a(newNet_268), .o(newNet_269) );
na02f80 g759917 ( .a(n_21051), .b(n_21105), .o(n_21106) );
in01f80 g770832 ( .a(n_9933), .o(n_10018) );
ao12f80 g743681 ( .a(n_37434), .b(n_37363), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_37435) );
ao12f80 g746566 ( .a(n_33237), .b(n_33254), .c(n_33236), .o(n_34096) );
na02f80 g761433 ( .a(n_18898), .b(n_18336), .o(n_18947) );
in01f80 g761196 ( .a(n_19166), .o(n_19167) );
no02f80 g750729 ( .a(n_29196), .b(n_28735), .o(n_29197) );
na02f80 g742909 ( .a(n_36961), .b(n_37075), .o(n_37122) );
na02f80 g764460 ( .a(n_16218), .b(FE_OCP_RBN2591_n_14460), .o(n_16436) );
na02f80 g767648 ( .a(n_12808), .b(n_12770), .o(n_12829) );
in01f80 g748409 ( .a(n_31787), .o(n_31821) );
in01f80 newInst_3011 ( .a(newNet_3010), .o(newNet_3011) );
in01f80 newInst_2378 ( .a(newNet_2377), .o(newNet_2378) );
in01f80 g750633 ( .a(FE_OCP_RBN2328_n_29378), .o(n_29398) );
no02f80 g748263 ( .a(FE_OCP_RBN3731_n_31819), .b(n_30557), .o(n_32326) );
no03m80 FE_RC_2916_0 ( .a(FE_RN_1268_0), .b(n_39607), .c(n_39596), .o(FE_RN_1269_0) );
in01f80 g755073 ( .a(n_25615), .o(n_25616) );
na02f80 g764326 ( .a(n_16322), .b(n_16274), .o(n_16372) );
na02f80 g766544 ( .a(n_14059), .b(FE_OCP_RBN2245_n_13017), .o(n_14240) );
na02f80 g761833 ( .a(n_19097), .b(n_19070), .o(n_19071) );
no02f80 g780833 ( .a(n_498), .b(n_508), .o(n_511) );
ao12f80 g761083 ( .a(n_20016), .b(n_19912), .c(n_19980), .o(n_21101) );
in01f80 g769147 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_5_), .o(n_11659) );
no02f80 g751154 ( .a(n_29932), .b(n_30030), .o(n_30059) );
in01f80 g773026 ( .a(n_8166), .o(n_8167) );
in01f80 newInst_1570 ( .a(newNet_1569), .o(newNet_1570) );
oa12f80 g749618 ( .a(n_31645), .b(n_31644), .c(n_31643), .o(n_31691) );
in01f80 newInst_3178 ( .a(newNet_3177), .o(newNet_3178) );
no02f80 g778483 ( .a(n_2431), .b(n_2348), .o(n_2479) );
na02f80 g737040 ( .a(n_43082), .b(n_43129), .o(n_43184) );
in01f80 g778383 ( .a(n_47024), .o(n_2869) );
no02f80 g774748 ( .a(n_6287), .b(n_6213), .o(n_6288) );
in01f80 g772824 ( .a(n_7905), .o(n_7943) );
no02f80 g741206 ( .a(FE_OCP_RBN3626_n_38870), .b(FE_OCP_RBN3504_n_38592), .o(n_39180) );
in01f80 FE_OCP_RBC2257_n_37844 ( .a(FE_OCP_RBN2255_n_37844), .o(FE_OCP_RBN2257_n_37844) );
no02f80 g749570 ( .a(n_30489), .b(n_30488), .o(n_30490) );
na02f80 g748765 ( .a(n_31328), .b(n_31327), .o(n_31441) );
no02f80 g776780 ( .a(FE_OCP_RBN2676_n_4061), .b(n_3966), .o(n_4164) );
na02f80 g784784 ( .a(n_5746), .b(FE_OCP_RBN2788_n_4294), .o(n_47270) );
no02f80 g778308 ( .a(n_2796), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_), .o(n_2849) );
in01f80 g754112 ( .a(n_26911), .o(n_26978) );
in01f80 newInst_2175 ( .a(newNet_2174), .o(newNet_2175) );
in01f80 FE_OFC807_n_46195 ( .a(n_46195), .o(FE_OFN807_n_46195) );
in01f80 g752009 ( .a(n_28192), .o(n_28146) );
in01f80 newInst_422 ( .a(newNet_421), .o(newNet_422) );
na02f80 g778270 ( .a(n_2633), .b(n_3125), .o(n_2646) );
in01f80 FE_OCP_RBC2487_n_3338 ( .a(n_3338), .o(FE_OCP_RBN2487_n_3338) );
na02f80 g776696 ( .a(n_4134), .b(n_4133), .o(n_4220) );
na02f80 g763252 ( .a(n_17005), .b(n_16904), .o(n_17047) );
in01f80 newInst_3004 ( .a(newNet_3003), .o(newNet_3004) );
na02f80 g760180 ( .a(n_20489), .b(n_20458), .o(n_20568) );
no02f80 g758052 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n_23181) );
oa12f80 g759958 ( .a(n_21374), .b(n_21591), .c(n_20699), .o(n_21592) );
oa22f80 FE_RC_781_0 ( .a(n_33492), .b(n_33060), .c(n_45627), .d(n_33059), .o(n_33567) );
no02f80 g741142 ( .a(n_38909), .b(n_38955), .o(n_38956) );
no02f80 g739464 ( .a(n_40668), .b(n_40667), .o(n_40672) );
na02f80 g767495 ( .a(FE_OCP_RBN2230_n_13141), .b(n_12910), .o(n_13234) );
no02f80 g741526 ( .a(n_38707), .b(FE_OCP_RBN2542_n_38721), .o(n_38720) );
na02f80 g759293 ( .a(n_20857), .b(n_45024), .o(n_20924) );
oa12f80 g784685 ( .a(n_3569), .b(n_3557), .c(n_3444), .o(n_47015) );
oa12f80 g772974 ( .a(n_7681), .b(n_7803), .c(n_7727), .o(n_7902) );
na02f80 g747662 ( .a(n_33298), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_33299) );
in01f80 g741035 ( .a(n_38895), .o(n_38896) );
in01f80 g759838 ( .a(FE_OCPN1482_n_22207), .o(n_22280) );
oa12f80 g780752 ( .a(n_400), .b(n_576), .c(n_416), .o(n_584) );
no02f80 g744159 ( .a(n_35566), .b(n_35546), .o(n_35709) );
no02f80 g758762 ( .a(n_21582), .b(n_20019), .o(n_21741) );
na02f80 g745291 ( .a(n_35890), .b(n_36122), .o(n_36172) );
in01f80 newInst_1890 ( .a(newNet_1889), .o(newNet_1890) );
no02f80 g752960 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .o(n_28176) );
ao12f80 g752014 ( .a(n_28793), .b(n_28862), .c(n_28856), .o(n_28877) );
no02f80 g777312 ( .a(n_3938), .b(n_3902), .o(n_4108) );
in01f80 g742571 ( .a(n_37535), .o(n_37556) );
oa22f80 FE_RC_1467_0 ( .a(n_17584), .b(n_17688), .c(n_16339), .d(n_44150), .o(n_17750) );
in01f80 g780491 ( .a(n_895), .o(n_896) );
in01f80 g738134 ( .a(n_42107), .o(n_42081) );
in01f80 FE_OCPC928_n_26231 ( .a(FE_OCPN927_n_26231), .o(FE_OCPN928_n_26231) );
no02f80 FE_RC_92_0 ( .a(FE_RN_29_0), .b(n_17084), .o(n_17072) );
no02f80 g774243 ( .a(n_6600), .b(n_6550), .o(n_6652) );
in01f80 g779450 ( .a(n_1438), .o(n_1439) );
in01f80 g770367 ( .a(n_10615), .o(n_10616) );
na02f80 g746418 ( .a(n_33331), .b(n_33024), .o(n_33388) );
na02f80 g743171 ( .a(n_36932), .b(n_36931), .o(n_36986) );
na02f80 g738434 ( .a(n_41431), .b(n_41430), .o(n_41432) );
in01f80 g764834 ( .a(n_15843), .o(n_15844) );
oa22f80 FE_RC_798_0 ( .a(FE_OCP_RBN3524_n_8242), .b(FE_OCP_RBN2479_n_8530), .c(n_8530), .d(FE_OCP_RBN3522_n_8242), .o(n_8580) );
in01f80 newInst_710 ( .a(newNet_709), .o(newNet_710) );
in01f80 FE_OCP_DRV_C1610_n_20146 ( .a(FE_OCP_DRV_N1609_n_20146), .o(FE_OCP_DRV_N1610_n_20146) );
no02f80 g752676 ( .a(n_28082), .b(n_27876), .o(n_28138) );
no02f80 g749709 ( .a(n_31414), .b(n_31407), .o(n_31415) );
in01f80 g743964 ( .a(n_35865), .o(n_35866) );
no02f80 g769257 ( .a(FE_OCP_RBN3093_n_11475), .b(n_10915), .o(n_11622) );
na02f80 g780482 ( .a(n_1111), .b(n_750), .o(n_1148) );
no02f80 g779616 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .o(n_2083) );
na02f80 g764165 ( .a(n_16494), .b(n_16564), .o(n_16555) );
in01f80 g765239 ( .a(n_15026), .o(n_15059) );
in01f80 g740988 ( .a(n_39135), .o(n_39252) );
na02f80 g775078 ( .a(n_6051), .b(n_5175), .o(n_6070) );
no04s80 g757003 ( .a(FE_OCPN1017_n_23307), .b(n_23023), .c(n_23138), .d(n_23308), .o(n_23237) );
no02f80 g760864 ( .a(n_19333), .b(n_18540), .o(n_19364) );
no02f80 g773004 ( .a(n_7752), .b(n_8444), .o(n_7753) );
no02f80 g767802 ( .a(n_13038), .b(n_13113), .o(n_13256) );
no02f80 g737343 ( .a(n_42854), .b(n_42433), .o(n_42867) );
in01f80 g773637 ( .a(n_7330), .o(n_7331) );
oa22f80 g751086 ( .a(n_30097), .b(n_30038), .c(n_30156), .d(n_30104), .o(n_30288) );
in01f80 g738118 ( .a(n_42043), .o(n_42044) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_5_ ( .ck(newNet_3001), .d(n_1010), .o(delay_add_ln22_unr2_stage2_stallmux_q_5_) );
in01f80 newInst_3051 ( .a(newNet_3050), .o(newNet_3051) );
na02f80 g772940 ( .a(n_7912), .b(n_7866), .o(n_8004) );
in01f80 g754186 ( .a(n_26045), .o(n_26114) );
no02f80 g757299 ( .a(n_44066), .b(delay_xor_ln22_unr15_stage6_stallmux_q_11_), .o(n_23077) );
in01f80 FE_OFC783_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN781_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
no02f80 g754481 ( .a(n_26314), .b(n_26419), .o(n_26386) );
in01f80 g738195 ( .a(n_41980), .o(n_41981) );
no02f80 g764285 ( .a(n_16230), .b(n_14588), .o(n_16296) );
no02f80 g747000 ( .a(n_32822), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .o(n_32835) );
in01f80 FE_OCPC3768_FE_OCP_RBN2375_n_8221 ( .a(FE_OCP_RBN2375_n_8221), .o(FE_OCPN3768_FE_OCP_RBN2375_n_8221) );
oa22f80 FE_RC_2956_0 ( .a(FE_OFN803_n_46285), .b(n_11873), .c(FE_OCP_RBN3043_n_46337), .d(n_11841), .o(n_46359) );
oa12f80 g764812 ( .a(n_15887), .b(n_15888), .c(n_15886), .o(n_15978) );
na02f80 g742134 ( .a(n_38348), .b(n_38302), .o(n_38406) );
na02f80 g763472 ( .a(n_16987), .b(delay_add_ln22_unr11_stage5_stallmux_q_1_), .o(n_17025) );
no02f80 FE_RC_2775_0 ( .a(n_38167), .b(n_38187), .o(FE_RN_1183_0) );
in01f80 fopt783971 ( .a(FE_OCP_RBN2121_n_45224), .o(n_45685) );
in01f80 FE_RC_3304_0 ( .a(n_17970), .o(FE_RN_1455_0) );
in01f80 newInst_1514 ( .a(newNet_1513), .o(newNet_1514) );
in01f80 g739253 ( .a(n_41079), .o(n_41080) );
no02f80 g757444 ( .a(n_22987), .b(n_22934), .o(n_23036) );
no02f80 g768454 ( .a(n_12394), .b(n_12393), .o(n_12395) );
in01f80 FE_OCP_RBC2420_n_24505 ( .a(n_24505), .o(FE_OCP_RBN2420_n_24505) );
in01f80 g777680 ( .a(n_5109), .o(n_3381) );
na02f80 g765571 ( .a(n_15140), .b(n_15139), .o(n_15141) );
na02f80 g749099 ( .a(n_30881), .b(n_30861), .o(n_30960) );
na02f80 g741210 ( .a(n_38841), .b(n_38828), .o(n_38883) );
in01f80 g747495 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_31_), .o(n_32335) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_18_ ( .ck(newNet_3326), .d(n_32113), .o(delay_add_ln22_unr20_stage8_stallmux_q_18_) );
in01f80 g746944 ( .a(n_32961), .o(n_33021) );
oa22f80 FE_RC_3307_0 ( .a(n_36770), .b(n_36832), .c(n_36769), .d(n_36833), .o(n_36874) );
no02f80 g759474 ( .a(n_20884), .b(n_20936), .o(n_21000) );
in01f80 newInst_2734 ( .a(newNet_2733), .o(newNet_2734) );
in01f80 newInst_131 ( .a(newNet_130), .o(newNet_131) );
na02f80 g771647 ( .a(n_8972), .b(n_8970), .o(n_9074) );
no02f80 g759093 ( .a(n_21350), .b(n_21389), .o(n_21537) );
ao12f80 g749753 ( .a(n_30211), .b(n_30242), .c(FE_OCPN1786_n_30134), .o(n_30297) );
na02f80 g749635 ( .a(n_30226), .b(n_30225), .o(n_30227) );
in01f80 newInst_755 ( .a(newNet_600), .o(newNet_755) );
na02f80 g753283 ( .a(FE_OCPN964_n_27287), .b(FE_OCP_RBN2968_n_26398), .o(n_27410) );
no02f80 g760926 ( .a(n_19416), .b(n_18913), .o(n_19424) );
oa22f80 g737264 ( .a(n_42876), .b(n_42679), .c(n_42918), .d(n_42680), .o(n_42954) );
na02f80 g779528 ( .a(n_1358), .b(n_1369), .o(n_1404) );
no03m80 FE_RC_1537_0 ( .a(n_40932), .b(n_41229), .c(n_41216), .o(n_41294) );
ao12f80 g750913 ( .a(n_29013), .b(n_29012), .c(n_29011), .o(n_29081) );
na02f80 g737042 ( .a(n_43046), .b(n_43104), .o(n_43128) );
ao12f80 g751074 ( .a(n_30092), .b(n_30303), .c(n_30063), .o(n_30412) );
na02f80 g737922 ( .a(n_42201), .b(n_41961), .o(n_42328) );
in01f80 newInst_2739 ( .a(newNet_2738), .o(newNet_2739) );
in01f80 g740431 ( .a(n_40238), .o(n_40239) );
in01f80 g777293 ( .a(n_5188), .o(n_5189) );
no02f80 FE_RC_2259_0 ( .a(FE_RN_835_0), .b(n_28401), .o(n_28399) );
na02f80 g749136 ( .a(n_30935), .b(n_30936), .o(n_30956) );
in01f80 g742246 ( .a(n_37867), .o(n_37868) );
in01f80 g759079 ( .a(n_21195), .o(n_21227) );
na02f80 g766082 ( .a(n_14515), .b(n_14471), .o(n_14616) );
oa12f80 g770657 ( .a(n_9985), .b(n_10068), .c(FE_OCP_RBN3635_n_47260), .o(n_10200) );
in01f80 g763379 ( .a(n_17329), .o(n_17326) );
no02f80 g763936 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .o(n_17572) );
no02f80 g764566 ( .a(n_15915), .b(n_14419), .o(n_15954) );
na02f80 g764688 ( .a(n_15896), .b(n_15737), .o(n_15986) );
in01f80 g747275 ( .a(n_33724), .o(n_33725) );
no02f80 g741863 ( .a(n_38287), .b(n_38026), .o(n_38413) );
in01f80 g757661 ( .a(n_22746), .o(n_22747) );
in01f80 newInst_2611 ( .a(newNet_232), .o(newNet_2611) );
in01f80 newInst_875 ( .a(newNet_874), .o(newNet_875) );
no02f80 g783847 ( .a(n_25707), .b(n_25678), .o(n_45533) );
no02f80 g739148 ( .a(n_40989), .b(n_40963), .o(n_41026) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_2_ ( .ck(newNet_1815), .d(n_16408), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_) );
in01f80 g746946 ( .a(n_32942), .o(n_32943) );
in01f80 newInst_1064 ( .a(newNet_628), .o(newNet_1064) );
na02f80 g746378 ( .a(n_33411), .b(n_32958), .o(n_33475) );
na02f80 g771761 ( .a(n_8980), .b(n_44575), .o(n_9005) );
oa22f80 g746429 ( .a(n_33346), .b(n_33302), .c(n_33347), .d(n_33301), .o(n_33426) );
na02f80 g760358 ( .a(n_20224), .b(n_20190), .o(n_20236) );
in01f80 g756389 ( .a(n_23973), .o(n_24016) );
ao12f80 g756317 ( .a(n_24544), .b(n_24587), .c(n_24543), .o(n_25129) );
na02f80 FE_RC_1864_0 ( .a(n_28182), .b(n_28234), .o(FE_RN_573_0) );
no02f80 g767894 ( .a(n_12905), .b(n_12914), .o(n_13064) );
na02f80 g737894 ( .a(n_42270), .b(n_42122), .o(n_42406) );
oa12f80 g747090 ( .a(n_34001), .b(n_34000), .c(n_33999), .o(n_34611) );
in01f80 newInst_1264 ( .a(newNet_1263), .o(newNet_1264) );
in01f80 g760498 ( .a(n_20026), .o(n_20078) );
no02f80 FE_RC_1186_0 ( .a(FE_RN_357_0), .b(FE_RN_358_0), .o(FE_RN_359_0) );
no02f80 g771848 ( .a(n_9694), .b(n_9591), .o(n_10576) );
in01f80 g771989 ( .a(n_9225), .o(n_9226) );
in01f80 g776945 ( .a(n_3977), .o(n_4498) );
na02f80 g736744 ( .a(n_43189), .b(n_43165), .o(n_43225) );
in01f80 g742721 ( .a(n_37398), .o(n_37910) );
in01f80 g741586 ( .a(n_38655), .o(n_38681) );
oa22f80 g775690 ( .a(n_5410), .b(n_5224), .c(n_5332), .d(n_5225), .o(n_5527) );
na02f80 g769967 ( .a(n_10957), .b(n_10995), .o(n_10996) );
in01f80 fopt782821 ( .a(n_44223), .o(n_44222) );
na02f80 g778704 ( .a(FE_OCP_RBN2290_n_2438), .b(n_2562), .o(n_2701) );
ao12f80 g773439 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .c(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n_7537) );
na02f80 g750425 ( .a(n_29596), .b(n_29549), .o(n_29612) );
in01f80 g775703 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n_5471) );
ao12f80 g769198 ( .a(n_12003), .b(n_10458), .c(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11632) );
no02f80 g770908 ( .a(FE_OCPN1255_n_8499), .b(n_9864), .o(n_9930) );
na02f80 g751552 ( .a(n_28460), .b(n_28523), .o(n_28600) );
in01f80 FE_OCP_RBC2916_n_10644 ( .a(n_10644), .o(FE_OCP_RBN2916_n_10644) );
in01f80 g772009 ( .a(n_9385), .o(n_9386) );
ao22s80 FE_RC_366_0 ( .a(n_47212), .b(n_11816), .c(n_47213), .d(n_11815), .o(n_12261) );
na02f80 g745522 ( .a(n_34320), .b(n_33385), .o(n_34346) );
in01f80 FE_OCP_RBC3845_FE_RN_1242_0 ( .a(FE_OCP_RBN3844_FE_RN_1242_0), .o(FE_OCP_RBN3845_FE_RN_1242_0) );
in01f80 FE_OCPC1530_n_26090 ( .a(FE_OCPN1529_n_26090), .o(FE_OCPN1530_n_26090) );
na02f80 g757094 ( .a(n_23301), .b(n_23214), .o(n_23346) );
in01f80 g741957 ( .a(n_38185), .o(n_38186) );
in01f80 newInst_3210 ( .a(newNet_3209), .o(newNet_3210) );
na02f80 g776196 ( .a(FE_OCP_RBN2790_n_4462), .b(n_4237), .o(n_4534) );
na02f80 g773404 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .o(n_7569) );
no02f80 g762452 ( .a(FE_OCP_RBN2147_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .o(n_17977) );
na02f80 g742495 ( .a(n_37656), .b(n_37655), .o(n_37715) );
ao12f80 g780768 ( .a(n_559), .b(n_558), .c(n_557), .o(n_678) );
na02f80 g779550 ( .a(n_1365), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1426) );
oa12f80 g778399 ( .a(n_2081), .b(n_2400), .c(n_2059), .o(n_2524) );
no02f80 g738589 ( .a(n_41876), .b(n_41532), .o(n_42083) );
ao22s80 g781007 ( .a(n_272), .b(n_142), .c(n_259), .d(n_141), .o(n_485) );
oa12f80 g762298 ( .a(n_18015), .b(n_18130), .c(n_17964), .o(n_18194) );
na02f80 g758031 ( .a(n_22227), .b(n_22266), .o(n_22379) );
na02f80 g768739 ( .a(n_12129), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_), .o(n_12248) );
in01f80 g760656 ( .a(n_19775), .o(n_19776) );
in01f80 FE_OFC76_n_5397 ( .a(n_5398), .o(FE_OFN76_n_5397) );
in01f80 g773735 ( .a(n_7262), .o(n_7263) );
ao12f80 g738312 ( .a(n_41822), .b(n_41648), .c(n_41820), .o(n_42191) );
na02f80 g784756 ( .a(n_8073), .b(n_47239), .o(n_47242) );
no02f80 g738538 ( .a(n_41508), .b(n_41507), .o(n_41509) );
in01f80 newInst_1546 ( .a(newNet_1545), .o(newNet_1546) );
oa12f80 g766695 ( .a(n_13789), .b(n_13836), .c(FE_OCP_RBN2246_n_13017), .o(n_13887) );
in01f80 g776042 ( .a(n_5032), .o(n_5033) );
in01f80 g774534 ( .a(n_6491), .o(n_6513) );
in01f80 g771946 ( .a(n_9693), .o(n_9694) );
ao12f80 g757910 ( .a(n_23084), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .o(n_23591) );
in01f80 newInst_795 ( .a(newNet_794), .o(newNet_795) );
in01f80 g751115 ( .a(n_30546), .o(n_30614) );
in01f80 g750788 ( .a(n_29215), .o(n_29216) );
in01f80 g751336 ( .a(n_29938), .o(n_29534) );
no02f80 g761539 ( .a(n_18754), .b(n_18716), .o(n_18798) );
in01f80 g737827 ( .a(n_42367), .o(n_42392) );
in01f80 FE_OCP_RBC3709_n_46337 ( .a(FE_OCP_RBN3039_n_46337), .o(FE_OCP_RBN3709_n_46337) );
no02f80 g762349 ( .a(n_45120), .b(n_18448), .o(n_18497) );
oa22f80 g739870 ( .a(n_40164), .b(n_40320), .c(n_40165), .d(n_40321), .o(n_40416) );
in01f80 g749555 ( .a(n_31502), .o(n_30553) );
no02f80 g741450 ( .a(n_38763), .b(n_38707), .o(n_38784) );
na02f80 g757307 ( .a(n_23438), .b(n_23437), .o(n_23450) );
oa12f80 g753699 ( .a(n_26527), .b(n_26526), .c(n_26525), .o(n_26582) );
no02f80 g742552 ( .a(n_37527), .b(n_37709), .o(n_37659) );
no02f80 g740884 ( .a(n_39373), .b(n_39343), .o(n_39844) );
in01f80 g756911 ( .a(n_23328), .o(n_23379) );
na02f80 g747737 ( .a(n_33357), .b(n_33334), .o(n_33358) );
oa12f80 g750959 ( .a(n_28509), .b(n_28967), .c(n_28510), .o(n_29012) );
oa12f80 g758566 ( .a(n_21799), .b(n_22525), .c(n_21753), .o(n_22604) );
ao12f80 g777714 ( .a(n_3315), .b(n_3326), .c(n_3314), .o(n_5168) );
na02f80 g739012 ( .a(n_41124), .b(n_41438), .o(n_41125) );
na02f80 g770233 ( .a(FE_OCP_RBN2890_n_10568), .b(FE_OCP_RBN3645_n_44490), .o(n_10622) );
in01f80 g765807 ( .a(n_14830), .o(n_14889) );
na02f80 g770055 ( .a(n_10851), .b(n_10832), .o(n_10908) );
no02f80 g755538 ( .a(n_24712), .b(n_24775), .o(n_24832) );
na02f80 g738155 ( .a(n_42005), .b(n_41908), .o(n_42070) );
ao12f80 g740765 ( .a(FE_OCP_RBN2602_n_39126), .b(n_39493), .c(n_39121), .o(n_39514) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_21_ ( .ck(newNet_3222), .d(n_36430), .o(delay_add_ln22_unr23_stage9_stallmux_q_21_) );
na02f80 FE_RC_1947_0 ( .a(n_24458), .b(n_25486), .o(FE_RN_623_0) );
no02f80 g779739 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .o(n_1643) );
in01f80 g780781 ( .a(n_545), .o(n_546) );
in01f80 newInst_3030 ( .a(newNet_3029), .o(newNet_3030) );
na02f80 g759107 ( .a(n_21386), .b(n_21147), .o(n_21420) );
no02f80 g745586 ( .a(n_34291), .b(n_34323), .o(n_34354) );
no02f80 FE_RC_270_0 ( .a(n_44277), .b(n_22082), .o(FE_RN_81_0) );
in01f80 g781150 ( .a(n_202), .o(n_203) );
no02f80 FE_RC_3025_0 ( .a(n_20744), .b(n_21067), .o(FE_RN_1325_0) );
na02f80 g773974 ( .a(n_6918), .b(n_5139), .o(n_7010) );
in01f80 g767313 ( .a(n_13413), .o(n_13410) );
na02f80 g757336 ( .a(n_23105), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .o(n_23188) );
in01f80 newInst_3636 ( .a(newNet_3635), .o(newNet_3636) );
in01f80 newInst_338 ( .a(newNet_337), .o(newNet_338) );
in01f80 newInst_3534 ( .a(newNet_2131), .o(newNet_3534) );
in01f80 g775970 ( .a(n_5152), .o(n_5201) );
no02f80 g755997 ( .a(n_25160), .b(n_25129), .o(n_25570) );
na02f80 g778352 ( .a(n_2585), .b(n_2474), .o(n_2633) );
in01f80 FE_OCPC1383_n_18345 ( .a(n_18345), .o(FE_OCPN1383_n_18345) );
in01f80 FE_RC_3533_0 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .o(FE_RN_1528_0) );
in01f80 FE_OCPC1800_FE_OFN780_n_17093 ( .a(FE_OCPN1799_FE_OFN780_n_17093), .o(FE_OCPN1800_FE_OFN780_n_17093) );
in01f80 newInst_631 ( .a(newNet_293), .o(newNet_631) );
in01f80 g754585 ( .a(n_26894), .o(n_26895) );
no02f80 g762027 ( .a(n_18426), .b(n_18425), .o(n_18458) );
in01f80 g764409 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .o(n_16617) );
in01f80 g743976 ( .a(n_36196), .o(n_36197) );
in01f80 g769086 ( .a(n_11808), .o(n_11809) );
ao12f80 g749812 ( .a(n_31322), .b(n_31311), .c(n_31251), .o(n_31567) );
in01f80 FE_OCPC1425_n_18099 ( .a(n_18099), .o(FE_OCPN1425_n_18099) );
oa12f80 g742718 ( .a(n_37149), .b(n_37409), .c(n_37038), .o(n_37457) );
na02f80 g762384 ( .a(n_45118), .b(n_18441), .o(n_18664) );
in01f80 g748724 ( .a(n_31142), .o(n_31160) );
in01f80 g744559 ( .a(n_36683), .o(n_36684) );
no02f80 FE_RC_768_0 ( .a(n_33810), .b(FE_RN_239_0), .o(n_46955) );
in01f80 newInst_1643 ( .a(newNet_1642), .o(newNet_1643) );
oa12f80 g777824 ( .a(n_3242), .b(n_3260), .c(n_2759), .o(n_3321) );
na02f80 g758678 ( .a(n_21792), .b(n_21687), .o(n_21813) );
no02f80 g737740 ( .a(n_42285), .b(n_41917), .o(n_42377) );
in01f80 g768538 ( .a(n_12368), .o(n_12348) );
in01f80 FE_OCP_RBC2680_n_14768 ( .a(n_14768), .o(FE_OCP_RBN2680_n_14768) );
na02f80 g772594 ( .a(n_8305), .b(n_7860), .o(n_8372) );
in01f80 g736947 ( .a(n_43255), .o(n_43307) );
no02f80 g744500 ( .a(n_35411), .b(n_35404), .o(n_35470) );
in01f80 g744015 ( .a(n_36299), .o(n_36300) );
na02f80 g767777 ( .a(n_12791), .b(n_12836), .o(n_12837) );
na02f80 g764868 ( .a(n_15557), .b(FE_OCPN1007_n_13962), .o(n_15591) );
no02f80 g778324 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_30_), .o(n_4073) );
no02f80 g775308 ( .a(n_5636), .b(n_5469), .o(n_5637) );
no02f80 g771545 ( .a(n_9781), .b(n_9605), .o(n_9443) );
no02f80 g767698 ( .a(n_13088), .b(n_13040), .o(n_13156) );
no02f80 FE_RC_2867_0 ( .a(n_33882), .b(FE_RN_1236_0), .o(n_33969) );
na02f80 g744671 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_36557) );
na02f80 g781340 ( .a(n_7), .b(beta_23), .o(n_72) );
no02f80 g766615 ( .a(n_13915), .b(n_13894), .o(n_14018) );
in01f80 FE_OCP_RBC2465_n_4336 ( .a(FE_OCP_RBN2464_n_4336), .o(FE_OCP_RBN2465_n_4336) );
in01f80 newInst_1730 ( .a(newNet_1729), .o(newNet_1730) );
ao12f80 g768273 ( .a(n_12568), .b(n_12573), .c(n_12567), .o(n_12964) );
oa12f80 g756068 ( .a(n_24284), .b(n_24306), .c(n_24283), .o(n_24390) );
na02f80 g752661 ( .a(n_28138), .b(n_27904), .o(n_28205) );
in01f80 newInst_560 ( .a(newNet_367), .o(newNet_560) );
in01f80 g736521 ( .a(n_43722), .o(n_43735) );
in01f80 newInst_1321 ( .a(newNet_1320), .o(newNet_1321) );
na02f80 g739413 ( .a(FE_OCPN897_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n_41013) );
ao12f80 g769238 ( .a(n_12082), .b(n_45659), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n_12429) );
no02f80 g754080 ( .a(n_26069), .b(n_25651), .o(n_26070) );
in01f80 g754722 ( .a(n_26637), .o(n_26638) );
in01f80 g753469 ( .a(n_26786), .o(n_26787) );
na02f80 g739237 ( .a(n_41040), .b(n_40691), .o(n_41116) );
na02f80 g739953 ( .a(n_39960), .b(n_39927), .o(n_40049) );
in01f80 newInst_1860 ( .a(newNet_632), .o(newNet_1860) );
na02f80 g773705 ( .a(n_7272), .b(n_6123), .o(n_7355) );
na02f80 FE_RC_3067_0 ( .a(FE_RN_1346_0), .b(FE_RN_1348_0), .o(n_20926) );
no02f80 g771816 ( .a(n_8868), .b(n_8867), .o(n_8869) );
na02f80 g751916 ( .a(n_29099), .b(n_29305), .o(n_29711) );
in01f80 g744548 ( .a(n_35385), .o(n_35386) );
in01f80 g770067 ( .a(n_10932), .o(n_10933) );
no02f80 g766325 ( .a(n_14199), .b(n_14182), .o(n_14281) );
in01f80 g755915 ( .a(n_25708), .o(n_25709) );
oa12f80 g768727 ( .a(n_12126), .b(n_12125), .c(n_12124), .o(n_12247) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_16_ ( .ck(newNet_2306), .d(n_40433), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_) );
in01f80 g745706 ( .a(n_34245), .o(n_34246) );
in01f80 g778158 ( .a(n_2938), .o(n_2896) );
na02f80 g744882 ( .a(n_34978), .b(n_30633), .o(n_35010) );
na02f80 g741963 ( .a(n_44036), .b(n_37987), .o(n_37988) );
in01f80 g778739 ( .a(n_2758), .o(n_2834) );
na02f80 g755174 ( .a(n_25023), .b(n_25022), .o(n_25105) );
in01f80 g740537 ( .a(n_39698), .o(n_39699) );
na02f80 g768056 ( .a(FE_OCPN860_n_12880), .b(n_12850), .o(n_13159) );
no02f80 g760962 ( .a(n_19270), .b(n_18032), .o(n_19282) );
in01f80 g757494 ( .a(n_23040), .o(n_22985) );
no02f80 g754416 ( .a(n_25704), .b(n_25453), .o(n_25733) );
in01f80 g742428 ( .a(n_37707), .o(n_37719) );
no02f80 g759233 ( .a(n_21801), .b(n_21835), .o(n_21837) );
in01f80 g748339 ( .a(n_31893), .o(n_31894) );
in01f80 newInst_1886 ( .a(newNet_1885), .o(newNet_1886) );
na02f80 g770739 ( .a(n_10018), .b(n_10017), .o(n_10019) );
na02f80 g762195 ( .a(n_18194), .b(n_18168), .o(n_18169) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_24_ ( .ck(newNet_2465), .d(n_32463), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_) );
ao12f80 g750493 ( .a(n_30481), .b(n_30480), .c(n_30479), .o(n_31171) );
na02f80 g780689 ( .a(n_648), .b(n_515), .o(n_657) );
in01f80 g766338 ( .a(n_14398), .o(n_14399) );
in01f80 FE_OCP_RBC2758_FE_RN_722_0 ( .a(FE_RN_722_0), .o(FE_OCP_RBN2758_FE_RN_722_0) );
in01f80 newInst_1833 ( .a(newNet_1832), .o(newNet_1833) );
na02f80 g757249 ( .a(n_23469), .b(n_22852), .o(n_23492) );
ao12f80 g760383 ( .a(n_20743), .b(n_20742), .c(n_20741), .o(n_21370) );
oa12f80 g764335 ( .a(n_16018), .b(n_16673), .c(n_15967), .o(n_16742) );
no02f80 g754560 ( .a(n_26861), .b(n_26608), .o(n_26899) );
na02f80 FE_RC_2963_0 ( .a(FE_RN_1293_0), .b(FE_OCP_RBN2775_n_10100), .o(FE_RN_1294_0) );
in01f80 g771881 ( .a(n_8905), .o(n_8927) );
in01f80 newInst_1929 ( .a(newNet_1928), .o(newNet_1929) );
in01f80 g745106 ( .a(n_34788), .o(n_34858) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_9_ ( .ck(newNet_2038), .d(n_5527), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_) );
na02f80 g762697 ( .a(n_18237), .b(n_18211), .o(n_18212) );
in01f80 FE_OCP_RBC3613_n_20249 ( .a(FE_OCP_RBN2670_n_20249), .o(FE_OCP_RBN3613_n_20249) );
ao12f80 g766766 ( .a(n_13173), .b(n_13645), .c(n_13213), .o(n_13695) );
na02f80 g781062 ( .a(cos_out_26), .b(FE_OFN1_n_43918), .o(n_337) );
na02f80 g736751 ( .a(n_43529), .b(n_43113), .o(n_43114) );
in01f80 FE_OCP_RBC3514_n_13960 ( .a(FE_OCP_RBN3513_n_13960), .o(FE_OCP_RBN3514_n_13960) );
oa22f80 FE_RC_1668_0 ( .a(FE_OCP_RBN3466_n_7886), .b(n_8321), .c(FE_OCPN890_n_7802), .d(n_8322), .o(n_8462) );
no02f80 g764189 ( .a(n_16443), .b(n_16435), .o(n_16497) );
na02f80 g774377 ( .a(n_6944), .b(n_6721), .o(n_6962) );
no02f80 g778617 ( .a(n_2635), .b(n_2634), .o(n_2990) );
no02f80 g766890 ( .a(n_14259), .b(n_14758), .o(n_14300) );
in01f80 g760013 ( .a(n_21406), .o(n_21691) );
na02f80 g769696 ( .a(n_11243), .b(n_11157), .o(n_11295) );
ao12f80 g756256 ( .a(n_24630), .b(n_24629), .c(n_24628), .o(n_25133) );
na02f80 g747671 ( .a(n_32279), .b(n_32078), .o(n_32298) );
in01f80 g757695 ( .a(n_23244), .o(n_23220) );
in01f80 FE_OCP_RBC3529_n_13765 ( .a(FE_OCP_RBN3527_n_13765), .o(FE_OCP_RBN3529_n_13765) );
in01f80 g760770 ( .a(n_19715), .o(n_19716) );
in01f80 g750855 ( .a(n_29188), .o(n_29372) );
in01f80 newInst_1576 ( .a(newNet_1575), .o(newNet_1576) );
oa12f80 g768721 ( .a(n_11580), .b(n_11989), .c(n_11712), .o(n_11990) );
oa12f80 g750348 ( .a(n_29587), .b(n_29687), .c(n_29622), .o(n_29735) );
no02f80 g744844 ( .a(n_35005), .b(n_30612), .o(n_35035) );
in01f80 fopt783210 ( .a(FE_OCP_RBN3309_n_44722), .o(n_44763) );
oa12f80 g743891 ( .a(n_35565), .b(n_35573), .c(n_35599), .o(n_35712) );
oa22f80 FE_RC_827_0 ( .a(n_24051), .b(n_24406), .c(n_24050), .d(n_24405), .o(n_24505) );
in01f80 newInst_2644 ( .a(newNet_2643), .o(newNet_2644) );
oa12f80 g767451 ( .a(n_12951), .b(n_13462), .c(n_13033), .o(n_13521) );
in01f80 newInst_3141 ( .a(newNet_3140), .o(newNet_3141) );
in01f80 g759367 ( .a(n_20926), .o(n_20861) );
in01f80 g763149 ( .a(n_17579), .o(n_17616) );
oa12f80 g747763 ( .a(n_32028), .b(n_32188), .c(n_31902), .o(n_32277) );
ao22s80 g736686 ( .a(n_43055), .b(n_43041), .c(n_43056), .d(n_43040), .o(n_43115) );
na02f80 g737541 ( .a(n_42264), .b(n_42263), .o(n_42318) );
in01f80 g758616 ( .a(n_21921), .o(n_21936) );
na02f80 g737201 ( .a(n_42949), .b(n_42816), .o(n_42976) );
in01f80 g780992 ( .a(n_354), .o(n_357) );
in01f80 g746792 ( .a(n_33184), .o(n_33185) );
in01f80 g777366 ( .a(n_4193), .o(n_4194) );
na02f80 g766888 ( .a(n_14216), .b(n_14215), .o(n_14306) );
in01f80 fopt783481 ( .a(n_45091), .o(n_45070) );
no02f80 g765538 ( .a(FE_OCP_RBN2713_n_14982), .b(FE_OCP_RBN1170_n_13756), .o(n_15049) );
oa22f80 g737300 ( .a(n_42847), .b(n_42767), .c(n_42862), .d(n_42768), .o(n_42922) );
ao12f80 g784394 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .o(n_46205) );
in01f80 g752266 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .o(n_27871) );
in01f80 FE_OCP_RBC2476_n_8599 ( .a(n_8599), .o(FE_OCP_RBN2476_n_8599) );
no02f80 g776176 ( .a(n_4459), .b(FE_OCPN960_n_3951), .o(n_4523) );
na02f80 g777624 ( .a(n_3389), .b(n_3190), .o(n_3452) );
in01f80 FE_OCP_RBC3027_n_39942 ( .a(FE_OCP_RBN3023_n_39942), .o(FE_OCP_RBN3027_n_39942) );
in01f80 FE_OFC757_n_45813 ( .a(n_45813), .o(FE_OFN757_n_45813) );
na02f80 g769685 ( .a(n_11223), .b(n_44498), .o(n_11246) );
in01f80 g765389 ( .a(n_15055), .o(n_15056) );
no02f80 g759287 ( .a(n_21119), .b(n_21039), .o(n_21156) );
na02f80 g774914 ( .a(n_6101), .b(n_6102), .o(n_6151) );
in01f80 g743952 ( .a(n_36320), .o(n_36321) );
in01f80 FE_OCPC1400_n_8670 ( .a(FE_OCPN1399_n_8670), .o(FE_OCPN1400_n_8670) );
na02f80 g775624 ( .a(n_5736), .b(n_5662), .o(n_5761) );
no02f80 g780389 ( .a(n_860), .b(n_847), .o(n_950) );
no02f80 g761007 ( .a(n_19273), .b(n_19272), .o(n_19325) );
in01f80 g774965 ( .a(n_6203), .o(n_6204) );
oa12f80 g757866 ( .a(n_22445), .b(n_22448), .c(n_22352), .o(n_22472) );
in01f80 FE_RC_496_0 ( .a(n_28230), .o(FE_RN_148_0) );
na02f80 g767359 ( .a(n_13362), .b(n_13365), .o(n_13416) );
no02f80 g752622 ( .a(n_27568), .b(n_27275), .o(n_27593) );
no02f80 g759732 ( .a(n_20320), .b(n_20298), .o(n_20420) );
no02f80 g750337 ( .a(n_29730), .b(n_29551), .o(n_29762) );
ao12f80 g752153 ( .a(n_28010), .b(FE_OCPN877_n_44734), .c(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .o(n_28040) );
in01f80 g736972 ( .a(n_43342), .o(n_43343) );
no02f80 g764202 ( .a(n_47340), .b(n_14783), .o(n_16561) );
na02f80 g763917 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .o(n_17098) );
na02f80 g761341 ( .a(n_20219), .b(n_20254), .o(n_21020) );
in01f80 g768780 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .o(n_12254) );
in01f80 FE_OCPC888_n_42367 ( .a(FE_OCPN886_n_42367), .o(FE_OCPN888_n_42367) );
in01f80 g777657 ( .a(n_3528), .o(n_3529) );
no02f80 g776843 ( .a(n_3987), .b(FE_OCP_RBN2649_n_3840), .o(n_4061) );
na02f80 g751799 ( .a(n_28911), .b(n_28840), .o(n_28930) );
in01f80 g739127 ( .a(n_41028), .o(n_41401) );
in01f80 g775844 ( .a(n_4964), .o(n_4965) );
na02f80 g779181 ( .a(n_1939), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .o(n_2006) );
na02f80 g769362 ( .a(FE_OCPN867_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .o(n_11892) );
in01f80 g755418 ( .a(n_24760), .o(n_24878) );
in01f80 g748114 ( .a(n_31744), .o(n_31745) );
in01f80 newInst_1974 ( .a(newNet_912), .o(newNet_1974) );
na02f80 g766440 ( .a(n_14117), .b(n_14243), .o(n_14229) );
in01f80 g764385 ( .a(n_16677), .o(n_16678) );
oa12f80 g754598 ( .a(FE_OCP_RBN2966_n_26231), .b(n_26680), .c(n_26679), .o(n_26793) );
ao22s80 g781115 ( .a(n_226), .b(n_125), .c(n_225), .d(n_126), .o(n_549) );
oa12f80 g768604 ( .a(n_12130), .b(n_12292), .c(n_12041), .o(n_12341) );
ao22s80 g751931 ( .a(n_28186), .b(n_28180), .c(n_28141), .d(n_28179), .o(n_29375) );
in01f80 g763266 ( .a(n_17334), .o(n_17440) );
na02f80 g743129 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n_37149) );
in01f80 FE_OCPC1254_n_8499 ( .a(FE_OCP_RBN3519_n_8498), .o(FE_OCPN1254_n_8499) );
ao12f80 g753501 ( .a(n_26581), .b(n_26781), .c(n_26473), .o(n_26848) );
na02f80 g766538 ( .a(FE_OCP_RBN2401_n_13954), .b(n_13376), .o(n_14025) );
na02f80 g765309 ( .a(n_15961), .b(n_15874), .o(n_16017) );
in01f80 g776318 ( .a(n_4811), .o(n_4812) );
in01f80 newInst_909 ( .a(newNet_908), .o(newNet_909) );
in01f80 newInst_856 ( .a(newNet_855), .o(newNet_856) );
ao12f80 g736472 ( .a(n_43168), .b(FE_OCP_RBN3110_n_43711), .c(n_43515), .o(n_43752) );
in01f80 g748008 ( .a(n_33040), .o(n_33041) );
na02f80 g752028 ( .a(n_28086), .b(delay_add_ln22_unr17_stage7_stallmux_q_4_), .o(n_28183) );
in01f80 g740326 ( .a(n_40359), .o(n_40360) );
in01f80 g742937 ( .a(n_37061), .o(n_37062) );
no02f80 g772887 ( .a(n_7939), .b(n_7938), .o(n_7940) );
na02f80 g739906 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_5_), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40339) );
no02f80 g754376 ( .a(n_25807), .b(n_25778), .o(n_25889) );
no02f80 g784793 ( .a(n_15543), .b(n_15586), .o(n_47332) );
in01f80 g747285 ( .a(n_32784), .o(n_32785) );
oa22f80 FE_RC_1708_0 ( .a(n_17381), .b(n_17457), .c(n_17380), .d(n_17495), .o(n_17630) );
oa12f80 g772418 ( .a(n_7889), .b(n_8503), .c(n_7922), .o(n_8717) );
na02f80 g769725 ( .a(n_11170), .b(n_11114), .o(n_11224) );
ao12f80 g765370 ( .a(n_15829), .b(n_16245), .c(n_15833), .o(n_16249) );
in01f80 g753460 ( .a(n_27589), .o(n_27586) );
na02f80 g774845 ( .a(n_6202), .b(n_6208), .o(n_6313) );
na02f80 g745973 ( .a(n_33926), .b(n_33925), .o(n_33927) );
no02f80 g776863 ( .a(n_3630), .b(n_3624), .o(n_3732) );
in01f80 g748018 ( .a(n_32184), .o(n_32185) );
no02f80 g741160 ( .a(FE_OCP_RBN2639_n_38806), .b(n_38431), .o(n_38966) );
in01f80 g753993 ( .a(n_26184), .o(n_26185) );
no02f80 g755191 ( .a(n_25097), .b(n_25068), .o(n_25180) );
in01f80 g779765 ( .a(n_1543), .o(n_1549) );
in01f80 g775230 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .o(n_5999) );
na02f80 FE_RC_3896_0 ( .a(FE_RN_1690_0), .b(FE_RN_1691_0), .o(FE_RN_1692_0) );
ao12f80 g763078 ( .a(n_17547), .b(n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .o(n_17617) );
no02f80 g746532 ( .a(n_33168), .b(n_33166), .o(n_33167) );
in01f80 g756336 ( .a(n_24541), .o(n_25028) );
in01f80 g755304 ( .a(n_25528), .o(n_25529) );
na02f80 FE_RC_3154_0 ( .a(FE_RN_1399_0), .b(n_21186), .o(n_21470) );
in01f80 newInst_1025 ( .a(newNet_1024), .o(newNet_1025) );
in01f80 g768570 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n_12271) );
na02f80 g748133 ( .a(n_32782), .b(n_32781), .o(n_32804) );
in01f80 g767519 ( .a(n_13057), .o(n_13058) );
in01f80 g777884 ( .a(n_3309), .o(n_3310) );
in01f80 g740856 ( .a(n_39381), .o(n_39468) );
na02f80 g776978 ( .a(n_5356), .b(n_5355), .o(n_6304) );
in01f80 g751844 ( .a(n_29148), .o(n_29149) );
na02f80 g776721 ( .a(n_4075), .b(n_4088), .o(n_4247) );
na02f80 g736830 ( .a(n_43126), .b(n_46940), .o(n_43139) );
no02f80 g743434 ( .a(n_36569), .b(n_36750), .o(n_36570) );
in01f80 g747396 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .o(n_32402) );
in01f80 FE_OCP_RBC3106_n_22590 ( .a(n_22590), .o(FE_OCP_RBN3106_n_22590) );
na02f80 FE_RC_4148_0 ( .a(n_16988), .b(FE_RN_1803_0), .o(FE_RN_1804_0) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_0_ ( .ck(newNet_854), .d(n_1327), .o(delay_xor_ln21_unr3_stage2_stallmux_q_0_) );
no02f80 g769078 ( .a(n_11482), .b(n_11312), .o(n_11483) );
in01f80 g756442 ( .a(n_23775), .o(n_23739) );
no02f80 g773830 ( .a(n_7065), .b(n_6964), .o(n_7101) );
in01f80 g742063 ( .a(n_38008), .o(n_38009) );
no02f80 g771829 ( .a(n_9772), .b(n_9771), .o(n_9773) );
na02f80 g737193 ( .a(n_42977), .b(n_42988), .o(n_43000) );
in01f80 FE_OCP_RBC1851_n_22556 ( .a(n_22556), .o(FE_OCP_RBN1851_n_22556) );
no02f80 FE_RC_4195_0 ( .a(FE_RN_1837_0), .b(FE_RN_1838_0), .o(n_19107) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_25_ ( .ck(newNet_2933), .d(n_46993), .o(delay_add_ln22_unr5_stage3_stallmux_q_25_) );
in01f80 fopt782876 ( .a(n_44312), .o(n_44311) );
ao12f80 g760568 ( .a(n_19418), .b(n_19860), .c(n_19553), .o(n_19868) );
na02f80 FE_RC_2820_0 ( .a(FE_RN_1208_0), .b(n_34433), .o(FE_RN_1209_0) );
in01f80 g761368 ( .a(n_19988), .o(n_19902) );
no02f80 g774526 ( .a(n_6385), .b(n_6228), .o(n_6425) );
oa22f80 FE_RC_1109_0 ( .a(n_40643), .b(n_40659), .c(n_40644), .d(n_40664), .o(n_40715) );
in01f80 g739040 ( .a(n_41156), .o(n_41153) );
na02f80 g776837 ( .a(n_3855), .b(n_3863), .o(n_3871) );
no02f80 g741292 ( .a(n_44955), .b(n_38955), .o(n_38995) );
in01f80 newInst_1106 ( .a(newNet_1105), .o(newNet_1106) );
no02f80 g779568 ( .a(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .o(n_1385) );
na02f80 g773852 ( .a(n_7049), .b(n_7048), .o(n_7386) );
no02f80 g749468 ( .a(n_30472), .b(FE_OCP_RBN2633_n_30170), .o(n_30512) );
na02f80 g757545 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_18_), .b(delay_add_ln22_unr14_stage6_stallmux_q_19_), .o(n_22773) );
na02f80 g742369 ( .a(n_37792), .b(n_37241), .o(n_37916) );
in01f80 newInst_1956 ( .a(newNet_1955), .o(newNet_1956) );
in01f80 g768791 ( .a(n_11994), .o(n_11995) );
in01f80 newInst_3456 ( .a(newNet_3455), .o(newNet_3456) );
in01f80 FE_RC_1999_0 ( .a(n_19653), .o(FE_RN_655_0) );
in01f80 newInst_432 ( .a(newNet_288), .o(newNet_432) );
no02f80 g746386 ( .a(n_34779), .b(n_34911), .o(n_35043) );
na02f80 g756929 ( .a(n_23803), .b(n_24023), .o(n_24061) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_16_ ( .ck(newNet_2401), .d(n_36377), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_) );
in01f80 newInst_1016 ( .a(newNet_856), .o(newNet_1016) );
na02f80 g778537 ( .a(n_2817), .b(n_2769), .o(n_3353) );
no02f80 g776217 ( .a(n_4583), .b(n_4592), .o(n_4656) );
na02f80 g760230 ( .a(FE_OCPN1261_n_20242), .b(n_19345), .o(n_20395) );
in01f80 g778681 ( .a(n_2249), .o(n_2230) );
ao12f80 g760562 ( .a(n_20357), .b(n_20356), .c(n_20355), .o(n_21249) );
na02f80 g758148 ( .a(n_21973), .b(FE_OCP_RBN1371_n_20763), .o(n_22046) );
in01f80 g736879 ( .a(n_43601), .o(n_43602) );
na03f80 g743659 ( .a(n_37473), .b(n_37472), .c(n_37306), .o(n_37474) );
no02f80 FE_RC_3692_0 ( .a(n_39249), .b(FE_OCP_RBN2847_n_39479), .o(FE_RN_1624_0) );
in01f80 newInst_1968 ( .a(newNet_1967), .o(newNet_1968) );
in01f80 g744011 ( .a(n_36361), .o(n_36362) );
in01f80 g774327 ( .a(n_6633), .o(n_6634) );
no02f80 g780616 ( .a(n_779), .b(n_859), .o(n_913) );
oa12f80 g777012 ( .a(n_3594), .b(n_3593), .c(n_3592), .o(n_3595) );
in01f80 g762859 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .o(n_17724) );
na02f80 g779215 ( .a(n_1859), .b(n_1858), .o(n_1860) );
na02f80 g744316 ( .a(n_35505), .b(n_35504), .o(n_35519) );
oa22f80 FE_RC_3465_0 ( .a(n_32120), .b(n_32345), .c(n_32121), .d(n_32359), .o(n_32517) );
oa22f80 g753389 ( .a(n_26883), .b(n_26836), .c(n_26828), .d(n_26835), .o(n_26968) );
oa12f80 g742947 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37050), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n_37184) );
ao12f80 g757730 ( .a(n_22212), .b(n_22149), .c(FE_OCP_RBN1851_n_22556), .o(n_22612) );
na02f80 g770806 ( .a(n_10111), .b(n_10107), .o(n_10115) );
in01f80 FE_OCP_RBC3129_n_32266 ( .a(n_32266), .o(FE_OCP_RBN3129_n_32266) );
in01f80 g769039 ( .a(n_11694), .o(n_11695) );
no02f80 g754507 ( .a(n_26707), .b(n_26712), .o(n_26771) );
no02f80 g752231 ( .a(n_27918), .b(n_27919), .o(n_27941) );
in01f80 newInst_2567 ( .a(newNet_1371), .o(newNet_2567) );
no02f80 g776923 ( .a(n_5092), .b(n_5147), .o(n_5148) );
in01f80 g760139 ( .a(n_20667), .o(n_20668) );
in01f80 g743273 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .o(n_36828) );
no02f80 g736921 ( .a(n_43015), .b(n_43014), .o(n_43023) );
oa12f80 g765959 ( .a(n_14897), .b(n_14915), .c(n_14896), .o(n_14999) );
in01f80 g750579 ( .a(FE_OCP_RBN2347_n_29448), .o(n_30310) );
in01f80 FE_OCP_RBC3015_n_31117 ( .a(FE_OCP_RBN3009_n_31117), .o(FE_OCP_RBN3015_n_31117) );
in01f80 g778648 ( .a(n_2422), .o(n_3286) );
oa12f80 g737363 ( .a(n_42511), .b(n_42838), .c(n_42529), .o(n_42847) );
no02f80 g749305 ( .a(n_30659), .b(FE_OCP_RBN3675_FE_RN_1581_0), .o(n_30706) );
na02f80 g745228 ( .a(n_35682), .b(n_35809), .o(n_35770) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_7_ ( .ck(newNet_2338), .d(n_35626), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_) );
in01f80 g774776 ( .a(n_6442), .o(n_6443) );
in01f80 g771184 ( .a(n_9360), .o(n_9361) );
na02f80 g745515 ( .a(n_34486), .b(n_47255), .o(n_34511) );
in01f80 newInst_323 ( .a(newNet_322), .o(newNet_323) );
oa12f80 g774760 ( .a(n_6220), .b(n_45217), .c(n_6173), .o(n_6332) );
in01f80 g741824 ( .a(n_38510), .o(n_38526) );
in01f80 newInst_2337 ( .a(newNet_2336), .o(newNet_2337) );
in01f80 g743761 ( .a(n_36272), .o(n_36309) );
oa12f80 g741761 ( .a(n_38314), .b(n_38425), .c(n_38333), .o(n_38457) );
no02f80 g738862 ( .a(n_41299), .b(n_41320), .o(n_41321) );
na02f80 g759223 ( .a(n_20980), .b(n_20924), .o(n_21012) );
in01f80 g761619 ( .a(n_19609), .o(n_19649) );
no02f80 g776572 ( .a(n_4225), .b(n_4046), .o(n_4321) );
ao12f80 g753419 ( .a(n_26691), .b(n_26765), .c(n_26660), .o(n_26882) );
in01f80 FE_OCP_RBC2945_FE_RN_1269_0 ( .a(FE_RN_1269_0), .o(FE_OCP_RBN2945_FE_RN_1269_0) );
no02f80 g762318 ( .a(n_18077), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .o(n_18091) );
no02f80 g770929 ( .a(n_9581), .b(n_9472), .o(n_9675) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_28_ ( .ck(newNet_2077), .d(n_6670), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_) );
in01f80 FE_OCPC1422_n_35611 ( .a(FE_OCPN1421_n_35611), .o(FE_OCPN1422_n_35611) );
na02f80 g766486 ( .a(n_14024), .b(n_13440), .o(n_14095) );
oa22f80 FE_RC_3212_0 ( .a(n_921), .b(n_44659), .c(n_920), .d(n_44623), .o(n_1340) );
in01f80 g766807 ( .a(n_14489), .o(n_14490) );
ao12f80 g737535 ( .a(n_42509), .b(n_42508), .c(n_42507), .o(n_43052) );
oa12f80 g756306 ( .a(n_24235), .b(n_24587), .c(n_24256), .o(n_24629) );
in01f80 g739470 ( .a(n_40716), .o(n_40717) );
ao12f80 g775460 ( .a(n_4998), .b(n_45323), .c(n_5061), .o(n_5428) );
no02f80 g764822 ( .a(n_15627), .b(n_15592), .o(n_15696) );
na02f80 g741341 ( .a(FE_OCP_RBN3582_n_44944), .b(n_38603), .o(n_39183) );
no02f80 g760245 ( .a(FE_OCP_RBN3617_n_20249), .b(n_20523), .o(n_20565) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_9_ ( .ck(newNet_2695), .d(n_16105), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_) );
in01f80 g775217 ( .a(n_5693), .o(n_5732) );
oa12f80 g763778 ( .a(n_16373), .b(n_16609), .c(n_16232), .o(n_16649) );
in01f80 FE_OCP_RBC3628_n_38870 ( .a(FE_OCP_RBN3627_n_38870), .o(FE_OCP_RBN3628_n_38870) );
oa22f80 g780036 ( .a(n_1245), .b(n_930), .c(n_1246), .d(n_931), .o(n_1257) );
no02f80 g773399 ( .a(n_7562), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .o(n_8531) );
no02f80 g773823 ( .a(n_7180), .b(n_7170), .o(n_7171) );
oa12f80 g743558 ( .a(n_36007), .b(n_36514), .c(n_36035), .o(n_36535) );
in01f80 FE_OCP_RBC2544_n_9082 ( .a(n_9082), .o(FE_OCP_RBN2544_n_9082) );
oa12f80 g744707 ( .a(n_30633), .b(n_35155), .c(n_35029), .o(n_35211) );
in01f80 FE_OCP_RBC3089_FE_OCPN1052_n_31674 ( .a(FE_OCPN1052_n_31674), .o(FE_OCP_RBN3089_FE_OCPN1052_n_31674) );
ao12f80 g779308 ( .a(n_1709), .b(n_1708), .c(n_1707), .o(n_2442) );
ao12f80 g760477 ( .a(n_19887), .b(n_19950), .c(n_19835), .o(n_20033) );
na02f80 g758044 ( .a(n_22645), .b(n_22920), .o(n_22921) );
oa22f80 g739636 ( .a(n_40592), .b(n_40598), .c(n_40583), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40597) );
in01f80 g762358 ( .a(n_18583), .o(n_18532) );
no02f80 FE_RC_1868_0 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .b(FE_OCP_RBN3824_n_44061), .o(FE_RN_575_0) );
in01f80 FE_OCP_RBC3545_n_44575 ( .a(n_44575), .o(FE_OCP_RBN3545_n_44575) );
in01f80 newInst_1790 ( .a(newNet_1789), .o(newNet_1790) );
na02f80 g744520 ( .a(n_35402), .b(n_35414), .o(n_35403) );
no02f80 g740919 ( .a(n_39338), .b(n_39337), .o(n_39339) );
na02f80 g759047 ( .a(n_21163), .b(n_45024), .o(n_21200) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_12_ ( .ck(newNet_2681), .d(n_22044), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_) );
in01f80 newInst_354 ( .a(newNet_353), .o(newNet_354) );
in01f80 g769565 ( .a(n_11398), .o(n_11399) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_11_ ( .ck(newNet_2790), .d(n_16362), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_) );
in01f80 g779544 ( .a(n_1878), .o(n_1879) );
na02f80 g773884 ( .a(n_7061), .b(n_6969), .o(n_7127) );
in01f80 FE_OCP_RBC2391_n_19434 ( .a(FE_OCP_RBN2390_n_19434), .o(FE_OCP_RBN2391_n_19434) );
no02f80 g762351 ( .a(n_45002), .b(n_18252), .o(n_18766) );
in01f80 newInst_2581 ( .a(newNet_2580), .o(newNet_2581) );
in01f80 g755942 ( .a(n_24268), .o(n_24314) );
in01f80 g742116 ( .a(n_38158), .o(n_38159) );
in01f80 g737289 ( .a(n_42912), .o(n_42913) );
in01f80 g760971 ( .a(n_19382), .o(n_19383) );
oa12f80 g736548 ( .a(n_318), .b(n_43650), .c(FE_OFN4_n_43918), .o(n_43685) );
in01f80 g769795 ( .a(n_11307), .o(n_11282) );
in01f80 g759681 ( .a(n_21300), .o(n_21301) );
no02f80 g740382 ( .a(FE_OCP_RBN3028_n_39942), .b(n_39891), .o(n_40246) );
oa12f80 g772281 ( .a(n_7530), .b(n_8504), .c(n_7511), .o(n_8621) );
na02f80 g779635 ( .a(n_1463), .b(n_1462), .o(n_1817) );
in01f80 g775420 ( .a(n_5876), .o(n_5807) );
in01f80 g738667 ( .a(n_41779), .o(n_41780) );
in01f80 newInst_1332 ( .a(newNet_43), .o(newNet_1332) );
na02f80 g775235 ( .a(n_5691), .b(n_5667), .o(n_5782) );
no02f80 g760639 ( .a(n_19726), .b(FE_OCP_RBN3832_n_19204), .o(n_19755) );
in01f80 newInst_3194 ( .a(newNet_3193), .o(newNet_3194) );
na02f80 g760510 ( .a(n_19999), .b(n_20007), .o(n_20000) );
no02f80 g765828 ( .a(n_14872), .b(FE_OCP_RBN2504_n_13896), .o(n_14956) );
na02f80 g760109 ( .a(n_20340), .b(FE_OCP_RBN1342_n_19077), .o(n_20374) );
na02f80 g778151 ( .a(n_2885), .b(n_2813), .o(n_2940) );
ao12f80 g756834 ( .a(n_24354), .b(n_24150), .c(n_24059), .o(n_24903) );
oa12f80 g767657 ( .a(n_13317), .b(n_13377), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n_13422) );
na02f80 g768425 ( .a(n_12391), .b(n_12420), .o(n_12447) );
na02f80 g736858 ( .a(n_43324), .b(n_43456), .o(n_43543) );
in01f80 FE_OCP_RBC3691_n_10567 ( .a(n_10567), .o(FE_OCP_RBN3691_n_10567) );
na02f80 g772724 ( .a(n_8187), .b(n_7817), .o(n_8202) );
in01f80 FE_OCPC1855_n_33341 ( .a(n_33341), .o(FE_OCPN1855_n_33341) );
in01f80 g768132 ( .a(n_12645), .o(n_12646) );
oa22f80 FE_RC_2920_0 ( .a(n_12902), .b(FE_OCP_RBN3421_n_12879), .c(n_12879), .d(FE_OCP_RBN2224_n_12902), .o(n_13050) );
in01f80 g738679 ( .a(n_41604), .o(n_41901) );
in01f80 FE_OCP_DRV_C1550_n_19053 ( .a(FE_OCP_DRV_N1549_n_19053), .o(FE_OCP_DRV_N1550_n_19053) );
no02f80 g750310 ( .a(n_29720), .b(n_29706), .o(n_29707) );
na02f80 g748916 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .o(n_32407) );
oa22f80 g740031 ( .a(n_39899), .b(n_39829), .c(n_39898), .d(n_39830), .o(n_39986) );
na02f80 g765979 ( .a(n_14672), .b(n_13404), .o(n_14754) );
in01f80 g772203 ( .a(n_8857), .o(n_8895) );
no02f80 g740770 ( .a(n_39295), .b(n_39193), .o(n_39386) );
in01f80 g753917 ( .a(n_26358), .o(n_26433) );
in01f80 newInst_416 ( .a(newNet_415), .o(newNet_416) );
ao22s80 g765409 ( .a(n_16245), .b(n_14081), .c(n_15874), .d(n_14044), .o(n_16344) );
no02f80 g751478 ( .a(n_28627), .b(n_28626), .o(n_28643) );
no02f80 g751354 ( .a(n_28771), .b(n_28648), .o(n_28805) );
na02f80 g771671 ( .a(n_10073), .b(n_44516), .o(n_11266) );
ao22s80 FE_RC_1155_0 ( .a(n_7802), .b(FE_OCP_RBN2406_n_8242), .c(FE_OCP_RBN3455_FE_OCPN1240_n_7721), .d(n_8242), .o(n_8335) );
in01f80 FE_RC_2349_0 ( .a(n_1645), .o(FE_RN_902_0) );
no02f80 g766013 ( .a(n_14614), .b(n_14317), .o(n_14668) );
na02f80 g740656 ( .a(n_39598), .b(n_45841), .o(n_39618) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_12_ ( .ck(newNet_981), .d(n_22963), .o(delay_xor_ln21_unr15_stage6_stallmux_q_12_) );
in01f80 newInst_119 ( .a(newNet_118), .o(newNet_119) );
na02f80 g770070 ( .a(n_10791), .b(n_10792), .o(n_10883) );
in01f80 FE_OFC815_n_19807 ( .a(FE_OFN831_n_19807), .o(FE_OFN815_n_19807) );
ao12f80 g746496 ( .a(FE_OCP_DRV_N3148_n_33225), .b(n_33207), .c(n_32923), .o(n_33273) );
no02f80 g769059 ( .a(FE_OCP_RBN3268_n_45224), .b(n_11558), .o(n_11690) );
in01f80 g764861 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n_16503) );
no02f80 g776551 ( .a(n_4243), .b(FE_OCP_RBN2625_n_3848), .o(n_4309) );
in01f80 g761946 ( .a(n_18318), .o(n_18360) );
no02f80 g751588 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .o(n_28568) );
in01f80 newInst_349 ( .a(newNet_34), .o(newNet_349) );
no02f80 g750650 ( .a(n_29414), .b(n_29465), .o(n_29514) );
ao12f80 g773016 ( .a(FE_OCP_RBN3460_n_7886), .b(n_8110), .c(n_8062), .o(n_8151) );
oa12f80 g784663 ( .a(n_6349), .b(n_6332), .c(n_6215), .o(n_46993) );
in01f80 g763339 ( .a(n_17378), .o(n_17379) );
in01f80 FE_OCP_RBC2946_n_5428 ( .a(n_5428), .o(FE_OCP_RBN2946_n_5428) );
in01f80 newInst_1396 ( .a(newNet_1395), .o(newNet_1396) );
oa22f80 FE_RC_891_0 ( .a(n_45010), .b(n_20984), .c(n_45070), .d(n_20985), .o(n_21127) );
in01f80 g761450 ( .a(n_20084), .o(n_20085) );
in01f80 g747938 ( .a(n_33238), .o(n_33315) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_18_ ( .ck(newNet_1859), .d(n_16847), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_) );
in01f80 FE_OCP_RBC1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
oa22f80 g744941 ( .a(n_36386), .b(n_36168), .c(n_36356), .d(n_36167), .o(n_36418) );
na02f80 FE_RC_2323_0 ( .a(n_179), .b(n_28811), .o(FE_RN_884_0) );
no02f80 g771219 ( .a(n_9639), .b(n_9446), .o(n_9703) );
oa12f80 g780088 ( .a(n_742), .b(n_1184), .c(n_781), .o(n_1198) );
na02f80 g755462 ( .a(n_24625), .b(n_24604), .o(n_24765) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_31_ ( .ck(newNet_1581), .d(n_27678), .o(n_27923) );
no02f80 g767373 ( .a(n_13399), .b(n_12437), .o(n_13507) );
in01f80 g771182 ( .a(n_9496), .o(n_9510) );
no02f80 g744733 ( .a(n_35154), .b(n_30614), .o(n_35213) );
ao12f80 g781153 ( .a(n_112), .b(n_199), .c(n_130), .o(n_206) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_25_ ( .ck(newNet_3132), .d(n_40560), .o(delay_add_ln22_unr27_stage10_stallmux_q_25_) );
in01f80 g771973 ( .a(n_9951), .o(n_9952) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_8_ ( .ck(newNet_1357), .d(n_36418), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_) );
in01f80 g771905 ( .a(FE_OCP_RBN2468_n_8767), .o(n_10183) );
na02f80 g755128 ( .a(n_25373), .b(n_24450), .o(n_25476) );
na02f80 g776681 ( .a(n_4130), .b(n_4068), .o(n_4360) );
na02f80 g776080 ( .a(n_5048), .b(FE_OCP_RBN2659_n_4101), .o(n_5061) );
no02f80 FE_RC_3698_0 ( .a(FE_RN_1625_0), .b(FE_OCP_RBN3207_n_44365), .o(FE_RN_1627_0) );
no02f80 g742912 ( .a(n_36972), .b(n_36968), .o(n_37339) );
na02f80 g739060 ( .a(n_41151), .b(n_41150), .o(n_41152) );
in01f80 newInst_271 ( .a(newNet_270), .o(newNet_271) );
in01f80 g775563 ( .a(n_5641), .o(n_5642) );
oa12f80 g780526 ( .a(n_976), .b(n_890), .c(n_906), .o(n_1072) );
ao12f80 g759737 ( .a(n_20168), .b(n_20251), .c(n_20224), .o(n_20321) );
na02f80 g776255 ( .a(n_4950), .b(n_4932), .o(n_5207) );
na02f80 g764795 ( .a(n_15890), .b(n_15889), .o(n_15891) );
in01f80 g776505 ( .a(n_4532), .o(n_4533) );
oa12f80 g738285 ( .a(n_41800), .b(n_41799), .c(n_41798), .o(n_41867) );
in01f80 newInst_2081 ( .a(newNet_2080), .o(newNet_2081) );
na02f80 g768765 ( .a(n_11921), .b(n_11848), .o(n_12027) );
no02f80 g761191 ( .a(n_20050), .b(n_20009), .o(n_21019) );
in01f80 g739406 ( .a(n_40728), .o(n_40729) );
in01f80 g737210 ( .a(n_42992), .o(n_42993) );
na02f80 FE_RC_2236_0 ( .a(FE_RN_814_0), .b(FE_RN_815_0), .o(FE_RN_816_0) );
in01f80 g752852 ( .a(n_28021), .o(n_28022) );
in01f80 FE_RC_4215_0 ( .a(n_14988), .o(FE_RN_1845_0) );
in01f80 g772360 ( .a(n_8714), .o(n_8715) );
na02f80 g775407 ( .a(n_5469), .b(FE_OCP_RBN2733_n_4219), .o(n_5537) );
na02f80 g767369 ( .a(n_13389), .b(n_13386), .o(n_13496) );
no02f80 g765132 ( .a(FE_OCP_RBN2693_n_15083), .b(n_14758), .o(n_15162) );
ao12f80 g756354 ( .a(n_23798), .b(n_23827), .c(n_23797), .o(n_23892) );
in01f80 g756930 ( .a(n_23950), .o(n_23951) );
no02f80 g755299 ( .a(n_24939), .b(n_24938), .o(n_24940) );
in01f80 g763460 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_3_), .o(n_16881) );
no02f80 g754707 ( .a(n_26160), .b(n_25441), .o(n_26308) );
na02f80 g778952 ( .a(n_2158), .b(n_1969), .o(n_2159) );
no02f80 g751049 ( .a(n_30290), .b(n_30256), .o(n_30334) );
in01f80 FE_OCP_RBC2594_n_25181 ( .a(FE_OCP_RBN2592_n_25181), .o(FE_OCP_RBN2594_n_25181) );
no02f80 g775821 ( .a(n_5030), .b(n_5051), .o(n_5071) );
oa22f80 g762720 ( .a(n_17632), .b(n_17539), .c(n_18197), .d(n_17358), .o(n_18256) );
no02f80 g746544 ( .a(n_34608), .b(n_34544), .o(n_35126) );
in01f80 FE_OCP_DRV_C3149_n_12773 ( .a(n_12773), .o(FE_OCP_DRV_N3149_n_12773) );
in01f80 g743679 ( .a(n_36349), .o(n_36350) );
in01f80 g738342 ( .a(n_41755), .o(n_41756) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_15_ ( .ck(newNet_2780), .d(n_16757), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_) );
na02f80 g776067 ( .a(n_4940), .b(n_4994), .o(n_5095) );
in01f80 g742004 ( .a(n_38239), .o(n_38240) );
in01f80 newInst_85 ( .a(newNet_39), .o(newNet_85) );
ao12f80 g767294 ( .a(n_13080), .b(n_13678), .c(n_13115), .o(n_13718) );
na02f80 g749258 ( .a(n_30824), .b(n_30708), .o(n_30822) );
na02f80 g741270 ( .a(FE_OCP_RBN2546_n_44944), .b(n_39025), .o(n_39068) );
ao22s80 g784431 ( .a(n_36713), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .o(n_46243) );
na02f80 g769244 ( .a(n_11440), .b(n_11435), .o(n_11658) );
in01f80 FE_OCP_RBC1189_n_14911 ( .a(n_14911), .o(FE_OCP_RBN1189_n_14911) );
na02f80 g751156 ( .a(n_29800), .b(n_29799), .o(n_29821) );
in01f80 g741581 ( .a(n_38683), .o(n_38684) );
no02f80 g750596 ( .a(n_29395), .b(n_25738), .o(n_29446) );
oa22f80 FE_RC_3378_0 ( .a(n_45066), .b(n_20509), .c(n_45101), .d(n_20510), .o(n_20650) );
no02f80 g773095 ( .a(n_7721), .b(n_8676), .o(n_7722) );
in01f80 g746267 ( .a(n_47249), .o(n_33620) );
no02f80 g775050 ( .a(n_6020), .b(n_5740), .o(n_6082) );
in01f80 FE_RC_3729_0 ( .a(n_19565), .o(FE_RN_1641_0) );
ao12f80 g766280 ( .a(n_14121), .b(n_14286), .c(n_14240), .o(n_14287) );
no02f80 FE_RC_602_0 ( .a(n_40626), .b(n_40664), .o(FE_RN_190_0) );
no02f80 g766589 ( .a(n_13885), .b(n_13363), .o(n_13953) );
in01f80 g747314 ( .a(n_33910), .o(n_33911) );
in01f80 FE_OCP_RBC3647_n_44490 ( .a(FE_OCP_RBN3642_n_44490), .o(FE_OCP_RBN3647_n_44490) );
na02f80 g739293 ( .a(n_40729), .b(n_40820), .o(n_40846) );
in01f80 newInst_592 ( .a(newNet_591), .o(newNet_592) );
na02f80 g774957 ( .a(n_6000), .b(n_6064), .o(n_6084) );
na02f80 g751822 ( .a(n_28249), .b(n_28089), .o(n_28267) );
in01f80 g743902 ( .a(n_35627), .o(n_35671) );
in01f80 g766157 ( .a(n_14552), .o(n_14553) );
na02f80 g754752 ( .a(n_25383), .b(n_25490), .o(n_25512) );
in01f80 g737514 ( .a(n_46943), .o(n_43158) );
oa12f80 g752314 ( .a(n_28446), .b(n_28457), .c(n_28445), .o(n_28937) );
in01f80 FE_OCP_RBC1133_n_16041 ( .a(n_16041), .o(FE_OCP_RBN1133_n_16041) );
oa12f80 g778256 ( .a(n_2588), .b(n_2615), .c(n_2587), .o(n_3006) );
ao12f80 g773845 ( .a(n_7080), .b(n_7088), .c(n_7079), .o(n_8016) );
oa12f80 g742442 ( .a(n_37624), .b(n_37646), .c(n_37645), .o(n_37668) );
na02f80 g781052 ( .a(cos_out_28), .b(FE_OFN1_n_43918), .o(n_316) );
no02f80 g768929 ( .a(n_11646), .b(n_11560), .o(n_11776) );
no02f80 FE_RC_4205_0 ( .a(n_18117), .b(n_19561), .o(n_19736) );
no02f80 g763428 ( .a(n_16903), .b(n_16867), .o(n_16920) );
in01f80 fopt783248 ( .a(n_44812), .o(n_44811) );
in01f80 FE_RC_636_0 ( .a(n_6539), .o(FE_RN_199_0) );
in01f80 g754936 ( .a(n_25506), .o(n_25540) );
no02f80 g737597 ( .a(n_42589), .b(n_42474), .o(n_42631) );
no02f80 g773869 ( .a(n_7052), .b(n_7042), .o(n_7043) );
na02f80 g773162 ( .a(n_7817), .b(n_7885), .o(n_8045) );
no02f80 g781246 ( .a(n_43), .b(n_109), .o(n_217) );
in01f80 g738736 ( .a(n_41530), .o(n_41616) );
in01f80 newInst_995 ( .a(newNet_57), .o(newNet_995) );
no02f80 g757399 ( .a(FE_OCP_RBN3821_n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .o(n_23078) );
in01f80 g771929 ( .a(n_9110), .o(n_9061) );
in01f80 g741487 ( .a(n_38750), .o(n_38751) );
in01f80 newInst_1179 ( .a(newNet_1178), .o(newNet_1179) );
na02f80 g767001 ( .a(n_13497), .b(n_12914), .o(n_13534) );
oa22f80 g743634 ( .a(n_36347), .b(n_36259), .c(n_36348), .d(n_36258), .o(n_36415) );
na02f80 g745128 ( .a(n_34632), .b(n_34342), .o(n_34714) );
in01f80 g749328 ( .a(n_30733), .o(n_30759) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_0_ ( .ck(newNet_3660), .d(n_14740), .o(delay_add_ln22_unr11_stage5_stallmux_q_0_) );
in01f80 FE_OCP_RBC2497_n_8835 ( .a(n_8835), .o(FE_OCP_RBN2497_n_8835) );
no03m80 FE_RC_1072_0 ( .a(FE_RN_317_0), .b(n_12333), .c(n_12055), .o(n_12361) );
in01f80 g772233 ( .a(n_8678), .o(n_8679) );
oa12f80 g769625 ( .a(n_11249), .b(n_11294), .c(n_11131), .o(n_11349) );
oa22f80 g758601 ( .a(n_22485), .b(n_21855), .c(n_22486), .d(n_21856), .o(n_22567) );
oa12f80 g770105 ( .a(n_10634), .b(n_10821), .c(n_10678), .o(n_10874) );
no02f80 g779043 ( .a(n_45716), .b(n_1512), .o(n_2074) );
no02f80 g749726 ( .a(n_31311), .b(n_31410), .o(n_31414) );
in01f80 g761889 ( .a(n_18707), .o(n_18708) );
in01f80 g737293 ( .a(n_42886), .o(n_42887) );
in01f80 g761028 ( .a(n_19318), .o(n_19319) );
na02f80 g754320 ( .a(n_25817), .b(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .o(n_25856) );
no03m80 g737560 ( .a(n_42470), .b(n_42420), .c(n_42469), .o(n_42471) );
in01f80 g774582 ( .a(n_6556), .o(n_6586) );
oa12f80 g752595 ( .a(n_27439), .b(n_27568), .c(n_27146), .o(n_27632) );
na02f80 g756192 ( .a(n_24058), .b(n_23707), .o(n_24147) );
in01f80 newInst_2308 ( .a(newNet_2307), .o(newNet_2308) );
no02f80 g742077 ( .a(FE_OCP_RBN3445_n_37945), .b(n_37618), .o(n_38313) );
in01f80 g755277 ( .a(n_25095), .o(n_25096) );
na02f80 g751878 ( .a(n_28905), .b(n_28904), .o(n_28906) );
na02f80 g750845 ( .a(n_29019), .b(n_28700), .o(n_29064) );
ao12f80 g768437 ( .a(n_12400), .b(n_45659), .c(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .o(n_12631) );
oa12f80 g762121 ( .a(n_18668), .b(n_18703), .c(n_18667), .o(n_18777) );
no02f80 g749884 ( .a(n_29841), .b(n_29926), .o(n_29988) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_3_ ( .ck(newNet_302), .d(n_1360), .o(delay_xor_ln22_unr3_stage2_stallmux_q_3_) );
no02f80 g757204 ( .a(n_23225), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_), .o(n_23245) );
ao22s80 FE_RC_740_0 ( .a(n_7541), .b(n_8547), .c(n_8546), .d(n_7540), .o(n_8664) );
oa22f80 FE_RC_394_0 ( .a(n_12997), .b(n_13533), .c(n_12998), .d(n_13532), .o(n_13616) );
oa12f80 g775634 ( .a(n_5116), .b(n_5455), .c(n_5203), .o(n_5551) );
in01f80 g775388 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_12_), .o(n_5777) );
oa12f80 g742016 ( .a(n_37955), .b(FE_OCP_RBN3445_n_37945), .c(n_37894), .o(n_38365) );
in01f80 newInst_705 ( .a(newNet_102), .o(newNet_705) );
in01f80 g767445 ( .a(n_13266), .o(n_13267) );
in01f80 g765328 ( .a(n_15113), .o(n_15114) );
in01f80 g763723 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .o(n_17212) );
no02f80 g768093 ( .a(n_12914), .b(n_12887), .o(n_13210) );
in01f80 g758263 ( .a(n_22645), .o(n_22730) );
no02f80 g761549 ( .a(n_18938), .b(FE_OCP_DRV_N1548_n_17643), .o(n_18996) );
no02f80 g742811 ( .a(n_37297), .b(n_37028), .o(n_37331) );
no02f80 g758895 ( .a(n_21433), .b(n_21428), .o(n_21500) );
na02f80 g778448 ( .a(n_2419), .b(n_2371), .o(n_2453) );
in01f80 g737206 ( .a(n_42973), .o(n_42974) );
no02f80 g747802 ( .a(n_33208), .b(n_32585), .o(n_33258) );
in01f80 newInst_765 ( .a(newNet_764), .o(newNet_765) );
ao12f80 FE_RC_4029_0 ( .a(FE_RN_1750_0), .b(n_14419), .c(n_15900), .o(n_16074) );
in01f80 g756620 ( .a(n_23815), .o(n_23816) );
in01f80 FE_OCPC942_n_44925 ( .a(FE_OCPN941_n_44925), .o(FE_OCPN942_n_44925) );
in01f80 g767838 ( .a(n_12800), .o(n_14003) );
no02f80 g741017 ( .a(n_38863), .b(FE_OCP_RBN2635_n_38806), .o(n_38933) );
in01f80 fopt783138 ( .a(n_44636), .o(n_44623) );
na02f80 g780772 ( .a(n_471), .b(n_456), .o(n_490) );
in01f80 FE_RC_2586_0 ( .a(FE_RN_1069_0), .o(n_17954) );
in01f80 g760929 ( .a(n_19333), .o(n_19334) );
ao12f80 g773776 ( .a(n_6753), .b(n_7206), .c(n_6705), .o(n_7264) );
no02f80 g742967 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_26_), .o(n_37471) );
in01f80 g751145 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30545) );
in01f80 FE_OCPC3781_n_16440 ( .a(FE_OCPN3780_n_16440), .o(FE_OCPN3781_n_16440) );
oa22f80 FE_RC_538_0 ( .a(n_29348), .b(n_28821), .c(n_28820), .d(n_29347), .o(n_29448) );
no02f80 g736651 ( .a(n_43374), .b(n_43233), .o(n_43442) );
in01f80 newInst_2601 ( .a(newNet_2600), .o(newNet_2601) );
no02f80 g770759 ( .a(n_10212), .b(n_10067), .o(n_10256) );
oa22f80 g768622 ( .a(n_12204), .b(n_12225), .c(n_12205), .d(n_12292), .o(n_13264) );
in01f80 g765670 ( .a(n_15132), .o(n_15133) );
in01f80 newInst_208 ( .a(newNet_206), .o(newNet_208) );
ao12f80 g757520 ( .a(n_22196), .b(FE_OCP_RBN1849_n_22639), .c(n_22129), .o(n_22756) );
in01f80 newInst_895 ( .a(newNet_460), .o(newNet_895) );
ao12f80 g771033 ( .a(n_9787), .b(n_9822), .c(n_9698), .o(n_10049) );
in01f80 g777692 ( .a(n_3468), .o(n_3469) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_9_ ( .ck(newNet_870), .d(n_32373), .o(delay_xor_ln21_unr21_stage8_stallmux_q_9_) );
na02f80 g743361 ( .a(n_36593), .b(n_36617), .o(n_36673) );
no02f80 g775278 ( .a(n_5808), .b(n_5743), .o(n_5778) );
na02f80 g754902 ( .a(FE_OCP_RBN2597_n_25181), .b(FE_OCP_RBN2280_n_24199), .o(n_25399) );
in01f80 g758740 ( .a(n_22286), .o(n_22287) );
oa22f80 g779893 ( .a(n_44652), .b(n_1189), .c(n_44637), .d(n_1179), .o(n_1334) );
na02f80 g746455 ( .a(n_35017), .b(n_35016), .o(n_35018) );
in01f80 g746217 ( .a(n_35045), .o(n_35089) );
na02f80 g741600 ( .a(n_38616), .b(n_38778), .o(n_38652) );
no02f80 g775255 ( .a(n_5836), .b(n_5773), .o(n_5856) );
in01f80 g752941 ( .a(n_27876), .o(n_27877) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_21_ ( .ck(newNet_816), .d(n_1302), .o(delay_xor_ln21_unr3_stage2_stallmux_q_21_) );
no02f80 g749018 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .o(n_32312) );
no02f80 g762113 ( .a(n_18242), .b(n_17568), .o(n_18309) );
in01f80 newInst_2994 ( .a(newNet_2993), .o(newNet_2994) );
in01f80 newInst_367 ( .a(newNet_108), .o(newNet_367) );
ao22s80 FE_RC_772_0 ( .a(n_10150), .b(n_10195), .c(n_10149), .d(n_10196), .o(n_10369) );
na02f80 g763504 ( .a(FE_OCP_RBN3081_n_16977), .b(n_15651), .o(n_17171) );
oa12f80 g738818 ( .a(n_41333), .b(n_41356), .c(n_41332), .o(n_41386) );
in01f80 g760899 ( .a(n_19462), .o(n_19463) );
na02f80 g756348 ( .a(n_24453), .b(n_23988), .o(n_24480) );
na02f80 g756055 ( .a(n_24270), .b(n_24249), .o(n_24250) );
na02f80 g755348 ( .a(n_24964), .b(n_22484), .o(n_24965) );
in01f80 g747076 ( .a(n_33034), .o(n_33108) );
na02f80 FE_RC_4199_0 ( .a(n_19184), .b(n_18458), .o(n_19250) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_30_ ( .ck(newNet_1193), .d(n_6405), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_) );
no02f80 g771591 ( .a(n_8870), .b(FE_OCP_RBN3475_n_7886), .o(n_8913) );
in01f80 g743092 ( .a(n_36988), .o(n_37096) );
na02f80 g739890 ( .a(n_40379), .b(n_40068), .o(n_40400) );
in01f80 fopt783062 ( .a(n_44463), .o(n_44464) );
in01f80 g750733 ( .a(n_30337), .o(n_30338) );
no02f80 g775865 ( .a(n_5014), .b(n_5051), .o(n_5142) );
na02f80 g739652 ( .a(n_40547), .b(n_40556), .o(n_40578) );
oa12f80 g736578 ( .a(n_304), .b(n_43648), .c(FE_OFN5_n_43918), .o(n_43680) );
in01f80 g743504 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .o(n_36537) );
na02f80 g763812 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .o(n_17532) );
in01f80 g738442 ( .a(n_41766), .o(n_41767) );
no02f80 g749974 ( .a(n_30173), .b(n_30194), .o(n_30259) );
no02f80 FE_RC_4077_0 ( .a(n_16837), .b(n_16759), .o(FE_RN_1777_0) );
na02f80 g765551 ( .a(n_15142), .b(n_14191), .o(n_15143) );
no02f80 g742315 ( .a(n_37831), .b(n_37816), .o(n_37950) );
in01f80 FE_OCPC1456_n_18860 ( .a(FE_OCPN1455_n_18860), .o(FE_OCPN1456_n_18860) );
in01f80 newInst_3681 ( .a(newNet_3680), .o(newNet_3681) );
in01f80 g737734 ( .a(n_42434), .o(n_42435) );
no02f80 g775862 ( .a(n_5200), .b(n_5087), .o(n_5230) );
in01f80 FE_OCP_RBC2293_n_2438 ( .a(FE_OCP_RBN2290_n_2438), .o(FE_OCP_RBN2293_n_2438) );
in01f80 newInst_2429 ( .a(newNet_2428), .o(newNet_2429) );
in01f80 g766712 ( .a(FE_OCP_RBN1170_n_13756), .o(n_13833) );
no02f80 g754869 ( .a(n_25328), .b(n_25329), .o(n_25396) );
in01f80 newInst_3588 ( .a(newNet_3154), .o(newNet_3588) );
oa12f80 g775324 ( .a(n_5861), .b(n_5860), .c(n_5859), .o(n_5915) );
in01f80 FE_OCP_RBC2170_n_32892 ( .a(FE_OCP_RBN2167_n_32892), .o(FE_OCP_RBN2170_n_32892) );
no02f80 g754805 ( .a(n_26106), .b(n_26072), .o(n_26073) );
in01f80 FE_OCPC3172_n_34222 ( .a(FE_OCPN3171_n_34222), .o(FE_OCPN3172_n_34222) );
in01f80 g775001 ( .a(n_6153), .o(n_6220) );
oa12f80 g773119 ( .a(n_7917), .b(n_8362), .c(n_7923), .o(n_8724) );
in01f80 g763272 ( .a(FE_OCPN1454_n_18559), .o(n_18748) );
no02f80 g741231 ( .a(n_39069), .b(n_39094), .o(n_39176) );
in01f80 FE_RC_3402_0 ( .a(FE_RN_617_0), .o(FE_RN_1472_0) );
in01f80 newInst_302 ( .a(newNet_301), .o(newNet_302) );
oa12f80 g739732 ( .a(n_40229), .b(n_40466), .c(n_40119), .o(n_40491) );
in01f80 g741404 ( .a(n_38868), .o(n_38869) );
in01f80 fopt783533 ( .a(n_45144), .o(n_45146) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_0_ ( .ck(newNet_2501), .d(n_30813), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_) );
in01f80 g746235 ( .a(n_33752), .o(n_33769) );
na02f80 g736392 ( .a(n_43801), .b(n_43658), .o(n_43848) );
in01f80 newInst_3047 ( .a(newNet_1863), .o(newNet_3047) );
oa12f80 g767998 ( .a(n_12704), .b(n_12703), .c(n_12702), .o(n_12990) );
no02f80 g752937 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_), .o(n_27929) );
in01f80 g768452 ( .a(n_12396), .o(n_12397) );
in01f80 FE_OCP_RBC2145_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2143_FE_OCPN861_n_45450), .o(FE_OCP_RBN2145_FE_OCPN861_n_45450) );
na02f80 g781041 ( .a(sin_out_26), .b(FE_OFN4_n_43918), .o(n_302) );
in01f80 g775290 ( .a(n_5667), .o(n_5714) );
na02f80 g761621 ( .a(n_19495), .b(n_19406), .o(n_19609) );
in01f80 g780560 ( .a(n_869), .o(n_844) );
in01f80 g744994 ( .a(n_34880), .o(n_34881) );
in01f80 FE_OCP_RBC2235_n_29055 ( .a(n_29055), .o(FE_OCP_RBN2235_n_29055) );
no02f80 g779342 ( .a(FE_OCP_RBN2156_n_1602), .b(n_1385), .o(n_1675) );
in01f80 g743957 ( .a(n_36318), .o(n_36319) );
na02f80 g781306 ( .a(n_1), .b(n_51), .o(n_59) );
ao12f80 g750267 ( .a(n_30894), .b(n_30893), .c(n_30892), .o(n_31213) );
oa12f80 g779799 ( .a(n_2115), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .o(n_2137) );
in01f80 FE_OFC840_n_3500 ( .a(n_3500), .o(FE_OFN840_n_3500) );
in01f80 newInst_807 ( .a(newNet_806), .o(newNet_807) );
na02f80 g739371 ( .a(n_40917), .b(n_40928), .o(n_40949) );
no02f80 g750104 ( .a(FE_OCP_RBN3566_n_29857), .b(FE_OCP_RBN1153_n_29053), .o(n_30356) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_15_ ( .ck(newNet_658), .d(n_46355), .o(delay_xor_ln21_unr9_stage4_stallmux_q_15_) );
in01f80 g779678 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .o(n_1374) );
no02f80 g772921 ( .a(n_7953), .b(n_7849), .o(n_8028) );
in01f80 g758723 ( .a(n_21910), .o(n_21911) );
in01f80 g755025 ( .a(FE_OCP_RBN2594_n_25181), .o(n_25210) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_15_ ( .ck(newNet_1868), .d(n_16744), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_) );
na02f80 g749129 ( .a(n_30871), .b(n_27130), .o(n_30912) );
no02f80 g741313 ( .a(n_38830), .b(n_38468), .o(n_38852) );
in01f80 FE_RC_3310_0 ( .a(n_13833), .o(FE_RN_1456_0) );
no02f80 g767675 ( .a(n_13281), .b(n_13278), .o(n_13351) );
na02f80 g742827 ( .a(n_37230), .b(n_37129), .o(n_37231) );
no02f80 g742708 ( .a(n_37379), .b(n_37017), .o(n_37371) );
in01f80 g774357 ( .a(n_6868), .o(n_6869) );
no02f80 g778542 ( .a(n_2335), .b(n_2237), .o(n_2336) );
in01f80 newInst_3565 ( .a(newNet_3564), .o(newNet_3565) );
in01f80 g763712 ( .a(n_16736), .o(n_16737) );
in01f80 newInst_1942 ( .a(newNet_857), .o(newNet_1942) );
in01f80 FE_RC_4048_0 ( .a(n_36075), .o(FE_RN_1759_0) );
in01f80 g778964 ( .a(n_2140), .o(n_2611) );
in01f80 g762427 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_17_), .o(n_18009) );
in01f80 FE_OCP_RBC2278_n_24173 ( .a(n_24173), .o(FE_OCP_RBN2278_n_24173) );
no02f80 g777351 ( .a(n_3938), .b(n_3911), .o(n_3990) );
in01f80 g762863 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n_17748) );
na02f80 g776474 ( .a(n_4392), .b(n_4317), .o(n_4511) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_26_ ( .ck(newNet_3035), .d(n_1211), .o(delay_add_ln22_unr2_stage2_stallmux_q_26_) );
na02f80 g776363 ( .a(n_4579), .b(n_4659), .o(n_4714) );
in01f80 newInst_2416 ( .a(newNet_2415), .o(newNet_2416) );
no02f80 g761143 ( .a(n_19798), .b(n_19913), .o(n_19853) );
na02f80 g775010 ( .a(n_6082), .b(n_5845), .o(n_6152) );
oa22f80 FE_RC_3225_0 ( .a(n_18032), .b(n_19353), .c(n_19218), .d(FE_OCP_RBN1698_n_19353), .o(n_19462) );
ao12f80 g754816 ( .a(n_25245), .b(n_25282), .c(n_25244), .o(n_26956) );
in01f80 fopt784015 ( .a(n_11914), .o(n_45748) );
in01f80 FE_RC_2589_0 ( .a(n_12107), .o(FE_RN_1071_0) );
oa22f80 FE_RC_329_0 ( .a(n_22496), .b(n_22744), .c(n_22497), .d(n_22706), .o(n_22902) );
ao22s80 g736561 ( .a(n_43628), .b(n_43594), .c(n_43627), .d(n_43593), .o(n_43660) );
oa12f80 g775101 ( .a(n_5247), .b(n_6062), .c(n_5111), .o(n_6076) );
in01f80 g767571 ( .a(n_12981), .o(n_13010) );
no02f80 g771385 ( .a(n_9370), .b(FE_OCP_RBN3572_n_44563), .o(n_9446) );
in01f80 g761739 ( .a(n_18713), .o(n_18746) );
na02f80 g753309 ( .a(n_27167), .b(n_26247), .o(n_27291) );
na02f80 g753089 ( .a(n_27231), .b(n_27230), .o(n_27267) );
in01f80 g751602 ( .a(n_28773), .o(n_28800) );
na02f80 g756703 ( .a(n_23483), .b(n_23111), .o(n_23563) );
na02f80 g746033 ( .a(n_33959), .b(n_33958), .o(n_33978) );
ao12f80 g740674 ( .a(n_39485), .b(n_39484), .c(n_39483), .o(n_39543) );
no02f80 g771704 ( .a(n_9236), .b(n_9105), .o(n_9284) );
no02f80 g740756 ( .a(n_39385), .b(n_39077), .o(n_39443) );
oa12f80 g740013 ( .a(n_39771), .b(n_39824), .c(n_39751), .o(n_39849) );
in01f80 g764997 ( .a(n_15537), .o(n_15538) );
no02f80 g775987 ( .a(n_4800), .b(n_4669), .o(n_4844) );
in01f80 g773184 ( .a(n_45825), .o(n_7644) );
no02f80 g776330 ( .a(n_4809), .b(n_3717), .o(n_4931) );
in01f80 FE_OCPC894_n_6521 ( .a(n_6521), .o(FE_OCPN894_n_6521) );
na02f80 g758798 ( .a(n_21586), .b(n_45073), .o(n_21616) );
oa12f80 g767363 ( .a(n_13621), .b(n_13620), .c(n_13150), .o(n_13652) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_5_ ( .ck(newNet_617), .d(n_46377), .o(delay_xor_ln21_unr9_stage4_stallmux_q_5_) );
oa22f80 FE_RC_3872_0 ( .a(n_28604), .b(n_28969), .c(n_28603), .d(n_28968), .o(n_29056) );
na02f80 g774494 ( .a(n_6556), .b(n_5984), .o(n_6887) );
in01f80 g764298 ( .a(n_47268), .o(n_16293) );
na02f80 g772034 ( .a(n_8793), .b(n_8686), .o(n_8825) );
na02f80 g753784 ( .a(n_26467), .b(n_26372), .o(n_26493) );
in01f80 newInst_982 ( .a(newNet_879), .o(newNet_982) );
ao12f80 g768988 ( .a(n_11694), .b(FE_OCP_RBN2117_n_45224), .c(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .o(n_12038) );
na02f80 g764248 ( .a(n_16377), .b(n_16441), .o(n_16464) );
na02f80 g748814 ( .a(n_32448), .b(n_32555), .o(n_33115) );
in01f80 FE_OCP_RBC1913_n_20965 ( .a(FE_OCP_RBN1912_n_20965), .o(FE_OCP_RBN1913_n_20965) );
in01f80 FE_OCP_RBC1296_n_30451 ( .a(n_30451), .o(FE_OCP_RBN1296_n_30451) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_26_ ( .ck(newNet_1094), .d(n_11305), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_) );
no02f80 g749940 ( .a(n_30356), .b(n_30076), .o(n_30145) );
in01f80 g746968 ( .a(n_33075), .o(n_33157) );
in01f80 g772556 ( .a(n_8403), .o(n_8375) );
no02f80 g760463 ( .a(n_20093), .b(n_20092), .o(n_20146) );
in01f80 g738309 ( .a(n_41916), .o(n_41909) );
no02f80 g738203 ( .a(n_41966), .b(n_41965), .o(n_41967) );
in01f80 g753078 ( .a(n_27528), .o(n_27529) );
no02f80 g746922 ( .a(FE_OCP_RBN3390_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n_33401) );
na02f80 g777371 ( .a(n_3794), .b(n_3902), .o(n_3997) );
na02f80 g767391 ( .a(n_13310), .b(n_13244), .o(n_13390) );
na02f80 g740223 ( .a(n_39993), .b(FE_OCP_RBN3027_n_39942), .o(n_40063) );
in01f80 FE_OCP_RBC2807_n_30643 ( .a(n_30643), .o(FE_OCP_RBN2807_n_30643) );
in01f80 FE_OCPC1393_n_962 ( .a(n_962), .o(FE_OCPN1393_n_962) );
in01f80 g737214 ( .a(n_42990), .o(n_42991) );
oa12f80 g773228 ( .a(n_7604), .b(n_7603), .c(n_7602), .o(n_7950) );
oa22f80 FE_RC_3874_0 ( .a(FE_RN_1513_0), .b(FE_OCP_RBN2308_n_29298), .c(n_29379), .d(n_29298), .o(n_29399) );
oa22f80 g784553 ( .a(FE_OFN801_n_46285), .b(n_11356), .c(FE_OCP_RBN3044_n_46337), .d(n_11334), .o(n_46374) );
na02f80 g764260 ( .a(n_16388), .b(n_16456), .o(n_16488) );
oa22f80 g752758 ( .a(n_27851), .b(n_186), .c(n_27852), .d(n_179), .o(n_27957) );
na02f80 g740940 ( .a(n_39215), .b(n_39161), .o(n_39216) );
na02f80 g774947 ( .a(n_6103), .b(n_6084), .o(n_6196) );
in01f80 g751329 ( .a(n_29597), .o(n_29636) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_24_ ( .ck(newNet_2641), .d(FE_OCP_RBN3117_n_22710), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_) );
na02f80 g772667 ( .a(n_8255), .b(n_8245), .o(n_8246) );
na02f80 g737228 ( .a(n_42932), .b(n_42945), .o(n_43002) );
ao12f80 g779810 ( .a(n_2109), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .o(n_2124) );
in01f80 newInst_3266 ( .a(newNet_3265), .o(newNet_3266) );
oa12f80 g775688 ( .a(n_5108), .b(n_5084), .c(n_5032), .o(n_5192) );
oa12f80 g766829 ( .a(n_14427), .b(n_14947), .c(n_14299), .o(n_14428) );
no02f80 g756094 ( .a(n_24202), .b(n_24246), .o(n_24262) );
no02f80 g746342 ( .a(n_33475), .b(n_33474), .o(n_33476) );
no02f80 g738927 ( .a(n_41247), .b(n_41027), .o(n_41307) );
na02f80 g756714 ( .a(n_23543), .b(n_23571), .o(n_23595) );
na02f80 g771780 ( .a(n_9325), .b(n_9324), .o(n_9326) );
na02f80 g753323 ( .a(n_27125), .b(FE_RN_1356_0), .o(n_27101) );
in01f80 newInst_1819 ( .a(newNet_360), .o(newNet_1819) );
ao12f80 g751309 ( .a(n_28661), .b(n_28685), .c(n_28660), .o(n_29812) );
oa12f80 g770918 ( .a(n_10005), .b(n_10049), .c(n_10004), .o(n_10088) );
ao12f80 g752831 ( .a(n_28108), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n_28619) );
in01f80 FE_OCP_RBC2664_n_20333 ( .a(FE_OCP_RBN2663_n_20333), .o(FE_OCP_RBN2664_n_20333) );
in01f80 g737421 ( .a(n_42802), .o(n_42803) );
na02f80 g770127 ( .a(n_10809), .b(n_10791), .o(n_10850) );
ao12f80 g762933 ( .a(n_17745), .b(n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .o(n_17796) );
in01f80 g762784 ( .a(n_17964), .o(n_17965) );
in01f80 FE_OCPC858_n_45697 ( .a(FE_OCPN857_n_45697), .o(FE_OCPN858_n_45697) );
oa22f80 g743778 ( .a(n_36369), .b(n_36316), .c(n_36370), .d(n_36317), .o(n_36421) );
oa12f80 g750022 ( .a(n_29919), .b(FE_OCP_RBN3561_n_29857), .c(n_28995), .o(n_30460) );
oa12f80 g781165 ( .a(n_118), .b(n_182), .c(n_63), .o(n_189) );
na02f80 g755441 ( .a(n_24754), .b(n_24618), .o(n_24755) );
in01f80 FE_OCPC1458_n_18426 ( .a(FE_OCPN1457_n_18426), .o(FE_OCPN1458_n_18426) );
in01f80 FE_OCP_RBC2889_n_46957 ( .a(n_46957), .o(FE_OCP_RBN2889_n_46957) );
na02f80 g771079 ( .a(n_9907), .b(n_9906), .o(n_10034) );
na02f80 g755803 ( .a(n_24310), .b(n_22111), .o(n_24367) );
in01f80 g750056 ( .a(n_29958), .o(n_29959) );
no02f80 g766552 ( .a(n_13957), .b(n_13001), .o(n_13995) );
na02f80 g774213 ( .a(n_6813), .b(n_6766), .o(n_6814) );
na02f80 g763491 ( .a(n_16814), .b(FE_OCPN3180_FE_OCP_RBN2744_n_15319), .o(n_16838) );
in01f80 FE_OCPC1787_n_36034 ( .a(n_36034), .o(FE_OCPN1787_n_36034) );
na02f80 g737451 ( .a(n_42669), .b(n_42402), .o(n_42689) );
in01f80 newInst_1826 ( .a(newNet_988), .o(newNet_1826) );
in01f80 g748091 ( .a(n_31614), .o(n_31668) );
in01f80 fopt782857 ( .a(n_44288), .o(n_44287) );
in01f80 g773479 ( .a(n_7584), .o(n_7608) );
in01f80 g751313 ( .a(n_29649), .o(n_29708) );
na02f80 g781149 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_4_), .o(n_209) );
in01f80 newInst_3281 ( .a(newNet_3280), .o(newNet_3281) );
no02f80 g774167 ( .a(n_6565), .b(n_6415), .o(n_6576) );
ao12f80 g744201 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n_46215), .c(n_36747), .o(n_36863) );
in01f80 g743717 ( .a(n_36280), .o(n_36329) );
na02f80 g737576 ( .a(n_42332), .b(n_42402), .o(n_42376) );
in01f80 g746442 ( .a(n_36111), .o(n_35602) );
in01f80 newInst_760 ( .a(newNet_759), .o(newNet_760) );
in01f80 g775881 ( .a(n_5276), .o(n_5277) );
no02f80 g766581 ( .a(n_14087), .b(n_14050), .o(n_16111) );
na02f80 g760917 ( .a(n_19454), .b(n_18119), .o(n_19460) );
in01f80 FE_OCP_RBC2332_n_29380 ( .a(n_29380), .o(FE_OCP_RBN2332_n_29380) );
no02f80 g742236 ( .a(n_44881), .b(n_37653), .o(n_38079) );
in01f80 newInst_2675 ( .a(newNet_2528), .o(newNet_2675) );
no02f80 g773125 ( .a(n_7646), .b(n_7644), .o(n_7692) );
na02f80 g743400 ( .a(n_36671), .b(n_36652), .o(n_36715) );
in01f80 g751462 ( .a(n_28737), .o(n_28738) );
in01f80 newInst_1619 ( .a(newNet_1618), .o(newNet_1619) );
no02f80 g754522 ( .a(n_26513), .b(FE_OCPN928_n_26231), .o(n_26611) );
in01f80 g780222 ( .a(n_1134), .o(n_1120) );
in01f80 g737224 ( .a(n_42933), .o(n_42934) );
no02f80 g767290 ( .a(n_13511), .b(n_13510), .o(n_13517) );
in01f80 g749020 ( .a(n_31097), .o(n_31098) );
no02f80 g769329 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n_11863) );
na02f80 g756581 ( .a(n_23821), .b(n_23658), .o(n_23733) );
in01f80 g739741 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_19_), .o(n_40702) );
na02f80 g771363 ( .a(n_9149), .b(n_9047), .o(n_9150) );
no02f80 g760487 ( .a(n_19978), .b(n_19919), .o(n_19979) );
na02f80 g775086 ( .a(n_4904), .b(n_6035), .o(n_6157) );
oa12f80 g770296 ( .a(n_10641), .b(n_10650), .c(n_10640), .o(n_10739) );
oa22f80 g784371 ( .a(FE_OFN774_n_46137), .b(n_6392), .c(FE_OFN806_n_46196), .d(n_6419), .o(n_46177) );
in01f80 g743772 ( .a(n_36206), .o(n_36207) );
no02f80 g738490 ( .a(FE_OCP_RBN2316_n_41420), .b(n_41310), .o(n_41707) );
na02f80 g775929 ( .a(n_5394), .b(n_5289), .o(n_5579) );
na02f80 g759891 ( .a(n_20273), .b(FE_OFN751_n_45003), .o(n_20297) );
na02f80 g778361 ( .a(n_2493), .b(n_2520), .o(n_2559) );
na02f80 g749164 ( .a(n_30856), .b(n_30830), .o(n_30933) );
in01f80 newInst_1906 ( .a(newNet_1530), .o(newNet_1906) );
ao12f80 g765162 ( .a(n_15119), .b(n_15151), .c(n_15117), .o(n_15276) );
ao12f80 g751200 ( .a(n_28468), .b(n_28791), .c(n_28504), .o(n_28853) );
no02f80 g737499 ( .a(n_42538), .b(n_42537), .o(n_42539) );
na02f80 g769840 ( .a(n_11136), .b(n_11103), .o(n_11190) );
no02f80 g754220 ( .a(n_25915), .b(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .o(n_25943) );
na02f80 g770755 ( .a(n_9970), .b(n_9927), .o(n_9984) );
in01f80 g761836 ( .a(n_18379), .o(n_18347) );
in01f80 FE_RC_2499_0 ( .a(n_41782), .o(FE_RN_1013_0) );
in01f80 g755514 ( .a(n_24750), .o(n_24751) );
oa12f80 g757456 ( .a(n_22951), .b(n_23299), .c(n_22921), .o(n_23400) );
no02f80 g741163 ( .a(FE_OCP_RBN2635_n_38806), .b(n_38430), .o(n_38833) );
na02f80 g750694 ( .a(n_29368), .b(n_30136), .o(n_29393) );
oa12f80 g738871 ( .a(n_41308), .b(n_41307), .c(n_41306), .o(n_41347) );
in01f80 newInst_1126 ( .a(newNet_1125), .o(newNet_1126) );
na02f80 g778330 ( .a(n_2528), .b(n_2084), .o(n_2529) );
in01f80 g753405 ( .a(n_27657), .o(n_27626) );
na02f80 g743391 ( .a(n_36732), .b(n_36702), .o(n_36748) );
ao12f80 g739098 ( .a(n_41000), .b(n_40999), .c(n_40998), .o(n_41444) );
no02f80 g775416 ( .a(n_5540), .b(n_5500), .o(n_5575) );
na02f80 g755597 ( .a(n_24683), .b(n_24682), .o(n_24711) );
oa22f80 g746477 ( .a(n_33223), .b(n_33261), .c(n_33224), .d(n_33260), .o(n_34323) );
oa12f80 g775483 ( .a(n_5698), .b(n_5755), .c(n_5697), .o(n_5841) );
in01f80 newInst_3347 ( .a(newNet_3346), .o(newNet_3347) );
no02f80 g778719 ( .a(n_2277), .b(n_2276), .o(n_2366) );
oa22f80 FE_RC_1272_0 ( .a(n_9543), .b(n_9638), .c(n_9569), .d(n_9628), .o(n_9864) );
in01f80 FE_OCP_RBC2999_n_11004 ( .a(FE_OCP_RBN2997_n_11004), .o(FE_OCP_RBN2999_n_11004) );
in01f80 g760756 ( .a(n_20156), .o(n_20157) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_1_ ( .ck(newNet_345), .d(n_1340), .o(delay_xor_ln22_unr3_stage2_stallmux_q_1_) );
na02f80 g737492 ( .a(n_42554), .b(n_42316), .o(n_42564) );
in01f80 newInst_214 ( .a(newNet_213), .o(newNet_214) );
in01f80 newInst_1248 ( .a(newNet_506), .o(newNet_1248) );
in01f80 g758649 ( .a(n_21916), .o(n_21917) );
na02f80 g740085 ( .a(n_39975), .b(n_39943), .o(n_40038) );
oa12f80 g780776 ( .a(n_377), .b(n_455), .c(FE_OCPN1386_n_470), .o(n_471) );
no02f80 g773967 ( .a(n_6900), .b(n_6620), .o(n_6959) );
no02f80 g740634 ( .a(n_39603), .b(n_39610), .o(n_39633) );
na02f80 g740547 ( .a(n_39706), .b(n_39662), .o(n_39734) );
in01f80 FE_RC_2575_0 ( .a(FE_OFN817_n_2285), .o(FE_RN_1059_0) );
no02f80 g760821 ( .a(n_19517), .b(n_19469), .o(n_19537) );
na02f80 g743508 ( .a(n_37713), .b(n_46241), .o(n_37678) );
in01f80 FE_RC_2870_0 ( .a(n_23964), .o(FE_RN_1239_0) );
in01f80 g777618 ( .a(n_3542), .o(n_3543) );
ao12f80 g771493 ( .a(n_47244), .b(n_8922), .c(n_47243), .o(n_9093) );
in01f80 FE_OCP_RBC2684_n_35213 ( .a(n_35213), .o(FE_OCP_RBN2684_n_35213) );
in01f80 g758080 ( .a(n_22027), .o(n_22084) );
in01f80 g746411 ( .a(n_33534), .o(n_34143) );
oa12f80 g753465 ( .a(n_26764), .b(n_26788), .c(n_26658), .o(n_26808) );
in01f80 g749143 ( .a(n_32206), .o(n_32207) );
in01f80 g781311 ( .a(n_60), .o(n_61) );
oa12f80 g751817 ( .a(n_28225), .b(n_28255), .c(n_28224), .o(n_29420) );
na02f80 g742636 ( .a(n_37501), .b(n_37500), .o(n_37502) );
no02f80 g755791 ( .a(n_24396), .b(n_23878), .o(n_24445) );
in01f80 newInst_210 ( .a(newNet_209), .o(newNet_210) );
no02f80 g755362 ( .a(n_24785), .b(n_24837), .o(n_24879) );
in01f80 g778519 ( .a(n_2541), .o(n_2542) );
no02f80 g757105 ( .a(n_23536), .b(n_22980), .o(n_23619) );
oa22f80 g739202 ( .a(n_40840), .b(n_40846), .c(n_40892), .d(n_40847), .o(n_41389) );
ao22s80 g779074 ( .a(n_2087), .b(n_1854), .c(n_2067), .d(n_1855), .o(n_2119) );
na02f80 g750061 ( .a(n_29896), .b(FE_OCP_RBN2281_n_29111), .o(n_30114) );
in01f80 FE_OCP_RBC1358_FE_RN_677_0 ( .a(FE_RN_677_0), .o(FE_OCP_RBN1358_FE_RN_677_0) );
no02f80 g776089 ( .a(n_4842), .b(n_4657), .o(n_4763) );
na02f80 g758892 ( .a(FE_OCP_RBN3218_n_21358), .b(n_45026), .o(n_21437) );
na02f80 g756344 ( .a(n_24480), .b(n_24479), .o(n_24481) );
oa12f80 g755714 ( .a(n_24493), .b(n_24492), .c(n_24491), .o(n_24590) );
in01f80 g748363 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_7_), .o(n_32952) );
no02f80 g737470 ( .a(n_42686), .b(n_42701), .o(n_43070) );
no02f80 g775236 ( .a(n_5692), .b(n_5714), .o(n_5779) );
oa12f80 g757626 ( .a(n_22047), .b(n_22564), .c(n_22164), .o(n_22603) );
no02f80 g758761 ( .a(n_21581), .b(n_20018), .o(n_21620) );
in01f80 g775017 ( .a(n_6160), .o(n_6184) );
in01f80 g765738 ( .a(n_15441), .o(n_15514) );
in01f80 newInst_360 ( .a(newNet_359), .o(newNet_360) );
oa12f80 g752124 ( .a(n_27964), .b(n_28096), .c(n_28095), .o(n_28097) );
no02f80 g744936 ( .a(FE_OCP_RBN2562_n_34905), .b(n_30504), .o(n_34957) );
na02f80 g754564 ( .a(n_26710), .b(n_26639), .o(n_26681) );
no02f80 g771501 ( .a(n_9483), .b(n_9445), .o(n_9643) );
in01f80 g751003 ( .a(n_28872), .o(n_28873) );
no02f80 g738184 ( .a(n_41969), .b(n_41968), .o(n_41970) );
na02f80 g780141 ( .a(n_1147), .b(n_832), .o(n_1194) );
in01f80 FE_RC_2273_0 ( .a(n_17572), .o(FE_RN_846_0) );
na02f80 g736994 ( .a(n_43082), .b(n_43134), .o(n_43315) );
no02f80 g764738 ( .a(n_15847), .b(n_14588), .o(n_15946) );
oa12f80 g750983 ( .a(n_28632), .b(n_28933), .c(n_28485), .o(n_28974) );
in01f80 g766916 ( .a(n_14110), .o(n_14008) );
in01f80 g769738 ( .a(n_11287), .o(n_11288) );
no02f80 g745199 ( .a(n_36228), .b(n_36023), .o(n_36283) );
in01f80 FE_OCP_DRV_C3743_n_25400 ( .a(FE_OCP_DRV_N3742_n_25400), .o(FE_OCP_DRV_N3743_n_25400) );
in01f80 newInst_2845 ( .a(newNet_2844), .o(newNet_2845) );
in01f80 g781287 ( .a(state_cordic_1_), .o(n_66) );
no02f80 g777272 ( .a(n_3578), .b(n_2913), .o(n_3659) );
oa12f80 g756839 ( .a(n_23752), .b(n_23751), .c(n_23750), .o(n_23836) );
oa12f80 g745231 ( .a(n_36224), .b(n_36223), .c(n_36222), .o(n_36281) );
no02f80 g740793 ( .a(n_39350), .b(n_39364), .o(n_39407) );
oa12f80 g784660 ( .a(n_8520), .b(n_8421), .c(n_8466), .o(n_46990) );
oa22f80 g776957 ( .a(n_3781), .b(FE_OCP_RBN2535_n_47018), .c(n_3780), .d(FE_OCP_RBN2533_n_47018), .o(n_3968) );
no02f80 g746855 ( .a(n_33474), .b(n_32992), .o(n_33059) );
in01f80 FE_RC_4087_0 ( .a(n_16923), .o(FE_RN_1787_0) );
no02f80 g772956 ( .a(n_7927), .b(n_7913), .o(n_7928) );
in01f80 g765136 ( .a(n_15344), .o(n_15345) );
no02f80 g743385 ( .a(n_36585), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36634) );
no02f80 g741238 ( .a(FE_OCP_RBN2635_n_38806), .b(n_38435), .o(n_38882) );
in01f80 newInst_1276 ( .a(newNet_96), .o(newNet_1276) );
na02f80 g754433 ( .a(n_25635), .b(n_25399), .o(n_25636) );
na02f80 g750389 ( .a(n_29634), .b(n_29616), .o(n_29617) );
oa22f80 g746629 ( .a(n_33068), .b(n_32893), .c(n_33113), .d(n_32894), .o(n_34288) );
in01f80 g778897 ( .a(n_2256), .o(n_2277) );
in01f80 g760190 ( .a(n_20526), .o(n_20527) );
oa22f80 g776617 ( .a(n_4160), .b(n_3106), .c(n_4080), .d(n_3082), .o(n_4313) );
in01f80 newInst_2123 ( .a(newNet_942), .o(newNet_2123) );
oa22f80 g784350 ( .a(FE_OCP_RBN3075_FE_OFN807_n_46195), .b(n_5483), .c(FE_OFN775_n_46137), .d(n_5418), .o(n_46156) );
in01f80 g780197 ( .a(n_1167), .o(n_1154) );
na02f80 g770330 ( .a(FE_OCP_RBN2870_n_10480), .b(n_10542), .o(n_10544) );
in01f80 g743103 ( .a(n_37048), .o(n_37148) );
na02f80 g747153 ( .a(n_32856), .b(n_32853), .o(n_32854) );
in01f80 FE_RC_2289_0 ( .a(n_17611), .o(FE_RN_859_0) );
na02f80 FE_RC_2389_0 ( .a(FE_RN_932_0), .b(FE_RN_935_0), .o(FE_RN_936_0) );
in01f80 g762094 ( .a(n_18278), .o(n_18279) );
oa12f80 g765810 ( .a(n_14973), .b(n_14972), .c(n_14971), .o(n_15033) );
no02f80 g780453 ( .a(n_1203), .b(n_845), .o(n_798) );
na02f80 g777903 ( .a(n_3147), .b(n_2328), .o(n_3148) );
oa22f80 g744658 ( .a(n_36498), .b(n_36216), .c(n_36499), .d(n_36215), .o(n_36542) );
na02f80 g746609 ( .a(n_34388), .b(n_33910), .o(n_34499) );
ao12f80 g742940 ( .a(n_36998), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n_37059) );
oa12f80 g748663 ( .a(n_31205), .b(n_31204), .c(n_31203), .o(n_31267) );
in01f80 newInst_979 ( .a(newNet_978), .o(newNet_979) );
in01f80 g742227 ( .a(n_38291), .o(n_38292) );
no02f80 g755257 ( .a(n_25040), .b(n_25015), .o(n_25114) );
na02f80 g753108 ( .a(n_27143), .b(n_27142), .o(n_27184) );
na02f80 g749858 ( .a(FE_OCP_RBN3019_n_31117), .b(n_31184), .o(n_31289) );
na02f80 g777347 ( .a(FE_OCP_RBN2730_n_4219), .b(FE_OFN821_n_4632), .o(n_4702) );
oa12f80 g772906 ( .a(n_7871), .b(n_7902), .c(n_7870), .o(n_9151) );
no02f80 g778187 ( .a(n_2860), .b(n_2675), .o(n_2932) );
ao12f80 g745728 ( .a(n_34866), .b(n_35390), .c(n_34888), .o(n_35432) );
no02f80 g780541 ( .a(n_713), .b(n_46055), .o(n_767) );
in01f80 g764899 ( .a(n_15652), .o(n_15598) );
in01f80 newInst_567 ( .a(newNet_566), .o(newNet_567) );
na02f80 g768553 ( .a(n_12313), .b(n_12263), .o(n_12328) );
in01f80 g749809 ( .a(n_31621), .o(n_31622) );
in01f80 newInst_405 ( .a(newNet_404), .o(newNet_405) );
na02f80 g737916 ( .a(n_42277), .b(n_42276), .o(n_42577) );
in01f80 newInst_3086 ( .a(newNet_3085), .o(newNet_3086) );
no02f80 g753261 ( .a(n_27377), .b(n_25915), .o(n_27378) );
in01f80 g751905 ( .a(n_29069), .o(n_29124) );
na02f80 g743548 ( .a(n_37585), .b(n_46203), .o(n_37673) );
in01f80 FE_OCP_RBC2289_n_2314 ( .a(n_2314), .o(FE_OCP_RBN2289_n_2314) );
no02f80 g757032 ( .a(n_23803), .b(n_23978), .o(n_23955) );
no02f80 FE_RC_1761_0 ( .a(n_12170), .b(FE_RN_502_0), .o(FE_RN_503_0) );
oa12f80 g745038 ( .a(n_34856), .b(n_34855), .c(n_34854), .o(n_35567) );
no02f80 g744727 ( .a(n_35155), .b(FE_OCPN1796_n_30546), .o(n_35294) );
na02f80 FE_RC_440_0 ( .a(FE_RN_123_0), .b(FE_RN_124_0), .o(FE_RN_125_0) );
no02f80 g746605 ( .a(n_34612), .b(n_34611), .o(n_34635) );
na02f80 g755472 ( .a(n_24582), .b(n_25316), .o(n_24625) );
in01f80 FE_OCPC3763_n_34222 ( .a(FE_OCPN3762_n_34222), .o(FE_OCPN3763_n_34222) );
no02f80 g774470 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .o(n_6620) );
in01f80 g746638 ( .a(n_33368), .o(n_33407) );
in01f80 FE_OCP_RBC3728_FE_RN_1787_0 ( .a(FE_RN_1787_0), .o(FE_OCP_RBN3728_FE_RN_1787_0) );
in01f80 newInst_2024 ( .a(newNet_1740), .o(newNet_2024) );
in01f80 g767736 ( .a(FE_OCP_RBN2202_n_12808), .o(n_12846) );
no02f80 g757017 ( .a(n_24188), .b(n_23804), .o(n_24234) );
oa12f80 g739045 ( .a(n_41076), .b(n_41075), .c(n_41074), .o(n_41124) );
na02f80 g744650 ( .a(n_35251), .b(n_35121), .o(n_35273) );
in01f80 newInst_1288 ( .a(newNet_1287), .o(newNet_1288) );
in01f80 FE_RC_3529_0 ( .a(n_45224), .o(FE_RN_1526_0) );
in01f80 newInst_3231 ( .a(newNet_3230), .o(newNet_3231) );
in01f80 FE_OCP_RBC2914_n_42947 ( .a(n_42947), .o(FE_OCP_RBN2914_n_42947) );
in01f80 newInst_818 ( .a(newNet_817), .o(newNet_818) );
in01f80 FE_OCP_RBC2200_n_13889 ( .a(n_13889), .o(FE_OCP_RBN2200_n_13889) );
in01f80 g761006 ( .a(n_19325), .o(n_19326) );
in01f80 FE_OCPC1459_n_37232 ( .a(n_37232), .o(FE_OCPN1459_n_37232) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_15_ ( .ck(newNet_186), .d(n_46356), .o(delay_xor_ln22_unr9_stage4_stallmux_q_15_) );
na02f80 g759766 ( .a(n_21624), .b(n_21668), .o(n_21669) );
in01f80 g741057 ( .a(n_39189), .o(n_39190) );
no02f80 FE_RC_2811_0 ( .a(n_9726), .b(FE_RN_1202_0), .o(FE_RN_1203_0) );
no02f80 g760532 ( .a(n_20450), .b(n_20424), .o(n_20425) );
ao12f80 g758774 ( .a(n_21473), .b(n_21679), .c(n_21544), .o(n_21707) );
in01f80 FE_OCP_RBC1184_n_14638 ( .a(n_14638), .o(FE_OCP_RBN1184_n_14638) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_13_ ( .ck(newNet_922), .d(n_27855), .o(delay_xor_ln21_unr18_stage7_stallmux_q_13_) );
na02f80 g753631 ( .a(n_26630), .b(n_26319), .o(n_26661) );
no02f80 g740806 ( .a(n_39293), .b(n_39140), .o(n_39356) );
na02f80 g739750 ( .a(n_40466), .b(n_40196), .o(n_40475) );
no02f80 g750821 ( .a(n_29210), .b(n_29055), .o(n_29212) );
in01f80 g745542 ( .a(n_35511), .o(n_35540) );
in01f80 g764198 ( .a(n_16535), .o(n_16494) );
in01f80 FE_OFC735_n_22641 ( .a(FE_OFN734_n_22641), .o(FE_OFN735_n_22641) );
no02f80 g762981 ( .a(n_17938), .b(n_17431), .o(n_18034) );
no02f80 g778620 ( .a(n_2273), .b(n_2266), .o(n_2295) );
na02f80 g755102 ( .a(n_25173), .b(n_24098), .o(n_25323) );
in01f80 newInst_2763 ( .a(newNet_2762), .o(newNet_2763) );
in01f80 newInst_3289 ( .a(newNet_1709), .o(newNet_3289) );
na02f80 g741060 ( .a(n_38832), .b(n_38894), .o(n_38969) );
in01f80 g748739 ( .a(n_32584), .o(n_32585) );
na02f80 g736677 ( .a(n_43281), .b(n_43229), .o(n_43413) );
na02f80 g749652 ( .a(n_30155), .b(n_30179), .o(n_32076) );
in01f80 newInst_3364 ( .a(newNet_282), .o(newNet_3364) );
in01f80 newInst_3543 ( .a(newNet_3542), .o(newNet_3543) );
ao12f80 FE_RC_2035_0 ( .a(FE_RN_679_0), .b(n_25824), .c(n_25893), .o(n_25982) );
oa12f80 g761797 ( .a(n_18815), .b(n_19125), .c(n_18655), .o(n_19232) );
oa12f80 g747767 ( .a(n_33413), .b(n_33571), .c(n_33441), .o(n_33889) );
in01f80 FE_OCP_RBC3407_n_28597 ( .a(FE_OCP_RBN3405_n_28597), .o(FE_OCP_RBN3407_n_28597) );
na02f80 g780185 ( .a(n_1116), .b(n_1148), .o(n_1117) );
in01f80 newInst_1585 ( .a(newNet_1584), .o(newNet_1585) );
in01f80 g758563 ( .a(n_22585), .o(n_22586) );
oa22f80 FE_RC_1243_0 ( .a(FE_OCP_RBN3517_n_8498), .b(FE_OCP_RBN2495_n_8641), .c(FE_OCP_RBN3518_n_8498), .d(FE_OCP_RBN2496_n_8641), .o(n_8838) );
na02f80 g743346 ( .a(n_36655), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36712) );
oa12f80 g766986 ( .a(n_13763), .b(n_13762), .c(n_13761), .o(n_14303) );
no02f80 g762681 ( .a(n_17928), .b(n_17926), .o(n_17927) );
in01f80 FE_OCP_RBC2242_n_13017 ( .a(n_13017), .o(FE_OCP_RBN2242_n_13017) );
in01f80 g780117 ( .a(n_1205), .o(n_1200) );
na02f80 g755318 ( .a(n_25472), .b(n_25471), .o(n_25473) );
no02f80 g742751 ( .a(n_37393), .b(n_37392), .o(n_37391) );
in01f80 FE_OCP_RBC3060_FE_RN_640_0 ( .a(FE_RN_640_0), .o(FE_OCP_RBN3060_FE_RN_640_0) );
in01f80 FE_RC_3552_0 ( .a(n_18343), .o(FE_RN_1541_0) );
na02f80 g746962 ( .a(n_32836), .b(n_32878), .o(n_32893) );
in01f80 newInst_1635 ( .a(newNet_1634), .o(newNet_1635) );
in01f80 g778419 ( .a(n_2728), .o(n_3594) );
in01f80 newInst_3244 ( .a(newNet_2325), .o(newNet_3244) );
na02f80 g740184 ( .a(FE_OCP_RBN3715_n_39913), .b(n_39553), .o(n_40069) );
in01f80 FE_RC_2946_0 ( .a(n_22063), .o(FE_RN_1286_0) );
in01f80 newInst_1876 ( .a(newNet_900), .o(newNet_1876) );
in01f80 g771694 ( .a(n_9070), .o(n_9071) );
na02f80 g751453 ( .a(n_28722), .b(n_28721), .o(n_28739) );
na02f80 g764321 ( .a(n_16678), .b(n_16103), .o(n_16798) );
na02f80 g738748 ( .a(n_41384), .b(n_41383), .o(n_41443) );
in01f80 FE_OCP_RBC3426_n_44881 ( .a(n_44881), .o(FE_OCP_RBN3426_n_44881) );
in01f80 g767022 ( .a(n_14108), .o(n_14109) );
na02f80 g749412 ( .a(n_30535), .b(n_30292), .o(n_30564) );
in01f80 FE_OCP_RBC3737_n_12027 ( .a(n_12027), .o(FE_OCP_RBN3737_n_12027) );
na02f80 g736915 ( .a(FE_OCPN912_n_43022), .b(n_42802), .o(n_43110) );
na02f80 FE_RC_2037_0 ( .a(n_26727), .b(FE_RN_680_0), .o(FE_RN_681_0) );
in01f80 newInst_2110 ( .a(newNet_290), .o(newNet_2110) );
no02f80 g752957 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .o(n_28018) );
no02f80 g766019 ( .a(n_14706), .b(n_14782), .o(n_14808) );
ao22s80 g740520 ( .a(n_39734), .b(n_39735), .c(n_39744), .d(n_39743), .o(n_39769) );
in01f80 FE_OCP_RBC3306_n_44722 ( .a(FE_OCP_RBN3307_n_44722), .o(FE_OCP_RBN3306_n_44722) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_23_ ( .ck(newNet_3220), .d(n_36487), .o(delay_add_ln22_unr23_stage9_stallmux_q_23_) );
in01f80 newInst_1022 ( .a(newNet_912), .o(newNet_1022) );
na02f80 g742676 ( .a(n_37454), .b(n_37270), .o(n_37522) );
no02f80 g780872 ( .a(n_521), .b(n_7), .o(n_532) );
na02f80 g781016 ( .a(cos_out_25), .b(n_43918), .o(n_339) );
in01f80 newInst_1448 ( .a(newNet_1447), .o(newNet_1448) );
in01f80 newInst_1380 ( .a(newNet_1379), .o(newNet_1380) );
in01f80 FE_OCP_RBC3682_n_26171 ( .a(n_26171), .o(FE_OCP_RBN3682_n_26171) );
in01f80 newInst_429 ( .a(newNet_428), .o(newNet_429) );
no03m80 FE_RC_77_0 ( .a(n_17684), .b(n_17655), .c(n_17683), .o(n_17720) );
na02f80 g764871 ( .a(FE_OCP_RBN2878_n_15553), .b(n_15648), .o(n_15688) );
na03f80 FE_RC_591_0 ( .a(n_41978), .b(n_41774), .c(n_41973), .o(n_42005) );
na02f80 g743864 ( .a(n_46250), .b(n_46229), .o(n_37025) );
in01f80 FE_OCP_RBC1836_FE_RN_1542_0 ( .a(FE_RN_1542_0), .o(FE_OCP_RBN1836_FE_RN_1542_0) );
in01f80 g768370 ( .a(n_12520), .o(n_12521) );
in01f80 g759849 ( .a(FE_OCPN1482_n_22207), .o(n_22393) );
na02f80 g750808 ( .a(n_29092), .b(n_28701), .o(n_29122) );
ao12f80 g744626 ( .a(n_35883), .b(n_36574), .c(n_35961), .o(n_36638) );
no02f80 g771229 ( .a(n_9837), .b(n_9905), .o(n_10002) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_28_ ( .ck(newNet_1587), .d(n_27625), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_) );
no02f80 g775179 ( .a(FE_OCP_RBN3045_n_5881), .b(FE_OCPN1028_n_4182), .o(n_5964) );
no02f80 g747591 ( .a(n_31704), .b(n_32200), .o(n_32244) );
in01f80 g749107 ( .a(n_31026), .o(n_31081) );
oa22f80 g747888 ( .a(n_31884), .b(n_31917), .c(n_31883), .d(n_31916), .o(n_31999) );
in01f80 g740762 ( .a(n_39516), .o(n_39517) );
in01f80 g769430 ( .a(n_11439), .o(n_11455) );
in01f80 FE_OCP_RBC3494_n_19390 ( .a(FE_OCP_RBN3493_n_19390), .o(FE_OCP_RBN3494_n_19390) );
no02f80 g766989 ( .a(n_13572), .b(n_13592), .o(n_13689) );
no02f80 g774146 ( .a(n_6590), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n_6896) );
in01f80 g745102 ( .a(n_34728), .o(n_34753) );
in01f80 g741641 ( .a(n_38912), .o(n_38588) );
no02f80 g745967 ( .a(n_33946), .b(n_33945), .o(n_34013) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_1_ ( .ck(newNet_564), .d(n_16636), .o(delay_xor_ln22_unr12_stage5_stallmux_q_1_) );
na02f80 g770561 ( .a(n_10278), .b(n_9121), .o(n_10279) );
ao12f80 g754963 ( .a(n_25840), .b(n_25868), .c(n_25839), .o(n_26509) );
no02f80 g741287 ( .a(n_44954), .b(n_38471), .o(n_38909) );
na02f80 g754346 ( .a(n_25821), .b(n_25788), .o(n_25893) );
na02f80 g780164 ( .a(n_1162), .b(n_1155), .o(n_1156) );
in01f80 g761068 ( .a(n_19181), .o(n_19182) );
ao12f80 g756064 ( .a(n_25026), .b(n_24541), .c(n_25109), .o(n_25119) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_11_ ( .ck(newNet_1038), .d(n_17731), .o(delay_xor_ln21_unr12_stage5_stallmux_q_11_) );
in01f80 g750014 ( .a(n_31044), .o(n_31040) );
oa12f80 g738245 ( .a(n_41826), .b(n_41919), .c(n_41879), .o(n_41944) );
no02f80 g752143 ( .a(n_28068), .b(n_28067), .o(n_28121) );
na02f80 g751178 ( .a(n_29909), .b(n_29908), .o(n_30000) );
oa12f80 g776148 ( .a(n_4649), .b(n_4806), .c(n_4735), .o(n_4942) );
ao22s80 g777961 ( .a(n_3673), .b(FE_OCP_RBN2297_n_2438), .c(n_3155), .d(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(n_3189) );
no02f80 g764660 ( .a(n_15811), .b(n_15516), .o(n_15907) );
in01f80 g776374 ( .a(n_4787), .o(n_4918) );
in01f80 g753775 ( .a(n_26495), .o(n_26496) );
in01f80 g753472 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_5_), .o(n_28124) );
na02f80 g773144 ( .a(FE_OCP_RBN2229_n_7598), .b(n_7714), .o(n_7768) );
in01f80 FE_OCP_RBC2759_n_9843 ( .a(n_9843), .o(FE_OCP_RBN2759_n_9843) );
ao12f80 g749668 ( .a(n_29888), .b(n_30057), .c(n_29955), .o(n_30080) );
in01f80 g778145 ( .a(n_2884), .o(n_2942) );
no02f80 g773210 ( .a(n_7802), .b(n_7853), .o(n_7997) );
no02f80 g779587 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .o(n_1759) );
in01f80 g776334 ( .a(n_4319), .o(n_4320) );
in01f80 newInst_600 ( .a(newNet_599), .o(newNet_600) );
no02f80 g748398 ( .a(n_31730), .b(n_31599), .o(n_31733) );
no02f80 g769589 ( .a(n_11381), .b(n_11380), .o(n_11405) );
no02f80 g754274 ( .a(n_26689), .b(n_26384), .o(n_26909) );
na02f80 g753831 ( .a(n_26370), .b(n_26369), .o(n_26371) );
in01f80 g750619 ( .a(n_29418), .o(n_29419) );
na02f80 g760151 ( .a(n_20432), .b(n_20430), .o(n_20482) );
in01f80 newInst_2056 ( .a(newNet_2055), .o(newNet_2056) );
ao22s80 g772269 ( .a(n_8760), .b(n_8087), .c(n_8690), .d(n_8086), .o(n_9994) );
no02f80 g769896 ( .a(n_10970), .b(n_11011), .o(n_11128) );
na02f80 g742878 ( .a(n_37228), .b(n_37227), .o(n_37229) );
in01f80 newInst_3751 ( .a(newNet_3750), .o(newNet_3751) );
no02f80 g747747 ( .a(n_33762), .b(n_33571), .o(n_33989) );
in01f80 g772820 ( .a(n_8074), .o(n_8075) );
ao12f80 g768996 ( .a(n_11780), .b(FE_OCP_RBN2116_n_45224), .c(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .o(n_11815) );
in01f80 newInst_1665 ( .a(newNet_1664), .o(newNet_1665) );
na02f80 g740035 ( .a(n_39802), .b(n_39822), .o(n_39823) );
na02f80 g738163 ( .a(n_41979), .b(n_41860), .o(n_42030) );
in01f80 FE_RC_151_0 ( .a(n_17888), .o(FE_RN_45_0) );
in01f80 g770351 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .o(n_10708) );
in01f80 g756513 ( .a(n_23714), .o(n_23715) );
in01f80 FE_OCP_RBC3690_n_16146 ( .a(n_16146), .o(FE_OCP_RBN3690_n_16146) );
na02f80 g737391 ( .a(n_42751), .b(n_42465), .o(n_42791) );
no02f80 g741109 ( .a(n_39043), .b(n_39000), .o(n_39001) );
in01f80 g756686 ( .a(n_23572), .o(n_23843) );
na02f80 g773834 ( .a(n_7053), .b(n_5671), .o(n_7116) );
ao12f80 g763790 ( .a(n_16854), .b(n_16853), .c(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n_18483) );
in01f80 newInst_3494 ( .a(newNet_3493), .o(newNet_3494) );
in01f80 g745274 ( .a(n_36681), .o(n_35725) );
in01f80 FE_OCPC1770_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(FE_OCPN1769_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
no02f80 g774466 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n_6826) );
no02f80 g766320 ( .a(n_14703), .b(n_14076), .o(n_14780) );
in01f80 g745068 ( .a(n_36313), .o(n_36314) );
in01f80 g760737 ( .a(n_19736), .o(n_19693) );
in01f80 g776465 ( .a(n_4671), .o(n_4646) );
no02f80 g781307 ( .a(beta_31), .b(beta_14), .o(n_81) );
in01f80 g764512 ( .a(n_16095), .o(n_16013) );
in01f80 FE_RC_3946_0 ( .a(FE_RN_1708_0), .o(FE_RN_1707_0) );
in01f80 newInst_1475 ( .a(newNet_201), .o(newNet_1475) );
in01f80 g755536 ( .a(n_24776), .o(n_24777) );
in01f80 g775659 ( .a(n_5266), .o(n_5267) );
na02f80 g737386 ( .a(n_42796), .b(n_42627), .o(n_42810) );
in01f80 g777732 ( .a(n_3509), .o(n_3510) );
in01f80 g771024 ( .a(n_9926), .o(n_9979) );
in01f80 FE_RC_4210_0 ( .a(FE_RN_1844_0), .o(n_14612) );
oa12f80 g746184 ( .a(n_33590), .b(n_33711), .c(n_33591), .o(n_33830) );
na02f80 g743220 ( .a(n_36873), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .o(n_36944) );
in01f80 newInst_1856 ( .a(newNet_1855), .o(newNet_1856) );
in01f80 FE_OCP_RBC3360_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(FE_OCP_RBN3296_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3360_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
in01f80 g760517 ( .a(n_19972), .o(n_19997) );
no02f80 g759242 ( .a(n_21156), .b(n_21078), .o(n_21266) );
na02f80 g749910 ( .a(n_29965), .b(n_29870), .o(n_30265) );
no02f80 g781215 ( .a(n_94), .b(n_93), .o(n_95) );
oa22f80 g739896 ( .a(n_40369), .b(n_40389), .c(n_40370), .d(n_40388), .o(n_40439) );
no02f80 g750472 ( .a(n_29574), .b(n_29573), .o(n_29590) );
in01f80 g769119 ( .a(n_11747), .o(n_11748) );
in01f80 FE_OCP_RBC3247_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3247_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01f80 FE_RC_1939_0 ( .a(n_28566), .o(FE_RN_618_0) );
in01f80 FE_OFC787_n_25834 ( .a(FE_OFN786_n_25834), .o(FE_OFN787_n_25834) );
oa12f80 g776263 ( .a(n_4480), .b(n_4786), .c(n_4582), .o(n_4806) );
in01f80 g751196 ( .a(n_29937), .o(n_29997) );
na02f80 g736617 ( .a(n_43194), .b(n_43093), .o(n_43334) );
no02f80 g744099 ( .a(n_35688), .b(n_44180), .o(n_35783) );
na02f80 g780210 ( .a(n_1069), .b(n_1180), .o(n_1030) );
in01f80 g773793 ( .a(n_7159), .o(n_7150) );
na02f80 g744849 ( .a(n_35095), .b(n_35136), .o(n_35137) );
no02f80 g776023 ( .a(n_4838), .b(n_4423), .o(n_4902) );
na02f80 g749088 ( .a(n_30941), .b(n_30935), .o(n_31018) );
in01f80 FE_OCP_RBC2492_n_8508 ( .a(n_8508), .o(FE_OCP_RBN2492_n_8508) );
in01f80 g768151 ( .a(n_13017), .o(n_13634) );
na02f80 g773558 ( .a(n_7402), .b(n_7401), .o(n_7444) );
in01f80 FE_OCPC941_n_44925 ( .a(FE_OCP_RBN2548_n_44944), .o(FE_OCPN941_n_44925) );
no02f80 g778235 ( .a(n_2763), .b(n_2828), .o(n_2748) );
no02f80 g767810 ( .a(n_12763), .b(n_13634), .o(n_13349) );
no02f80 FE_RC_2168_0 ( .a(FE_RN_769_0), .b(n_21157), .o(FE_RN_770_0) );
in01f80 FE_RC_3492_0 ( .a(FE_RN_1505_0), .o(FE_RN_1500_0) );
no02f80 FE_RC_2517_0 ( .a(FE_RN_1023_0), .b(FE_RN_1024_0), .o(n_31239) );
in01f80 g756228 ( .a(n_24813), .o(n_25132) );
na02f80 g753254 ( .a(n_27110), .b(n_27142), .o(n_27227) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_31_ ( .ck(newNet_2357), .d(n_36567), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_) );
in01f80 FE_OCP_RBC2993_n_35539 ( .a(FE_OCP_RBN2990_n_35539), .o(FE_OCP_RBN2993_n_35539) );
na02f80 g781336 ( .a(n_7), .b(beta_19), .o(n_70) );
in01f80 g775654 ( .a(n_5424), .o(n_5425) );
na02f80 g756710 ( .a(n_23480), .b(n_23479), .o(n_23481) );
no02f80 g761487 ( .a(n_19569), .b(n_18777), .o(n_19713) );
no02f80 g756925 ( .a(n_23778), .b(n_23748), .o(n_24113) );
in01f80 g740995 ( .a(n_38934), .o(n_39065) );
no02f80 g778685 ( .a(n_2438), .b(n_2432), .o(n_2651) );
no02f80 g758851 ( .a(n_21475), .b(n_45081), .o(n_21505) );
in01f80 FE_OCPC3777_n_43019 ( .a(FE_OCPN3776_n_43019), .o(FE_OCPN3777_n_43019) );
no02f80 g767703 ( .a(n_13350), .b(n_13349), .o(n_13824) );
no02f80 g738943 ( .a(n_41171), .b(n_40908), .o(n_41172) );
in01f80 g767864 ( .a(n_12836), .o(n_12777) );
in01f80 FE_OCP_RBC2373_n_8221 ( .a(FE_OCP_RBN2371_n_8221), .o(FE_OCP_RBN2373_n_8221) );
in01f80 g746615 ( .a(n_34545), .o(n_34546) );
ao12f80 g742467 ( .a(n_37551), .b(n_37644), .c(n_37604), .o(n_37648) );
in01f80 g777880 ( .a(n_3261), .o(n_3262) );
no02f80 FE_RC_2133_0 ( .a(FE_RN_744_0), .b(n_25920), .o(FE_RN_745_0) );
in01f80 g766975 ( .a(n_13846), .o(n_13847) );
no02f80 g755407 ( .a(n_24808), .b(n_24759), .o(n_24830) );
na02f80 g776511 ( .a(n_4479), .b(FE_OCP_RBN2491_n_3338), .o(n_4542) );
in01f80 g738670 ( .a(n_41608), .o(n_41658) );
in01f80 g766658 ( .a(n_13931), .o(n_13988) );
in01f80 g737768 ( .a(n_42629), .o(n_42630) );
in01f80 newInst_3417 ( .a(newNet_1223), .o(newNet_3417) );
no02f80 g777776 ( .a(FE_OCP_RBN2486_n_3498), .b(n_2913), .o(n_3333) );
in01f80 g749576 ( .a(n_31780), .o(n_31752) );
in01f80 g781200 ( .a(n_362), .o(n_176) );
na02f80 g765332 ( .a(FE_OCP_RBN3620_n_15135), .b(n_15299), .o(n_15407) );
in01f80 newInst_955 ( .a(newNet_954), .o(newNet_955) );
ao12f80 g773931 ( .a(n_6843), .b(n_6984), .c(n_6891), .o(n_7055) );
no02f80 g744515 ( .a(n_35400), .b(n_35303), .o(n_35422) );
na02f80 g739233 ( .a(n_41053), .b(n_41039), .o(n_41070) );
ao22s80 g741483 ( .a(n_38749), .b(n_38726), .c(n_38748), .d(n_38727), .o(n_38792) );
no02f80 g742412 ( .a(n_37720), .b(n_37649), .o(n_37723) );
no02f80 g750705 ( .a(n_29365), .b(n_29135), .o(n_29412) );
in01f80 g757387 ( .a(n_22970), .o(n_22971) );
in01f80 g779431 ( .a(n_2116), .o(n_2117) );
in01f80 g744256 ( .a(n_36135), .o(n_36136) );
in01f80 newInst_3078 ( .a(newNet_3077), .o(newNet_3078) );
in01f80 g744368 ( .a(n_46217), .o(n_36852) );
in01f80 FE_OCPC1764_n_13646 ( .a(FE_OCPN1763_n_13646), .o(FE_OCPN1764_n_13646) );
ao22s80 FE_RC_1954_0 ( .a(n_18032), .b(FE_OCP_RBN3837_n_19513), .c(n_19418), .d(n_19513), .o(n_19633) );
in01f80 FE_OCP_RBC3528_n_13765 ( .a(FE_OCP_RBN3527_n_13765), .o(FE_OCP_RBN3528_n_13765) );
na02f80 g777166 ( .a(n_4999), .b(n_4817), .o(n_5862) );
na02f80 g761830 ( .a(n_19097), .b(n_18697), .o(n_19126) );
in01f80 g770415 ( .a(n_10609), .o(n_10610) );
in01f80 g780928 ( .a(n_463), .o(n_464) );
in01f80 g778311 ( .a(n_2835), .o(n_2836) );
in01f80 g762431 ( .a(n_18090), .o(n_18074) );
no02f80 g741137 ( .a(n_39395), .b(n_39041), .o(n_39423) );
in01f80 newInst_3598 ( .a(newNet_3597), .o(newNet_3598) );
na02f80 g743202 ( .a(n_37175), .b(n_36944), .o(n_36928) );
ao12f80 g738446 ( .a(n_41471), .b(n_41660), .c(n_41156), .o(n_41869) );
no02f80 FE_RC_2821_0 ( .a(n_34316), .b(n_34377), .o(FE_RN_1210_0) );
in01f80 g741228 ( .a(n_39453), .o(n_39454) );
in01f80 g771909 ( .a(n_9020), .o(n_9021) );
no02f80 g761823 ( .a(n_18375), .b(n_18483), .o(n_18894) );
in01f80 FE_RC_3747_0 ( .a(FE_RN_1644_0), .o(FE_OCPN1748_n_23354) );
no02f80 g756748 ( .a(n_23991), .b(n_23990), .o(n_23992) );
no02f80 g780380 ( .a(n_907), .b(n_1203), .o(n_964) );
in01f80 newInst_6 ( .a(newNet_5), .o(newNet_6) );
in01f80 FE_OCP_DRV_C1574_n_28869 ( .a(FE_OCP_DRV_N1573_n_28869), .o(FE_OCP_DRV_N1574_n_28869) );
oa12f80 g758908 ( .a(n_21472), .b(n_21471), .c(n_21470), .o(n_21541) );
ao12f80 g745182 ( .a(n_34602), .b(n_34601), .c(n_34600), .o(n_34712) );
ao12f80 g784675 ( .a(n_4772), .b(n_4743), .c(n_4609), .o(n_47005) );
na02f80 FE_RC_3663_0 ( .a(FE_RN_1608_0), .b(n_21874), .o(n_21940) );
no02f80 g769212 ( .a(n_12011), .b(n_11934), .o(n_12087) );
in01f80 g766212 ( .a(n_14417), .o(n_14418) );
oa12f80 g755391 ( .a(n_22111), .b(n_24701), .c(n_24507), .o(n_24703) );
in01f80 g739844 ( .a(n_40301), .o(n_40302) );
na02f80 g778709 ( .a(n_2365), .b(n_2394), .o(n_2371) );
no02f80 g759538 ( .a(n_20881), .b(n_20906), .o(n_21029) );
na02f80 g742546 ( .a(n_37558), .b(n_37576), .o(n_37656) );
no02f80 g763236 ( .a(n_17243), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .o(n_17279) );
oa12f80 g762168 ( .a(n_18088), .b(n_18138), .c(n_18045), .o(n_18196) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_8_ ( .ck(newNet_2137), .d(n_928), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_) );
in01f80 g749394 ( .a(n_30729), .o(n_30757) );
in01f80 g748204 ( .a(n_33281), .o(n_32802) );
ao12f80 g739247 ( .a(n_40859), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n_41287) );
in01f80 g757549 ( .a(n_23322), .o(n_22984) );
in01f80 FE_OCP_RBC2468_n_8767 ( .a(n_8767), .o(FE_OCP_RBN2468_n_8767) );
ao12f80 g780690 ( .a(n_654), .b(n_653), .c(n_652), .o(n_906) );
in01f80 g776212 ( .a(n_5015), .o(n_5016) );
in01f80 g768170 ( .a(n_13515), .o(n_14376) );
no03m80 g738317 ( .a(n_41460), .b(n_41818), .c(n_41683), .o(n_41757) );
in01f80 FE_OFC805_n_46196 ( .a(FE_OFN804_n_46196), .o(FE_OFN805_n_46196) );
no02f80 g748165 ( .a(n_31863), .b(n_30738), .o(n_31904) );
no02f80 g746800 ( .a(n_32973), .b(n_32972), .o(n_33488) );
in01f80 g767323 ( .a(n_13436), .o(n_13456) );
in01f80 newInst_2935 ( .a(newNet_2934), .o(newNet_2935) );
in01f80 g748702 ( .a(n_33240), .o(n_33256) );
in01f80 newInst_1996 ( .a(newNet_1378), .o(newNet_1996) );
in01f80 g762390 ( .a(n_18608), .o(n_18609) );
in01f80 g772000 ( .a(n_9825), .o(n_9826) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_1_ ( .ck(newNet_1117), .d(n_9437), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_) );
na02f80 g778106 ( .a(n_2827), .b(n_2896), .o(n_2949) );
in01f80 FE_OFC813_n_2540 ( .a(FE_OFN830_n_2540), .o(FE_OFN813_n_2540) );
ao12f80 g777797 ( .a(n_2687), .b(n_3227), .c(n_2701), .o(n_3435) );
in01f80 g744348 ( .a(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41337) );
in01f80 FE_RC_2234_0 ( .a(n_23057), .o(FE_RN_814_0) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_12_ ( .ck(newNet_1140), .d(n_10549), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_) );
in01f80 g742977 ( .a(n_36973), .o(n_37073) );
in01f80 g760446 ( .a(n_20095), .o(n_20096) );
oa12f80 g744621 ( .a(n_35136), .b(n_35272), .c(n_35134), .o(n_35329) );
no02f80 g777861 ( .a(n_3212), .b(n_2713), .o(n_3227) );
na02f80 g762392 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18494), .o(n_18657) );
na02f80 g741409 ( .a(n_38800), .b(FE_OCPN3174_n_38799), .o(n_38804) );
oa12f80 g781086 ( .a(n_72), .b(n_258), .c(n_140), .o(n_267) );
in01f80 g764841 ( .a(n_15734), .o(n_15692) );
in01f80 g761160 ( .a(n_19168), .o(n_19169) );
na02f80 g744512 ( .a(n_35413), .b(n_35342), .o(n_35444) );
in01f80 g742903 ( .a(n_37124), .o(n_37125) );
no02f80 g755818 ( .a(n_24268), .b(n_23925), .o(n_24295) );
no02f80 g769377 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n_12007) );
no02f80 g768308 ( .a(n_12531), .b(n_12368), .o(n_12561) );
na02f80 g741457 ( .a(n_38793), .b(n_38789), .o(n_38811) );
in01f80 g775873 ( .a(n_5372), .o(n_5373) );
in01f80 g761350 ( .a(n_18952), .o(n_18982) );
no02f80 g742258 ( .a(n_44871), .b(n_37414), .o(n_37880) );
in01f80 g736296 ( .a(n_43882), .o(n_43883) );
na02f80 g767558 ( .a(n_13052), .b(n_12768), .o(n_13093) );
in01f80 g739902 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .o(n_40480) );
in01f80 newInst_2227 ( .a(newNet_1741), .o(newNet_2227) );
in01f80 g750572 ( .a(n_29450), .o(n_30214) );
oa12f80 g749602 ( .a(n_30484), .b(n_30483), .c(n_30482), .o(n_30572) );
na02f80 g744601 ( .a(FE_OCP_RBN1372_n_35275), .b(n_35237), .o(n_35297) );
in01f80 g741908 ( .a(n_38242), .o(n_38358) );
in01f80 g772838 ( .a(n_8057), .o(n_8124) );
na02f80 g755750 ( .a(n_24404), .b(n_24373), .o(n_24447) );
ao22s80 g776753 ( .a(n_3812), .b(n_2912), .c(n_3736), .d(n_2911), .o(n_3981) );
oa12f80 g757372 ( .a(n_23037), .b(n_23036), .c(n_23035), .o(n_24142) );
in01f80 FE_OCP_RBC1348_n_19270 ( .a(FE_OCP_RBN1347_n_19270), .o(FE_OCP_RBN1348_n_19270) );
in01f80 g757402 ( .a(n_22967), .o(n_22968) );
in01f80 g748355 ( .a(n_31827), .o(n_31828) );
no02f80 g756434 ( .a(n_23614), .b(n_23639), .o(n_23667) );
na02f80 g767476 ( .a(n_13229), .b(n_13098), .o(n_13230) );
in01f80 g766446 ( .a(n_14120), .o(n_14191) );
oa12f80 g761717 ( .a(n_19297), .b(n_19296), .c(n_19295), .o(n_19398) );
na02f80 g775662 ( .a(n_5565), .b(n_5584), .o(n_5566) );
no02f80 g778515 ( .a(n_2521), .b(n_3286), .o(n_2522) );
in01f80 g736602 ( .a(n_43335), .o(n_43378) );
in01f80 newInst_1357 ( .a(newNet_99), .o(newNet_1357) );
no02f80 g738476 ( .a(n_41387), .b(n_41412), .o(n_41426) );
oa22f80 g745342 ( .a(n_35956), .b(n_35583), .c(FE_OCP_RBN2995_n_35539), .d(n_35559), .o(n_36223) );
in01f80 FE_OCP_RBC2605_FE_OCPN899_n_44593 ( .a(FE_OCPN899_n_44593), .o(FE_OCP_RBN2605_FE_OCPN899_n_44593) );
no02f80 g737693 ( .a(n_42216), .b(n_42286), .o(n_42566) );
ao22s80 FE_RC_1438_0 ( .a(n_31802), .b(n_44358), .c(n_31803), .d(n_32169), .o(n_32254) );
in01f80 FE_OCP_RBC3550_n_44575 ( .a(FE_OCP_RBN3543_n_44575), .o(FE_OCP_RBN3550_n_44575) );
in01f80 g779478 ( .a(n_2028), .o(n_2029) );
in01f80 drc784142 ( .a(n_45890), .o(n_45891) );
in01f80 g764317 ( .a(n_16397), .o(n_16396) );
in01f80 fopt783438 ( .a(n_45013), .o(n_45032) );
na02f80 g752817 ( .a(n_27986), .b(n_27877), .o(n_28135) );
na02f80 g765498 ( .a(n_15664), .b(n_15823), .o(n_15867) );
in01f80 g738984 ( .a(n_41220), .o(n_41221) );
na02f80 g777649 ( .a(n_3468), .b(n_3498), .o(n_3499) );
na02f80 g766209 ( .a(n_14535), .b(n_14376), .o(n_14656) );
in01f80 g745852 ( .a(n_34114), .o(n_34115) );
in01f80 g736417 ( .a(n_43747), .o(n_43759) );
in01f80 FE_OCP_RBC3612_FE_OCPN1797_n_20333 ( .a(FE_OCP_RBN3611_FE_OCPN1797_n_20333), .o(FE_OCP_RBN3612_FE_OCPN1797_n_20333) );
in01f80 newInst_2929 ( .a(newNet_1564), .o(newNet_2929) );
na02f80 g741577 ( .a(n_38686), .b(n_38685), .o(n_38687) );
no02f80 g776699 ( .a(n_4115), .b(n_4222), .o(n_4273) );
in01f80 newInst_158 ( .a(newNet_157), .o(newNet_158) );
na02f80 g775825 ( .a(n_5076), .b(FE_OCPN846_n_4046), .o(n_5097) );
oa12f80 g747631 ( .a(n_32070), .b(n_32300), .c(n_31869), .o(n_32330) );
na02f80 g777097 ( .a(n_3605), .b(n_4759), .o(n_5355) );
no02f80 g761016 ( .a(n_19177), .b(FE_OFN780_n_17093), .o(n_19216) );
oa12f80 g756380 ( .a(n_23959), .b(n_24277), .c(n_23953), .o(n_24417) );
ao12f80 g738602 ( .a(n_41725), .b(n_41716), .c(n_41656), .o(n_42020) );
in01f80 newInst_1814 ( .a(newNet_1813), .o(newNet_1814) );
in01f80 g772782 ( .a(n_8127), .o(n_8128) );
in01f80 FE_OCP_RBC2712_n_35075 ( .a(FE_OCP_RBN2711_n_35075), .o(FE_OCP_RBN2712_n_35075) );
ao22s80 g742035 ( .a(FE_OCP_RBN3445_n_37945), .b(n_37554), .c(FE_OCP_RBN3441_n_37945), .d(n_37569), .o(n_38422) );
oa22f80 FE_RC_3440_0 ( .a(n_22339), .b(n_22722), .c(n_22338), .d(n_22756), .o(n_22914) );
in01f80 newInst_1423 ( .a(newNet_1163), .o(newNet_1423) );
no02f80 g740044 ( .a(n_39865), .b(n_39921), .o(n_39922) );
in01f80 g780441 ( .a(n_788), .o(n_762) );
no02f80 g764415 ( .a(n_16013), .b(n_14452), .o(n_16233) );
na02f80 g739584 ( .a(n_40604), .b(n_44610), .o(n_40617) );
ao12f80 g778560 ( .a(n_2440), .b(n_2441), .c(n_2439), .o(n_2570) );
no02f80 FE_RC_1242_0 ( .a(FE_RN_372_0), .b(FE_RN_373_0), .o(FE_RN_374_0) );
no02f80 g769809 ( .a(n_11132), .b(n_44511), .o(n_11194) );
in01f80 g736441 ( .a(n_43779), .o(n_43780) );
ao12f80 g773040 ( .a(n_7817), .b(n_7889), .c(n_7888), .o(n_8027) );
in01f80 g758429 ( .a(n_23259), .o(n_23317) );
na02f80 g753764 ( .a(n_26398), .b(n_23353), .o(n_26448) );
no02f80 g751480 ( .a(n_28678), .b(n_28599), .o(n_28703) );
in01f80 newInst_625 ( .a(newNet_22), .o(newNet_625) );
na02f80 g744306 ( .a(n_44180), .b(n_35165), .o(n_36096) );
in01f80 g780459 ( .a(n_846), .o(n_836) );
in01f80 FE_RC_3830_0 ( .a(FE_OCPN908_n_23227), .o(FE_RN_1670_0) );
na02f80 g769702 ( .a(n_11345), .b(n_11289), .o(n_11331) );
no02f80 g759677 ( .a(n_21409), .b(n_21450), .o(n_21451) );
oa12f80 g751292 ( .a(n_29050), .b(n_29649), .c(n_29308), .o(n_29724) );
na02f80 g771994 ( .a(n_44498), .b(n_9939), .o(n_10077) );
in01f80 g757849 ( .a(n_22356), .o(n_22357) );
oa12f80 g742014 ( .a(n_38006), .b(FE_OCP_RBN3445_n_37945), .c(n_37983), .o(n_38374) );
in01f80 newInst_2035 ( .a(newNet_466), .o(newNet_2035) );
in01f80 g744737 ( .a(n_35152), .o(n_35180) );
no02f80 g775996 ( .a(n_4729), .b(n_4591), .o(n_4736) );
in01f80 g767015 ( .a(n_14171), .o(n_14136) );
na02f80 g777405 ( .a(n_3649), .b(n_3701), .o(n_3727) );
in01f80 g746765 ( .a(n_33143), .o(n_33144) );
oa22f80 g758702 ( .a(n_21683), .b(n_21734), .c(n_21682), .d(n_21735), .o(n_21810) );
no02f80 g773082 ( .a(n_7886), .b(n_8150), .o(n_8118) );
na02f80 g750537 ( .a(n_29427), .b(n_29406), .o(n_29500) );
in01f80 g742043 ( .a(n_38201), .o(n_38202) );
no02f80 FE_RC_2816_0 ( .a(n_34423), .b(n_34908), .o(FE_RN_1206_0) );
in01f80 g767621 ( .a(n_12888), .o(n_12940) );
in01f80 FE_OCP_RBC2762_n_15200 ( .a(n_15200), .o(FE_OCP_RBN2762_n_15200) );
no02f80 g748315 ( .a(n_31787), .b(n_32149), .o(n_31842) );
no02f80 g754363 ( .a(n_25733), .b(n_25415), .o(n_25764) );
no02f80 g769654 ( .a(n_11258), .b(n_11194), .o(n_11323) );
na02f80 g747048 ( .a(n_34022), .b(n_34021), .o(n_34023) );
no02f80 g776242 ( .a(n_47006), .b(n_47341), .o(n_4962) );
oa12f80 g743495 ( .a(n_36624), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .c(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_37625) );
no02f80 g746580 ( .a(n_34810), .b(n_34613), .o(n_35070) );
na02f80 g762403 ( .a(FE_OCP_RBN3409_n_45120), .b(n_17786), .o(n_18614) );
na02f80 g760225 ( .a(FE_OCP_RBN1332_n_20249), .b(FE_OCP_RBN1351_n_19148), .o(n_20304) );
in01f80 FE_RC_3710_0 ( .a(FE_RN_635_0), .o(FE_RN_1631_0) );
no02f80 FE_RC_2028_0 ( .a(FE_RN_674_0), .b(n_25847), .o(FE_RN_675_0) );
oa22f80 g784541 ( .a(n_11759), .b(FE_OFN801_n_46285), .c(n_11669), .d(FE_OCP_RBN3043_n_46337), .o(n_46362) );
oa22f80 FE_RC_725_0 ( .a(n_7452), .b(n_8295), .c(n_8294), .d(n_7453), .o(n_8402) );
na02f80 g744293 ( .a(FE_OCP_RBN2902_n_44174), .b(n_34946), .o(n_35856) );
no02f80 g779631 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_16_), .o(n_1764) );
na02f80 g769181 ( .a(n_12050), .b(n_11862), .o(n_12066) );
na02f80 g761964 ( .a(n_18224), .b(n_17186), .o(n_18301) );
na02f80 g764697 ( .a(n_15853), .b(n_15374), .o(n_15855) );
na02f80 g760923 ( .a(n_19360), .b(n_18010), .o(n_19505) );
no02f80 g755724 ( .a(n_24325), .b(n_23885), .o(n_24327) );
oa22f80 FE_RC_949_0 ( .a(n_20231), .b(n_22835), .c(n_22580), .d(n_22804), .o(n_22913) );
no02f80 g753888 ( .a(n_26184), .b(n_24590), .o(n_26337) );
na02f80 g747092 ( .a(n_32928), .b(n_32665), .o(n_32930) );
na02f80 g745600 ( .a(n_34286), .b(n_34313), .o(n_34383) );
na02f80 g753757 ( .a(n_26378), .b(n_26175), .o(n_26379) );
no02f80 g774349 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_16_), .o(n_6998) );
na02f80 g740111 ( .a(n_40069), .b(n_40178), .o(n_40277) );
in01f80 g737445 ( .a(n_42731), .o(n_42732) );
in01f80 g775605 ( .a(n_5484), .o(n_5485) );
in01f80 FE_OCP_RBC2997_n_11004 ( .a(FE_OCP_RBN2996_n_11004), .o(FE_OCP_RBN2997_n_11004) );
in01f80 g768189 ( .a(FE_OCP_RBN2250_n_13017), .o(n_13469) );
in01f80 g763786 ( .a(n_16749), .o(n_16750) );
no02f80 g739131 ( .a(n_40962), .b(n_40832), .o(n_41014) );
in01f80 g777083 ( .a(n_3795), .o(n_3885) );
in01f80 g758380 ( .a(FE_OFN735_n_22641), .o(n_22782) );
na02f80 g759252 ( .a(n_21152), .b(n_21180), .o(n_21305) );
in01f80 FE_OCP_RBC3398_n_37624 ( .a(n_37624), .o(FE_OCP_RBN3398_n_37624) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_9_ ( .ck(newNet_3090), .d(n_40440), .o(delay_add_ln22_unr27_stage10_stallmux_q_9_) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_27_ ( .ck(newNet_1091), .d(n_11344), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_) );
na02f80 g773644 ( .a(n_7343), .b(n_7177), .o(n_7370) );
in01f80 fopt783454 ( .a(FE_OFN751_n_45003), .o(n_45060) );
no02f80 g775781 ( .a(n_5509), .b(FE_OCP_RBN3590_n_47014), .o(n_5877) );
in01f80 g764517 ( .a(n_16089), .o(n_16118) );
in01f80 newInst_2277 ( .a(newNet_255), .o(newNet_2277) );
no02f80 g740595 ( .a(n_39577), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39596) );
in01f80 g763814 ( .a(n_17574), .o(n_17531) );
in01f80 g767458 ( .a(n_14968), .o(n_14966) );
in01f80 g736534 ( .a(n_43696), .o(n_43697) );
in01f80 g780325 ( .a(n_984), .o(n_1040) );
no02f80 g760645 ( .a(n_19730), .b(n_18032), .o(n_19754) );
in01f80 g777174 ( .a(n_5191), .o(n_5329) );
no02f80 g779402 ( .a(n_1478), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n_1690) );
no02f80 g775711 ( .a(n_5426), .b(n_5310), .o(n_5449) );
na02f80 g762414 ( .a(FE_OCP_RBN3410_n_45120), .b(n_18422), .o(n_18522) );
ao12f80 g749715 ( .a(n_31346), .b(n_31255), .c(n_31311), .o(n_31347) );
na02f80 g769877 ( .a(n_11096), .b(n_10921), .o(n_11133) );
in01f80 FE_OCP_RBC2130_n_32647 ( .a(n_32647), .o(FE_OCP_RBN2130_n_32647) );
no02f80 g758717 ( .a(n_21741), .b(n_21620), .o(n_21766) );
no02f80 g770748 ( .a(FE_OCP_RBN3652_n_10100), .b(FE_OCP_RBN2524_n_8951), .o(n_10768) );
na02f80 g763361 ( .a(n_16938), .b(n_16753), .o(n_16999) );
no02f80 g768749 ( .a(n_12128), .b(n_12127), .o(n_12180) );
no02f80 g742682 ( .a(n_37518), .b(n_38235), .o(n_37519) );
na02f80 g774370 ( .a(n_6703), .b(n_6722), .o(n_7564) );
ao12f80 g742762 ( .a(n_37347), .b(n_37346), .c(n_37345), .o(n_37894) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_21_ ( .ck(newNet_1740), .d(n_22567), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_) );
no02f80 g751741 ( .a(n_29246), .b(n_28993), .o(n_28994) );
na02f80 g779753 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .o(n_1558) );
in01f80 g757289 ( .a(n_23204), .o(n_23205) );
oa22f80 g770543 ( .a(FE_OCP_RBN2794_n_10106), .b(n_10733), .c(n_10278), .d(n_9200), .o(n_10469) );
in01f80 FE_OCP_RBC3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN3361_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
na02f80 g770882 ( .a(n_9968), .b(n_9900), .o(n_10053) );
no02f80 g777090 ( .a(n_3890), .b(n_3698), .o(n_4025) );
in01f80 g775074 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .o(n_6123) );
na02f80 g759454 ( .a(n_20910), .b(n_45032), .o(n_20939) );
no02f80 g754356 ( .a(n_25730), .b(FE_OCPN1514_FE_OFN738_n_22641), .o(n_25791) );
in01f80 g742585 ( .a(n_37965), .o(n_38325) );
no02f80 g752281 ( .a(n_28098), .b(n_27865), .o(n_27866) );
ao12f80 g762305 ( .a(n_18387), .b(n_18386), .c(n_18385), .o(n_18773) );
in01f80 g780601 ( .a(n_690), .o(n_691) );
no02f80 g780498 ( .a(n_1027), .b(n_1026), .o(n_1043) );
na02f80 g769838 ( .a(n_11129), .b(n_10983), .o(n_11208) );
na02f80 g780511 ( .a(n_951), .b(n_914), .o(n_999) );
na02f80 FE_RC_308_0 ( .a(FE_RN_90_0), .b(FE_RN_91_0), .o(FE_RN_92_0) );
na02f80 FE_RC_1743_0 ( .a(n_12375), .b(n_12252), .o(n_12450) );
no02f80 g762275 ( .a(n_18692), .b(n_18765), .o(n_19575) );
in01f80 g738090 ( .a(n_42091), .o(n_42092) );
na02f80 g766273 ( .a(n_14153), .b(n_14196), .o(n_14288) );
in01f80 g752329 ( .a(n_27831), .o(n_27832) );
na02f80 g772404 ( .a(n_8526), .b(FE_OCPN1011_n_7802), .o(n_8595) );
in01f80 g762736 ( .a(n_17849), .o(n_17850) );
no02f80 g749315 ( .a(n_30626), .b(FE_OCP_RBN2804_n_30534), .o(n_30654) );
na02f80 g770284 ( .a(n_10485), .b(n_47263), .o(n_10517) );
no02f80 g762746 ( .a(FE_OCPN854_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .o(n_17920) );
in01f80 FE_OCP_RBC2593_n_25181 ( .a(n_25181), .o(FE_OCP_RBN2593_n_25181) );
in01f80 g770796 ( .a(n_10181), .o(n_10220) );
in01f80 newInst_2659 ( .a(newNet_2195), .o(newNet_2659) );
no02f80 FE_RC_55_0 ( .a(FE_RN_14_0), .b(n_4470), .o(n_47007) );
in01f80 FE_RC_4155_0 ( .a(n_32835), .o(FE_RN_1808_0) );
na02f80 g756429 ( .a(n_23997), .b(n_23994), .o(n_24039) );
na02f80 FE_RC_2251_0 ( .a(FE_RN_822_0), .b(FE_RN_829_0), .o(n_37353) );
in01f80 g767213 ( .a(n_14215), .o(n_14340) );
ao12f80 g739167 ( .a(n_40924), .b(n_40938), .c(n_40923), .o(n_41412) );
in01f80 newInst_1486 ( .a(newNet_1485), .o(newNet_1486) );
oa12f80 g742576 ( .a(n_37470), .b(n_37469), .c(n_37468), .o(n_37935) );
na02f80 g763932 ( .a(n_17015), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .o(n_17207) );
no02f80 g775208 ( .a(n_5856), .b(n_5858), .o(n_5955) );
in01f80 g751718 ( .a(n_28373), .o(n_28335) );
no02f80 g741867 ( .a(n_38206), .b(n_38123), .o(n_38288) );
ao12f80 g739257 ( .a(n_40705), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_15_), .o(n_41143) );
no02f80 g746538 ( .a(n_34475), .b(n_34418), .o(n_34527) );
oa12f80 g740945 ( .a(n_39246), .b(n_39252), .c(n_39199), .o(n_39283) );
na02f80 g760342 ( .a(n_20123), .b(n_20213), .o(n_20241) );
na02f80 g761728 ( .a(n_19296), .b(n_19295), .o(n_19297) );
no02f80 g744251 ( .a(n_35487), .b(n_34516), .o(n_35533) );
na02f80 g748446 ( .a(n_31720), .b(n_31719), .o(n_31799) );
na02f80 FE_RC_3473_0 ( .a(FE_RN_1492_0), .b(n_39220), .o(n_39293) );
no02f80 g749352 ( .a(n_30580), .b(n_30584), .o(n_30659) );
no02f80 g778909 ( .a(FE_OCP_RBN2288_n_2268), .b(n_1998), .o(n_2338) );
in01f80 g769777 ( .a(n_11303), .o(n_11304) );
oa12f80 g738903 ( .a(n_41284), .b(n_41283), .c(n_41282), .o(n_41543) );
na02f80 g775935 ( .a(n_5208), .b(n_5207), .o(n_5209) );
in01f80 g762322 ( .a(n_18185), .o(n_18186) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_12_ ( .ck(newNet_3650), .d(n_16602), .o(delay_add_ln22_unr11_stage5_stallmux_q_12_) );
oa22f80 g757914 ( .a(n_22110), .b(n_21998), .c(n_22086), .d(n_21997), .o(n_22236) );
in01f80 g756058 ( .a(n_25195), .o(n_25161) );
in01f80 g743650 ( .a(n_36412), .o(n_36413) );
in01f80 g769098 ( .a(n_11596), .o(n_11597) );
in01f80 FE_OCP_RBC2290_n_2438 ( .a(n_2438), .o(FE_OCP_RBN2290_n_2438) );
in01f80 FE_OCPC1861_n_30319 ( .a(n_30319), .o(FE_OCPN1861_n_30319) );
in01f80 g763545 ( .a(n_16912), .o(n_16919) );
in01f80 g771045 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_2_), .o(n_9949) );
no02f80 g769040 ( .a(FE_OCP_RBN2116_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_7_), .o(n_11694) );
na02f80 g762444 ( .a(n_18046), .b(n_18088), .o(n_18107) );
no02f80 g766498 ( .a(n_14118), .b(FE_OCP_RBN2208_n_12907), .o(n_14146) );
oa12f80 g738261 ( .a(n_41847), .b(n_41846), .c(n_41845), .o(n_41952) );
oa22f80 g749286 ( .a(n_32006), .b(n_31619), .c(n_32007), .d(n_31620), .o(n_32093) );
in01f80 g773489 ( .a(n_7502), .o(n_7503) );
no02f80 FE_RC_2117_0 ( .a(n_24142), .b(n_24341), .o(FE_RN_735_0) );
in01f80 newInst_3686 ( .a(newNet_3685), .o(newNet_3686) );
na02f80 g767680 ( .a(n_13370), .b(n_13421), .o(n_13463) );
in01f80 g750036 ( .a(n_30385), .o(n_30386) );
na02f80 g775494 ( .a(n_5608), .b(n_5650), .o(n_5684) );
in01f80 g741277 ( .a(n_38988), .o(n_38943) );
in01f80 FE_RC_3652_0 ( .a(FE_OCPN1491_n_22036), .o(FE_RN_1603_0) );
no02f80 g761182 ( .a(n_19080), .b(n_18674), .o(n_19150) );
in01f80 FE_RC_2303_0 ( .a(n_25199), .o(FE_RN_871_0) );
na02f80 g766127 ( .a(n_14573), .b(n_14593), .o(n_14658) );
in01f80 FE_OCP_RBC2573_n_29922 ( .a(FE_OCP_RBN2570_n_29922), .o(FE_OCP_RBN2573_n_29922) );
oa12f80 g766770 ( .a(n_13573), .b(n_13693), .c(FE_OCP_RBN2244_n_13017), .o(n_13725) );
in01f80 g774547 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_23_), .o(n_6413) );
in01f80 g760881 ( .a(n_19474), .o(n_19435) );
in01f80 g741604 ( .a(n_38629), .o(n_38643) );
na02f80 g754116 ( .a(n_26114), .b(n_26113), .o(n_26115) );
na02f80 g759110 ( .a(n_21317), .b(FE_OCP_RBN3684_FE_RN_770_0), .o(n_21351) );
in01f80 g738389 ( .a(n_41708), .o(n_41709) );
in01f80 newInst_2824 ( .a(newNet_987), .o(newNet_2824) );
oa12f80 g747301 ( .a(n_32791), .b(n_32529), .c(n_44962), .o(n_32711) );
no02f80 g744207 ( .a(n_36132), .b(n_35617), .o(n_36256) );
no02f80 g776745 ( .a(n_4056), .b(n_3961), .o(n_4229) );
in01f80 g746959 ( .a(n_33210), .o(n_33211) );
in01f80 FE_OCP_RBC2925_n_10525 ( .a(n_10525), .o(FE_OCP_RBN2925_n_10525) );
na02f80 g781236 ( .a(n_64), .b(n_118), .o(n_131) );
ao12f80 g774522 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_6733) );
no02f80 g756570 ( .a(n_23572), .b(n_23611), .o(n_23632) );
na02f80 g756846 ( .a(n_23393), .b(n_23374), .o(n_23557) );
no02f80 g755402 ( .a(n_24832), .b(n_24834), .o(n_24833) );
na02f80 g760454 ( .a(n_20559), .b(n_20558), .o(n_20560) );
no02f80 g755497 ( .a(n_24578), .b(n_24318), .o(n_24701) );
na02f80 g770406 ( .a(n_10479), .b(n_10331), .o(n_10567) );
in01f80 fopt783528 ( .a(n_15510), .o(n_45139) );
in01f80 FE_OCP_RBC3640_n_44490 ( .a(n_44490), .o(FE_OCP_RBN3640_n_44490) );
in01f80 FE_OCP_RBC3073_n_43230 ( .a(FE_OCP_RBN3069_n_43230), .o(FE_OCP_RBN3073_n_43230) );
no02f80 g751489 ( .a(n_28816), .b(n_28867), .o(n_28885) );
na02f80 g777171 ( .a(n_5001), .b(n_4884), .o(n_5990) );
no02f80 g754218 ( .a(n_26037), .b(n_23354), .o(n_26038) );
na02f80 g745621 ( .a(n_34369), .b(n_33735), .o(n_34621) );
na02f80 g758813 ( .a(n_22177), .b(n_22176), .o(n_22178) );
no02f80 g739432 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n_40771) );
na02f80 g743299 ( .a(n_37899), .b(n_37898), .o(n_37959) );
in01f80 g778086 ( .a(n_3597), .o(n_3080) );
na02f80 g763603 ( .a(n_16855), .b(n_16826), .o(n_16898) );
oa12f80 g772318 ( .a(n_8088), .b(n_8613), .c(n_8079), .o(n_8684) );
in01f80 g750405 ( .a(n_29657), .o(n_29695) );
in01f80 newInst_3665 ( .a(newNet_3664), .o(newNet_3665) );
na02f80 g758168 ( .a(FE_OCPN1249_n_44267), .b(FE_OCP_RBN1913_n_20965), .o(n_22271) );
in01f80 g741763 ( .a(FE_OCP_RBN2349_n_38515), .o(n_38917) );
in01f80 g737842 ( .a(n_42216), .o(n_42285) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_17_ ( .ck(newNet_2963), .d(n_6154), .o(delay_add_ln22_unr5_stage3_stallmux_q_17_) );
na02f80 g737314 ( .a(n_42860), .b(n_42473), .o(n_42876) );
in01f80 g770636 ( .a(n_10328), .o(n_10354) );
na02f80 g749868 ( .a(FE_OCP_RBN3011_n_31117), .b(n_31214), .o(n_31312) );
no02f80 g746826 ( .a(n_32957), .b(n_32996), .o(n_33019) );
in01f80 FE_OCP_DRV_C1602_n_21639 ( .a(FE_OCP_DRV_N1601_n_21639), .o(FE_OCP_DRV_N1602_n_21639) );
ao22s80 g775373 ( .a(n_5503), .b(n_5479), .c(n_5487), .d(n_5478), .o(n_5656) );
in01f80 FE_RC_2592_0 ( .a(FE_RN_1073_0), .o(n_6891) );
no02f80 g761652 ( .a(n_19496), .b(n_19049), .o(n_19548) );
na02f80 g766066 ( .a(n_14554), .b(FE_OCP_RBN3532_n_13765), .o(n_14586) );
in01f80 g752562 ( .a(n_27714), .o(n_27683) );
in01f80 FE_OCPC1045_n_13570 ( .a(n_13570), .o(FE_OCPN1045_n_13570) );
na02f80 g756920 ( .a(n_23932), .b(n_23952), .o(n_23953) );
in01f80 newInst_28 ( .a(newNet_5), .o(newNet_28) );
in01f80 g747037 ( .a(n_32863), .o(n_32860) );
in01f80 g737773 ( .a(n_42627), .o(n_42628) );
in01f80 g757959 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_), .o(n_23056) );
na02f80 FE_RC_2688_0 ( .a(FE_RN_1124_0), .b(n_9080), .o(FE_RN_1125_0) );
in01f80 newInst_2066 ( .a(newNet_2065), .o(newNet_2066) );
na02f80 g771110 ( .a(n_9795), .b(n_9844), .o(n_9989) );
in01f80 g756505 ( .a(n_23919), .o(n_23920) );
na03f80 g743439 ( .a(n_37614), .b(n_37730), .c(n_37539), .o(n_37731) );
na02f80 g754897 ( .a(n_25481), .b(n_24632), .o(n_25625) );
na02f80 FE_RC_4238_0 ( .a(FE_RN_1861_0), .b(n_31126), .o(n_31196) );
no02f80 g771877 ( .a(n_8748), .b(n_7570), .o(n_8863) );
in01f80 FE_RC_2601_0 ( .a(n_18051), .o(FE_RN_1079_0) );
oa12f80 g749739 ( .a(FE_OCP_RBN3017_n_31117), .b(n_31509), .c(n_31256), .o(n_31292) );
in01f80 FE_OCP_RBC2852_n_26169 ( .a(n_26169), .o(FE_OCP_RBN2852_n_26169) );
no02f80 g767039 ( .a(FE_OCP_RBN2457_n_13765), .b(n_13795), .o(n_13939) );
oa12f80 g776852 ( .a(n_2948), .b(n_3633), .c(n_2887), .o(n_3830) );
na02f80 g774725 ( .a(n_45474), .b(n_6292), .o(n_6363) );
oa12f80 g761296 ( .a(n_19129), .b(n_19128), .c(n_19127), .o(n_20885) );
ao22s80 g756894 ( .a(n_24188), .b(n_24088), .c(n_24059), .d(n_23641), .o(n_24907) );
na02f80 g748981 ( .a(n_31127), .b(n_31021), .o(n_31128) );
ao12f80 g741226 ( .a(n_38995), .b(FE_OCP_RBN3579_n_44944), .c(n_38955), .o(n_39391) );
in01f80 g759973 ( .a(n_20500), .o(n_20540) );
in01f80 newInst_2388 ( .a(newNet_2387), .o(newNet_2388) );
ao22s80 g737235 ( .a(n_42894), .b(n_42759), .c(n_42895), .d(n_42758), .o(n_42962) );
no02f80 g764466 ( .a(n_16571), .b(n_15974), .o(n_16632) );
no02f80 FE_RC_3559_0 ( .a(FE_RN_1544_0), .b(n_29628), .o(FE_RN_1545_0) );
in01f80 newInst_2446 ( .a(newNet_1981), .o(newNet_2446) );
no02f80 g776109 ( .a(n_5063), .b(n_5062), .o(n_5203) );
in01f80 FE_OCP_RBC2717_n_14982 ( .a(FE_OCP_RBN2716_n_14982), .o(FE_OCP_RBN2717_n_14982) );
in01f80 g778244 ( .a(n_2760), .o(n_2761) );
oa12f80 g776545 ( .a(n_4420), .b(n_4432), .c(n_4419), .o(n_4526) );
in01f80 FE_OCP_RBC3589_n_47014 ( .a(n_47014), .o(FE_OCP_RBN3589_n_47014) );
in01f80 g759425 ( .a(n_21114), .o(n_21115) );
no02f80 g746696 ( .a(n_34276), .b(n_33815), .o(n_34359) );
in01f80 FE_RC_3899_0 ( .a(FE_RN_1282_0), .o(FE_RN_1693_0) );
oa12f80 g762600 ( .a(n_18295), .b(n_18294), .c(n_18293), .o(n_18572) );
ao12f80 g738103 ( .a(n_42058), .b(n_42057), .c(n_42056), .o(n_42116) );
na02f80 g753148 ( .a(n_27334), .b(n_27227), .o(n_27457) );
na02f80 g765359 ( .a(n_15332), .b(n_15331), .o(n_15333) );
na02f80 g764241 ( .a(n_16493), .b(FE_OCP_RBN1184_n_14638), .o(n_16515) );
ao12f80 g752161 ( .a(n_27973), .b(n_28009), .c(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n_28099) );
in01f80 g777037 ( .a(n_3758), .o(n_3759) );
no02f80 g748728 ( .a(n_31242), .b(n_31243), .o(n_31329) );
na02f80 FE_RC_2752_0 ( .a(FE_RN_1169_0), .b(n_43833), .o(FE_RN_1170_0) );
no02f80 g760170 ( .a(n_20363), .b(n_20366), .o(n_20434) );
na02f80 g759623 ( .a(n_21301), .b(n_21454), .o(n_21380) );
ao12f80 g755166 ( .a(n_25690), .b(n_25714), .c(n_25689), .o(n_26507) );
na02f80 g743370 ( .a(n_37813), .b(n_36814), .o(n_37828) );
in01f80 g769353 ( .a(n_11798), .o(n_11611) );
in01f80 newInst_2951 ( .a(newNet_1435), .o(newNet_2951) );
in01f80 newInst_2549 ( .a(newNet_2548), .o(newNet_2549) );
no02f80 g777137 ( .a(n_3669), .b(n_3660), .o(n_3780) );
na02f80 g740951 ( .a(n_39333), .b(n_39305), .o(n_40177) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_27_ ( .ck(newNet_3401), .d(n_27835), .o(delay_add_ln22_unr17_stage7_stallmux_q_27_) );
na02f80 g766826 ( .a(n_14341), .b(n_14344), .o(n_15572) );
no02f80 g767890 ( .a(n_13116), .b(n_13017), .o(n_13241) );
in01f80 g759986 ( .a(n_20441), .o(n_20442) );
no02f80 g762347 ( .a(n_45002), .b(n_18529), .o(n_18725) );
in01f80 FE_RC_2902_0 ( .a(n_19653), .o(FE_RN_1259_0) );
ao12f80 g773008 ( .a(n_8027), .b(n_7924), .c(FE_OCP_RBN3461_n_7886), .o(n_8046) );
in01f80 g772989 ( .a(n_7810), .o(n_8003) );
oa12f80 g747343 ( .a(n_32665), .b(FE_OCP_RBN2102_n_44962), .c(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n_32682) );
na02f80 g753180 ( .a(n_27207), .b(n_25757), .o(n_27456) );
no02f80 g778700 ( .a(FE_OCP_RBN2290_n_2438), .b(n_2056), .o(n_2652) );
na02f80 g764684 ( .a(n_16480), .b(n_16479), .o(n_16481) );
no02f80 g741516 ( .a(n_38703), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38723) );
no02f80 g737252 ( .a(n_42941), .b(n_43211), .o(n_42942) );
in01f80 newInst_2172 ( .a(newNet_372), .o(newNet_2172) );
na02f80 g764949 ( .a(n_15504), .b(n_15348), .o(n_15547) );
in01f80 g779270 ( .a(n_1725), .o(n_1786) );
in01f80 g782628 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n_44021) );
in01f80 fopt783424 ( .a(n_45024), .o(n_45026) );
na02f80 g751709 ( .a(n_28363), .b(n_28362), .o(n_28364) );
no02f80 g770987 ( .a(n_9456), .b(n_9461), .o(n_9463) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_21_ ( .ck(newNet_634), .d(n_46342), .o(delay_xor_ln21_unr9_stage4_stallmux_q_21_) );
in01f80 FE_OCP_RBC2666_n_35207 ( .a(n_35207), .o(FE_OCP_RBN2666_n_35207) );
na02f80 g779202 ( .a(n_1892), .b(n_1891), .o(n_2062) );
no02f80 g753483 ( .a(n_27540), .b(n_26868), .o(n_27541) );
in01f80 g742847 ( .a(n_37276), .o(n_37268) );
na02f80 g741662 ( .a(n_39040), .b(n_38553), .o(n_38554) );
na02f80 g736943 ( .a(FE_OCPN912_n_43022), .b(n_43135), .o(n_43320) );
na02f80 g779337 ( .a(n_1594), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .o(n_1666) );
in01f80 g781097 ( .a(mux_while_ln12_psv_q_8_), .o(n_275) );
ao12f80 g767923 ( .a(n_12712), .b(n_12711), .c(n_12710), .o(n_13119) );
ao12f80 g779485 ( .a(n_1990), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .o(n_2253) );
in01f80 g740130 ( .a(n_39846), .o(n_39867) );
na02f80 g767538 ( .a(n_13140), .b(n_13093), .o(n_14742) );
no02f80 g778575 ( .a(n_2476), .b(delay_add_ln22_unr2_stage2_stallmux_q_23_), .o(n_2499) );
no02f80 g739995 ( .a(n_40150), .b(n_40193), .o(n_40194) );
na02f80 g761924 ( .a(n_18634), .b(n_17856), .o(n_18672) );
oa12f80 g738969 ( .a(n_41162), .b(n_41161), .c(n_41160), .o(n_41211) );
no02f80 g776690 ( .a(n_3858), .b(n_3857), .o(n_3859) );
na02f80 g761335 ( .a(n_19903), .b(n_19648), .o(n_19904) );
na02f80 g775505 ( .a(n_5823), .b(n_5702), .o(n_5844) );
in01f80 FE_OCPC1427_n_13510 ( .a(n_13510), .o(FE_OCPN1427_n_13510) );
na02f80 g776486 ( .a(n_4450), .b(n_4174), .o(n_4585) );
oa12f80 g736379 ( .a(n_350), .b(n_43795), .c(FE_OFN2_n_43918), .o(n_43850) );
oa12f80 g761209 ( .a(FE_OCP_RBN2209_n_18280), .b(FE_OCP_RBN3827_n_18951), .c(n_19014), .o(n_19041) );
in01f80 FE_OCPC952_n_41540 ( .a(FE_OCPN951_n_41540), .o(FE_OCPN952_n_41540) );
oa12f80 g740114 ( .a(n_39799), .b(n_39798), .c(n_39797), .o(n_39847) );
na02f80 g780295 ( .a(n_1113), .b(n_956), .o(n_1021) );
no02f80 g773242 ( .a(n_8742), .b(n_7577), .o(n_7600) );
ao12f80 g747949 ( .a(n_33117), .b(n_33116), .c(n_33115), .o(n_33511) );
oa12f80 g765396 ( .a(n_15141), .b(n_15140), .c(n_15139), .o(n_15221) );
in01f80 g765995 ( .a(n_14809), .o(n_14810) );
in01f80 g756813 ( .a(n_24171), .o(n_23814) );
na02f80 g776566 ( .a(n_4355), .b(n_4210), .o(n_4407) );
no02f80 g771750 ( .a(n_10123), .b(n_10120), .o(n_10161) );
oa12f80 g780816 ( .a(n_476), .b(n_441), .c(n_403), .o(n_468) );
na02f80 FE_RC_164_0 ( .a(FE_RN_48_0), .b(FE_RN_49_0), .o(FE_RN_50_0) );
no02f80 g751549 ( .a(n_28450), .b(n_28449), .o(n_28468) );
na02f80 g738292 ( .a(n_41799), .b(n_41798), .o(n_41800) );
in01f80 FE_OCP_RBC1910_n_20545 ( .a(n_20545), .o(FE_OCP_RBN1910_n_20545) );
in01f80 FE_OCP_RBC2782_n_25997 ( .a(n_25997), .o(FE_OCP_RBN2782_n_25997) );
na02f80 g770691 ( .a(n_10241), .b(n_10185), .o(n_10322) );
in01f80 FE_RC_4025_0 ( .a(n_34516), .o(FE_RN_1748_0) );
in01f80 g764878 ( .a(n_15725), .o(n_15726) );
na02f80 g741950 ( .a(n_38090), .b(n_38041), .o(n_38091) );
in01f80 g762207 ( .a(n_18837), .o(n_18838) );
na02f80 g757881 ( .a(n_22979), .b(n_22879), .o(n_22980) );
in01f80 FE_OCP_RBC2267_n_2430 ( .a(n_2430), .o(FE_OCP_RBN2267_n_2430) );
no02f80 g760579 ( .a(n_19939), .b(n_19938), .o(n_19940) );
in01f80 g741618 ( .a(n_38690), .o(n_38647) );
na02f80 g770937 ( .a(n_9926), .b(n_9804), .o(n_10006) );
no02f80 g778545 ( .a(n_2307), .b(n_2348), .o(n_2349) );
no02f80 g749798 ( .a(n_31311), .b(n_31416), .o(n_31454) );
na02f80 g749675 ( .a(n_31638), .b(n_31637), .o(n_31639) );
in01f80 newInst_101 ( .a(newNet_100), .o(newNet_101) );
na02f80 g736623 ( .a(n_43118), .b(n_43054), .o(n_43240) );
in01f80 g736969 ( .a(n_43248), .o(n_43349) );
in01f80 g752443 ( .a(n_27800), .o(n_27767) );
no02f80 g763806 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n_17211) );
in01f80 g771280 ( .a(n_9617), .o(n_9618) );
na02f80 g751629 ( .a(n_28405), .b(delay_add_ln22_unr17_stage7_stallmux_q_12_), .o(n_28448) );
in01f80 g768864 ( .a(n_11958), .o(n_11874) );
na02f80 g762793 ( .a(n_17910), .b(n_17909), .o(n_17911) );
no02f80 g762652 ( .a(n_18038), .b(delay_add_ln22_unr11_stage5_stallmux_q_12_), .o(n_18067) );
no02f80 g739882 ( .a(n_40478), .b(n_40480), .o(n_40479) );
ao12f80 g769194 ( .a(n_11640), .b(FE_OCP_RBN1992_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .c(FE_OCPN1001_n_45660), .o(n_12218) );
in01f80 FE_RC_3384_0 ( .a(n_12940), .o(FE_RN_1467_0) );
in01f80 g772421 ( .a(n_8542), .o(n_8543) );
na02f80 FE_RC_2338_0 ( .a(n_18966), .b(n_18612), .o(FE_RN_895_0) );
no02f80 FE_RC_2516_0 ( .a(n_27536), .b(FE_OCP_RBN2920_n_31107), .o(FE_RN_1024_0) );
no02f80 g766024 ( .a(n_14971), .b(n_14742), .o(n_14743) );
in01f80 FE_RC_3724_0 ( .a(FE_RN_1639_0), .o(n_15079) );
in01f80 newInst_2330 ( .a(newNet_2329), .o(newNet_2330) );
in01f80 FE_OCPC1224_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCPN1224_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01f80 g765222 ( .a(n_15878), .o(n_15879) );
na02f80 FE_RC_2314_0 ( .a(n_35962), .b(n_35847), .o(FE_RN_879_0) );
in01f80 newInst_522 ( .a(newNet_520), .o(newNet_522) );
in01f80 g770000 ( .a(n_11012), .o(n_11039) );
na02f80 g748185 ( .a(n_31505), .b(n_31518), .o(n_31563) );
oa22f80 g774257 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .c(FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(n_6510), .o(n_6590) );
oa12f80 g773628 ( .a(n_7387), .b(n_7389), .c(n_7386), .o(n_7726) );
in01f80 g757517 ( .a(n_22829), .o(n_22800) );
in01f80 g754656 ( .a(n_27130), .o(n_30823) );
na02f80 g779188 ( .a(n_1869), .b(n_1631), .o(n_1870) );
no02f80 g768257 ( .a(n_12566), .b(n_11391), .o(n_12620) );
in01f80 FE_OCP_RBC3417_n_12739 ( .a(FE_OCP_RBN3415_n_12739), .o(FE_OCP_RBN3417_n_12739) );
oa12f80 g745355 ( .a(n_34210), .b(n_34226), .c(n_34209), .o(n_34262) );
na02f80 g751769 ( .a(FE_OCPN1038_n_28318), .b(n_28289), .o(n_28329) );
oa12f80 g759703 ( .a(n_21691), .b(n_21721), .c(n_21720), .o(n_21752) );
no03m80 g759686 ( .a(n_21779), .b(n_21749), .c(n_21778), .o(n_21780) );
in01f80 FE_RC_3854_0 ( .a(n_20123), .o(FE_RN_1682_0) );
in01f80 newInst_107 ( .a(newNet_106), .o(newNet_107) );
oa22f80 FE_RC_3920_0 ( .a(n_27459), .b(n_45619), .c(n_27460), .d(n_27715), .o(n_27804) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_16_ ( .ck(newNet_503), .d(n_22913), .o(delay_xor_ln22_unr15_stage6_stallmux_q_16_) );
ao12f80 g778747 ( .a(n_1470), .b(n_2200), .c(n_1423), .o(n_2212) );
no02f80 g747180 ( .a(n_32702), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(n_32719) );
in01f80 newInst_2310 ( .a(newNet_1831), .o(newNet_2310) );
in01f80 g780531 ( .a(n_1062), .o(n_1063) );
oa12f80 g771548 ( .a(n_8887), .b(n_8911), .c(n_8861), .o(n_9046) );
no02f80 g752177 ( .a(FE_OCPN877_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_7_), .o(n_28010) );
no02f80 g749964 ( .a(n_29780), .b(n_29826), .o(n_29847) );
in01f80 g763145 ( .a(n_17406), .o(n_17407) );
no02f80 g780410 ( .a(n_796), .b(n_795), .o(n_797) );
na02f80 g761468 ( .a(n_19787), .b(n_19986), .o(n_20254) );
na02f80 g769705 ( .a(n_11209), .b(n_11167), .o(n_11210) );
na02f80 g751985 ( .a(n_28793), .b(n_28856), .o(n_29105) );
ao12f80 g751847 ( .a(n_28093), .b(n_28192), .c(n_28142), .o(n_28234) );
ao22s80 FE_RC_702_0 ( .a(n_6579), .b(n_6638), .c(n_6656), .d(n_6637), .o(n_6835) );
na02f80 g762281 ( .a(FE_OFN750_n_45003), .b(n_18415), .o(n_18813) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_7_ ( .ck(newNet_996), .d(n_17291), .o(delay_xor_ln21_unr12_stage5_stallmux_q_7_) );
oa12f80 g762764 ( .a(n_17911), .b(n_17910), .c(n_17909), .o(n_19436) );
in01f80 g739988 ( .a(n_40121), .o(n_40157) );
in01f80 FE_OCPC1431_n_29504 ( .a(n_29504), .o(FE_OCPN1431_n_29504) );
in01f80 newInst_1687 ( .a(newNet_1686), .o(newNet_1687) );
in01f80 g753910 ( .a(n_27063), .o(n_27064) );
no02f80 g746851 ( .a(n_32924), .b(n_32898), .o(n_32899) );
in01f80 g740233 ( .a(n_39782), .o(n_39783) );
na02f80 g744082 ( .a(n_44222), .b(n_34978), .o(n_36190) );
na02f80 g742129 ( .a(n_37972), .b(n_37888), .o(n_38069) );
in01f80 FE_OCP_RBC2930_n_5221 ( .a(n_5221), .o(FE_OCP_RBN2930_n_5221) );
in01f80 g737170 ( .a(n_43030), .o(n_43046) );
in01f80 g743994 ( .a(n_36363), .o(n_36364) );
ao22s80 g784427 ( .a(n_36578), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_46239) );
in01f80 g757029 ( .a(n_23832), .o(n_23908) );
in01f80 g773978 ( .a(n_6908), .o(n_6909) );
in01f80 g763370 ( .a(n_17331), .o(n_17390) );
in01f80 newInst_671 ( .a(newNet_670), .o(newNet_671) );
ao22s80 g780436 ( .a(n_1203), .b(n_855), .c(FE_OFN795_n_45813), .d(n_764), .o(n_822) );
no02f80 g771886 ( .a(n_8838), .b(FE_OCPN917_n_46991), .o(n_8936) );
no02f80 g743518 ( .a(n_36581), .b(n_36750), .o(n_36582) );
in01f80 newInst_2492 ( .a(newNet_2491), .o(newNet_2492) );
in01f80 g776056 ( .a(n_5041), .o(n_5042) );
in01f80 g761471 ( .a(n_19761), .o(n_19762) );
oa22f80 g774263 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .c(FE_OCP_RBN1986_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(FE_OCP_RBN3251_delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(n_6654) );
no02f80 g748808 ( .a(n_32489), .b(n_32488), .o(n_33069) );
na02f80 g739775 ( .a(n_40422), .b(n_40040), .o(n_40466) );
in01f80 g761373 ( .a(n_19055), .o(n_19052) );
oa12f80 g778222 ( .a(n_2505), .b(n_2709), .c(n_2573), .o(n_2753) );
no02f80 g759228 ( .a(n_21339), .b(n_45070), .o(n_21309) );
no02f80 g756275 ( .a(n_24629), .b(n_24628), .o(n_24630) );
na02f80 g737755 ( .a(n_42363), .b(n_42310), .o(n_42355) );
oa12f80 g751030 ( .a(n_29825), .b(n_29824), .c(n_29823), .o(n_30166) );
no02f80 g775591 ( .a(n_5590), .b(n_5579), .o(n_5580) );
in01f80 newInst_1056 ( .a(newNet_1055), .o(newNet_1056) );
in01f80 fopt783665 ( .a(n_6649), .o(n_45314) );
no03m80 FE_RC_3224_0 ( .a(n_11535), .b(n_11484), .c(n_11483), .o(n_11726) );
in01f80 g754232 ( .a(FE_OCP_RBN2826_FE_RN_1573_0), .o(n_26014) );
in01f80 g775570 ( .a(n_5397), .o(n_5398) );
in01f80 g770355 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .o(n_10715) );
no02f80 g739428 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n_40774) );
in01f80 FE_OFC761_n_45813 ( .a(FE_OFN757_n_45813), .o(FE_OFN761_n_45813) );
no02f80 g776593 ( .a(n_4438), .b(n_4437), .o(n_4482) );
na02f80 g743834 ( .a(n_35833), .b(n_35708), .o(n_36335) );
na02f80 g770735 ( .a(n_10026), .b(n_10094), .o(n_10112) );
na02f80 g743250 ( .a(n_36931), .b(n_36884), .o(n_36906) );
in01f80 g743670 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n_36429) );
na02f80 g764931 ( .a(n_15357), .b(n_15113), .o(n_15394) );
oa12f80 g773573 ( .a(n_45861), .b(n_7427), .c(n_6877), .o(n_7474) );
na02f80 g775280 ( .a(n_5751), .b(n_5735), .o(n_5773) );
in01f80 newInst_3424 ( .a(newNet_3423), .o(newNet_3424) );
in01f80 newInst_3376 ( .a(newNet_3375), .o(newNet_3376) );
no02f80 g755864 ( .a(n_25033), .b(n_25032), .o(n_25034) );
no02f80 g739923 ( .a(n_40336), .b(n_40120), .o(n_40337) );
in01f80 newInst_900 ( .a(newNet_899), .o(newNet_900) );
in01f80 FE_RC_1276_0 ( .a(n_2280), .o(FE_RN_375_0) );
in01f80 g778549 ( .a(n_2374), .o(n_2375) );
in01f80 g766662 ( .a(n_13884), .o(n_13885) );
no03m80 FE_RC_1723_0 ( .a(FE_OCPN1776_n_18263), .b(n_18317), .c(n_18602), .o(n_18652) );
ms00f80 sin_out_reg_25_ ( .ck(newNet_45), .d(n_43913), .o(sin_out_25) );
na02f80 g755883 ( .a(n_25003), .b(n_25002), .o(n_25004) );
na02f80 g736690 ( .a(n_43278), .b(n_43315), .o(n_43331) );
no02f80 g772736 ( .a(FE_RN_347_0), .b(n_8213), .o(n_8237) );
na02f80 g749309 ( .a(n_30655), .b(n_30371), .o(n_30678) );
in01f80 g780506 ( .a(n_987), .o(n_988) );
na02f80 g778127 ( .a(n_2872), .b(n_3361), .o(n_2890) );
in01f80 g778317 ( .a(n_2927), .o(n_2976) );
na02f80 g766026 ( .a(n_14643), .b(n_14600), .o(n_14694) );
no02f80 g762971 ( .a(n_17984), .b(n_17983), .o(n_17985) );
oa22f80 FE_RC_2849_0 ( .a(n_24920), .b(FE_RN_705_0), .c(n_24919), .d(FE_RN_706_0), .o(n_25074) );
in01f80 newInst_3603 ( .a(newNet_3602), .o(newNet_3603) );
na02f80 g770222 ( .a(n_10869), .b(n_10841), .o(n_10842) );
oa22f80 FE_RC_3834_0 ( .a(n_20434), .b(n_20799), .c(n_20460), .d(n_20819), .o(n_20941) );
oa12f80 g742622 ( .a(n_37523), .b(n_37522), .c(n_37521), .o(n_37587) );
ao12f80 g740904 ( .a(n_39203), .b(n_39088), .c(n_39251), .o(n_39288) );
in01f80 g744865 ( .a(n_35132), .o(n_35194) );
in01f80 g767919 ( .a(n_12763), .o(n_12764) );
no02f80 g738920 ( .a(n_41267), .b(n_41266), .o(n_41268) );
ao22s80 g762671 ( .a(n_17997), .b(n_17941), .c(n_17943), .d(n_17940), .o(n_19562) );
na02f80 g766435 ( .a(n_14100), .b(n_13122), .o(n_14163) );
in01f80 g752465 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .o(n_27719) );
no02f80 FE_RC_413_0 ( .a(FE_RN_122_0), .b(n_14242), .o(n_45521) );
na02f80 g758838 ( .a(n_21477), .b(n_21331), .o(n_21511) );
no02f80 g740420 ( .a(FE_OCP_RBN3022_n_39942), .b(FE_OCP_RBN2864_n_39523), .o(n_40097) );
in01f80 newInst_3352 ( .a(newNet_3351), .o(newNet_3352) );
na02f80 g777300 ( .a(n_4606), .b(n_3264), .o(n_4745) );
na02f80 g742391 ( .a(n_37736), .b(n_37692), .o(n_37769) );
no02f80 g755033 ( .a(n_25102), .b(n_23887), .o(n_25155) );
no02f80 g751414 ( .a(n_28609), .b(n_28608), .o(n_28893) );
oa22f80 g739824 ( .a(n_40261), .b(n_40289), .c(n_40262), .d(n_40290), .o(n_40404) );
in01f80 newInst_3128 ( .a(newNet_3127), .o(newNet_3128) );
in01f80 g763968 ( .a(n_16638), .o(n_16639) );
in01f80 g741833 ( .a(n_38321), .o(n_38322) );
na02f80 g751211 ( .a(n_28791), .b(n_28779), .o(n_28780) );
ao12f80 g780355 ( .a(n_877), .b(n_1155), .c(n_876), .o(n_947) );
na02f80 g775971 ( .a(n_5101), .b(n_3625), .o(n_5152) );
no02f80 g744540 ( .a(n_35387), .b(n_35284), .o(n_35413) );
no02f80 g741522 ( .a(n_38667), .b(n_38629), .o(n_38709) );
na02f80 g756734 ( .a(n_23397), .b(n_23287), .o(n_23431) );
oa22f80 g739670 ( .a(n_40517), .b(n_40114), .c(n_40518), .d(n_40115), .o(n_40553) );
na02f80 g769277 ( .a(n_11627), .b(FE_OCP_RBN3006_n_11087), .o(n_11619) );
no02f80 g760387 ( .a(n_20149), .b(n_18140), .o(n_20150) );
na02f80 g776568 ( .a(n_4225), .b(n_4219), .o(n_4393) );
no02f80 g763421 ( .a(n_16942), .b(n_16903), .o(n_17071) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_19_ ( .ck(newNet_177), .d(n_46357), .o(delay_xor_ln22_unr9_stage4_stallmux_q_19_) );
in01f80 newInst_3321 ( .a(newNet_3320), .o(newNet_3321) );
na02f80 g763191 ( .a(n_17401), .b(FE_RN_25_0), .o(n_17582) );
in01f80 g747151 ( .a(n_32870), .o(n_32871) );
ao12f80 g738933 ( .a(n_41167), .b(n_41166), .c(n_41165), .o(n_41217) );
no02f80 g753202 ( .a(n_27207), .b(n_25999), .o(n_27390) );
in01f80 g753291 ( .a(n_27677), .o(n_27678) );
na02f80 g749765 ( .a(n_31344), .b(n_31312), .o(n_31345) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_6_ ( .ck(newNet_2343), .d(n_35557), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_9_ ( .ck(newNet_1675), .d(n_22055), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_) );
in01f80 g756034 ( .a(n_24929), .o(n_24930) );
in01f80 g768359 ( .a(n_12554), .o(n_12555) );
na02f80 g753977 ( .a(FE_OCP_RBN2892_n_26152), .b(n_26048), .o(n_26213) );
na02f80 g758574 ( .a(n_21905), .b(n_21925), .o(n_21938) );
in01f80 newInst_1797 ( .a(newNet_1796), .o(newNet_1797) );
no02f80 g773646 ( .a(n_7288), .b(delay_add_ln22_unr5_stage3_stallmux_q_18_), .o(n_7307) );
in01f80 g756223 ( .a(n_25124), .o(n_24844) );
in01f80 g752667 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_), .o(n_28452) );
in01f80 FE_OCP_RBC3339_n_44610 ( .a(n_44610), .o(FE_OCP_RBN3339_n_44610) );
no02f80 g761721 ( .a(n_18647), .b(n_18214), .o(n_18653) );
in01f80 g776526 ( .a(n_4154), .o(n_4177) );
na02f80 g755373 ( .a(n_24829), .b(n_24692), .o(n_24895) );
no02f80 g747113 ( .a(n_32745), .b(n_32761), .o(n_32822) );
in01f80 g765667 ( .a(n_15170), .o(n_15171) );
in01f80 FE_OCP_DRV_C1553_n_19314 ( .a(n_19314), .o(FE_OCP_DRV_N1553_n_19314) );
ao22s80 FE_RC_1681_0 ( .a(n_13575), .b(n_12794), .c(n_13576), .d(n_12793), .o(n_13661) );
ao12f80 g761771 ( .a(n_18885), .b(n_19191), .c(n_18809), .o(n_19296) );
no02f80 g765564 ( .a(n_15142), .b(n_14317), .o(n_15806) );
ao12f80 g751350 ( .a(n_29411), .b(n_29410), .c(n_29409), .o(n_29935) );
na02f80 g748423 ( .a(n_31476), .b(n_30906), .o(n_31657) );
in01f80 FE_OCP_RBC2749_n_9629 ( .a(n_9629), .o(FE_OCP_RBN2749_n_9629) );
oa22f80 FE_RC_1485_0 ( .a(n_27499), .b(n_27605), .c(n_27498), .d(n_27604), .o(n_27686) );
in01f80 g765856 ( .a(n_14884), .o(n_14885) );
no02f80 g781160 ( .a(n_198), .b(n_264), .o(n_204) );
na02f80 g757995 ( .a(n_22698), .b(n_22621), .o(n_22765) );
in01f80 g767427 ( .a(n_13398), .o(n_13399) );
na02f80 g762242 ( .a(n_18451), .b(n_17427), .o(n_18501) );
in01f80 g760125 ( .a(n_20495), .o(n_20496) );
ao22s80 FE_RC_3166_0 ( .a(n_25935), .b(n_45329), .c(n_25919), .d(n_25964), .o(n_26085) );
in01f80 g739331 ( .a(n_40734), .o(n_40788) );
na02f80 g755333 ( .a(n_24810), .b(n_24829), .o(n_24881) );
no02f80 g744555 ( .a(n_35352), .b(n_35274), .o(n_35384) );
oa12f80 g739366 ( .a(n_40717), .b(n_44775), .c(n_40299), .o(n_41054) );
no02f80 g744812 ( .a(n_35118), .b(n_35080), .o(n_35139) );
na02f80 g739307 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n_41009) );
in01f80 g771683 ( .a(n_9238), .o(n_9239) );
in01f80 g741104 ( .a(n_39207), .o(n_39208) );
in01f80 g757467 ( .a(n_23954), .o(n_23979) );
in01f80 g743947 ( .a(n_36199), .o(n_36149) );
in01f80 newInst_1377 ( .a(newNet_1026), .o(newNet_1377) );
na02f80 g763402 ( .a(n_16975), .b(n_16084), .o(n_17217) );
in01f80 FE_OCPC1504_n_47257 ( .a(FE_OCPN1503_n_47257), .o(FE_OCPN1504_n_47257) );
no02f80 FE_RC_3000_0 ( .a(n_10542), .b(FE_OCP_RBN2870_n_10480), .o(FE_RN_1313_0) );
in01f80 g742665 ( .a(n_37547), .o(n_38315) );
na02f80 g775083 ( .a(n_5987), .b(n_5710), .o(n_6019) );
in01f80 g766783 ( .a(n_13751), .o(n_13750) );
na02f80 g748912 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .o(n_32457) );
ao12f80 g765375 ( .a(n_15920), .b(n_15874), .c(n_15869), .o(n_16302) );
oa22f80 FE_RC_833_0 ( .a(n_24048), .b(n_24468), .c(n_24049), .d(n_24467), .o(n_24621) );
in01f80 g780476 ( .a(n_1098), .o(n_1099) );
na02f80 g766284 ( .a(n_14245), .b(n_14155), .o(n_14246) );
in01f80 g744071 ( .a(n_35948), .o(n_36035) );
ao12f80 g772271 ( .a(n_8737), .b(n_8736), .c(n_8735), .o(n_8810) );
in01f80 g747373 ( .a(n_32600), .o(n_32439) );
in01f80 g739661 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_28_), .o(n_40590) );
in01f80 g737355 ( .a(n_42864), .o(n_42879) );
na02f80 g770171 ( .a(n_10754), .b(n_10724), .o(n_10803) );
in01f80 g775299 ( .a(n_5672), .o(n_5691) );
in01f80 g744992 ( .a(n_34990), .o(n_34991) );
na02f80 g764925 ( .a(n_15584), .b(n_15537), .o(n_15614) );
in01f80 g739918 ( .a(n_40260), .o(n_40297) );
in01f80 g769936 ( .a(n_11131), .o(n_11152) );
no02f80 g749065 ( .a(n_30996), .b(n_30995), .o(n_30997) );
no02f80 g740375 ( .a(n_39942), .b(n_39832), .o(n_39973) );
no02f80 g738733 ( .a(n_41483), .b(n_41613), .o(n_41912) );
in01f80 FE_OCP_RBC3430_n_13245 ( .a(n_13245), .o(FE_OCP_RBN3430_n_13245) );
in01f80 fopt782885 ( .a(n_22625), .o(n_44322) );
no02f80 g764839 ( .a(n_16139), .b(n_15744), .o(n_16211) );
in01f80 g776454 ( .a(n_4753), .o(n_4754) );
in01f80 g761955 ( .a(FE_OFN814_n_18287), .o(n_18288) );
na02f80 g777328 ( .a(n_3604), .b(n_3721), .o(n_3768) );
in01f80 newInst_3725 ( .a(newNet_3127), .o(newNet_3725) );
oa12f80 g754261 ( .a(n_26945), .b(n_26944), .c(n_26943), .o(n_27000) );
na02f80 g746930 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .o(n_32915) );
na02f80 g748210 ( .a(n_32019), .b(n_32051), .o(n_32120) );
in01f80 fopt783367 ( .a(n_38830), .o(n_44955) );
ao12f80 g751921 ( .a(n_29002), .b(n_28919), .c(n_28984), .o(n_29692) );
oa12f80 g738176 ( .a(n_41775), .b(n_41985), .c(n_41667), .o(n_42018) );
in01f80 g780591 ( .a(n_925), .o(n_898) );
oa12f80 g744448 ( .a(n_35450), .b(n_35449), .c(n_35460), .o(n_35474) );
na02f80 g758608 ( .a(n_21849), .b(n_21708), .o(n_21850) );
in01f80 g748029 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_11_), .o(n_31855) );
na02f80 FE_RC_1235_0 ( .a(FE_RN_369_0), .b(FE_RN_370_0), .o(FE_RN_371_0) );
in01f80 fopt782681 ( .a(n_44083), .o(n_44066) );
na02f80 g771333 ( .a(n_9295), .b(n_9254), .o(n_9450) );
oa12f80 g754757 ( .a(n_25176), .b(n_25248), .c(n_25146), .o(n_25365) );
oa22f80 FE_RC_1582_0 ( .a(n_4789), .b(n_5400), .c(n_4790), .d(n_5364), .o(n_5508) );
ao12f80 g756379 ( .a(n_23542), .b(n_23826), .c(n_23571), .o(n_23859) );
na02f80 g743087 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .o(n_37051) );
ms00f80 mux_while_ln12_psv_q_reg_7_ ( .ck(newNet_101), .d(n_243), .o(mux_while_ln12_psv_q_7_) );
oa12f80 g749041 ( .a(n_31543), .b(n_32231), .c(n_31541), .o(n_32292) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_16_ ( .ck(newNet_3243), .d(n_36407), .o(delay_add_ln22_unr23_stage9_stallmux_q_16_) );
no02f80 g773729 ( .a(n_7246), .b(n_7245), .o(n_7247) );
na02f80 g772994 ( .a(n_45846), .b(n_45871), .o(n_7773) );
no02f80 g756778 ( .a(n_23814), .b(n_23869), .o(n_23870) );
in01f80 g737486 ( .a(n_43061), .o(n_42730) );
no02f80 g751185 ( .a(n_29837), .b(n_29838), .o(n_29881) );
in01f80 g744962 ( .a(FE_OCP_RBN2712_n_35075), .o(n_35090) );
in01f80 g739853 ( .a(n_40429), .o(n_40430) );
no02f80 g749441 ( .a(n_30639), .b(n_30620), .o(n_30723) );
na02f80 g768061 ( .a(n_12790), .b(n_12789), .o(n_12841) );
in01f80 g755354 ( .a(n_24887), .o(n_24859) );
no02f80 g769818 ( .a(n_11165), .b(n_44453), .o(n_11217) );
na02f80 g759549 ( .a(n_20846), .b(FE_OCPN1444_n_45050), .o(n_20912) );
no02f80 g753516 ( .a(n_26804), .b(n_23564), .o(n_26824) );
ms00f80 cos_out_reg_2_ ( .ck(newNet_2), .d(n_43381), .o(cos_out_2) );
ao12f80 g764207 ( .a(n_16210), .b(n_16798), .c(n_15929), .o(n_16820) );
in01f80 g741282 ( .a(n_38942), .o(n_38978) );
na02f80 g758313 ( .a(n_22249), .b(n_21278), .o(n_22330) );
na02f80 g772450 ( .a(n_8490), .b(n_7851), .o(n_8561) );
na02f80 g769174 ( .a(n_11864), .b(n_11960), .o(n_11961) );
no02f80 g738685 ( .a(n_41537), .b(n_41212), .o(n_41614) );
no02f80 g764487 ( .a(n_16122), .b(n_14524), .o(n_16158) );
in01f80 g751785 ( .a(FE_OCPN1036_n_28288), .o(n_28289) );
no02f80 g757560 ( .a(n_22768), .b(n_44061), .o(n_22821) );
na02f80 g748528 ( .a(n_31697), .b(FE_RN_172_0), .o(n_31713) );
na02f80 g762621 ( .a(n_18070), .b(n_18041), .o(n_18042) );
no02f80 FE_RC_2393_0 ( .a(FE_RN_937_0), .b(FE_RN_939_0), .o(n_42790) );
in01f80 g744611 ( .a(n_36623), .o(n_36642) );
na02f80 g763523 ( .a(FE_OCP_RBN1210_n_16814), .b(n_16842), .o(n_16902) );
no02f80 g740831 ( .a(n_39219), .b(n_39302), .o(n_39383) );
na02f80 g763156 ( .a(n_17819), .b(n_17818), .o(n_17820) );
in01f80 newInst_2879 ( .a(newNet_2423), .o(newNet_2879) );
in01f80 g764856 ( .a(n_15755), .o(n_15756) );
oa12f80 g736399 ( .a(n_325), .b(n_43757), .c(FE_OFN3_n_43918), .o(n_43802) );
in01f80 g737554 ( .a(n_42590), .o(n_42591) );
in01f80 g770241 ( .a(n_10925), .o(n_10926) );
in01f80 FE_RC_3657_0 ( .a(FE_RN_1605_0), .o(n_21742) );
no02f80 g742020 ( .a(n_37911), .b(n_44872), .o(n_38042) );
na02f80 g754908 ( .a(n_25542), .b(n_24612), .o(n_25624) );
in01f80 g747130 ( .a(n_32983), .o(n_32984) );
in01f80 g764322 ( .a(n_16722), .o(n_16723) );
no02f80 g738232 ( .a(n_41897), .b(n_41754), .o(n_41939) );
in01f80 FE_RC_4_0 ( .a(n_1705), .o(FE_RN_0_0) );
na02f80 g755690 ( .a(n_24461), .b(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24497) );
in01f80 g767912 ( .a(n_13038), .o(n_13039) );
na02f80 g771259 ( .a(FE_RN_1125_0), .b(n_9372), .o(n_9452) );
in01f80 newInst_2810 ( .a(newNet_2809), .o(newNet_2810) );
oa12f80 g747703 ( .a(n_33372), .b(n_33418), .c(n_33169), .o(n_33419) );
in01f80 FE_OCP_RBC3831_n_19204 ( .a(FE_OCP_RBN3829_n_19204), .o(FE_OCP_RBN3831_n_19204) );
in01f80 newInst_276 ( .a(newNet_156), .o(newNet_276) );
na02f80 g754329 ( .a(n_25843), .b(n_25502), .o(n_25875) );
in01f80 g752565 ( .a(n_27661), .o(n_27681) );
na02f80 g746951 ( .a(n_32857), .b(n_32912), .o(n_32939) );
ao22s80 FE_RC_1687_0 ( .a(n_33664), .b(FE_OCP_RBN1356_n_44259), .c(n_44259), .d(FE_OCP_RBN3431_n_33664), .o(n_33780) );
no02f80 g781245 ( .a(n_111), .b(n_53), .o(n_228) );
in01f80 FE_OCPC1758_n_33213 ( .a(FE_OCPN1757_n_33213), .o(FE_OCPN1758_n_33213) );
ao12f80 g755454 ( .a(FE_OCPN1474_n_24624), .b(n_24602), .c(n_24601), .o(n_24659) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_19_ ( .ck(newNet_347), .d(n_1351), .o(delay_xor_ln22_unr3_stage2_stallmux_q_19_) );
oa22f80 g763872 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .c(n_16618), .d(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17983) );
in01f80 newInst_2250 ( .a(newNet_2249), .o(newNet_2250) );
na02f80 g754092 ( .a(n_26098), .b(n_23317), .o(n_26178) );
in01f80 g769950 ( .a(n_10880), .o(n_10881) );
in01f80 g765258 ( .a(n_15266), .o(n_15267) );
in01f80 FE_OFC799_n_46285 ( .a(n_46285), .o(FE_OFN799_n_46285) );
in01f80 g754677 ( .a(FE_OCPN1410_n_27014), .o(n_30790) );
in01f80 FE_OCP_RBC2510_n_13896 ( .a(FE_OCP_RBN2508_n_13896), .o(FE_OCP_RBN2510_n_13896) );
in01f80 g768041 ( .a(n_12782), .o(n_12759) );
na02f80 g776688 ( .a(n_3858), .b(n_2975), .o(n_3860) );
in01f80 FE_OCPC3759_n_2346 ( .a(FE_OCPN3758_n_2346), .o(FE_OCPN3759_n_2346) );
in01f80 FE_RC_848_0 ( .a(FE_OCPN1406_n_25859), .o(FE_RN_252_0) );
in01f80 g746847 ( .a(n_33301), .o(n_33302) );
na02f80 g756864 ( .a(n_23751), .b(n_23750), .o(n_23752) );
na03f80 g776383 ( .a(n_4547), .b(n_4386), .c(n_4366), .o(n_4548) );
oa12f80 g757062 ( .a(n_23803), .b(n_23979), .c(n_23978), .o(n_23980) );
in01f80 FE_RC_3850_0 ( .a(n_19645), .o(FE_RN_1680_0) );
na02f80 g763008 ( .a(n_17590), .b(n_17589), .o(n_17672) );
ao12f80 g743712 ( .a(n_35744), .b(n_36372), .c(n_36303), .o(n_36390) );
no02f80 g779553 ( .a(FE_OCP_RBN3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_2_), .o(n_1435) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_5_ ( .ck(newNet_3281), .d(n_31267), .o(delay_add_ln22_unr20_stage8_stallmux_q_5_) );
in01f80 g774951 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_), .o(n_7424) );
in01f80 g770510 ( .a(n_10556), .o(n_10557) );
in01f80 FE_OCP_RBC3250_delay_xor_ln22_unr6_stage3_stallmux_q_0_ ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(FE_OCP_RBN3250_delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
no02f80 g778000 ( .a(n_3066), .b(n_2828), .o(n_3086) );
in01f80 g770911 ( .a(n_9855), .o(n_9754) );
in01f80 g763223 ( .a(n_17785), .o(n_17786) );
in01f80 FE_OCP_RBC2611_n_3718 ( .a(n_3718), .o(FE_OCP_RBN2611_n_3718) );
na03f80 g766903 ( .a(n_14213), .b(n_14077), .c(n_14212), .o(n_14214) );
na02f80 g763900 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .o(n_17421) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_9_ ( .ck(newNet_2230), .d(n_40420), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_) );
no02f80 g740897 ( .a(n_39167), .b(n_38916), .o(n_39222) );
in01f80 FE_OCP_RBC2212_n_37720 ( .a(n_37720), .o(FE_OCP_RBN2212_n_37720) );
in01f80 g756618 ( .a(n_23972), .o(n_23885) );
na02f80 g777374 ( .a(n_4219), .b(n_4207), .o(n_4261) );
no02f80 g770930 ( .a(n_9580), .b(n_9456), .o(n_9671) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_5_ ( .ck(newNet_781), .d(n_1320), .o(delay_xor_ln21_unr3_stage2_stallmux_q_5_) );
in01f80 g766033 ( .a(n_14750), .o(n_14692) );
in01f80 g745086 ( .a(n_34966), .o(n_34967) );
no02f80 FE_RC_857_0 ( .a(FE_RN_255_0), .b(FE_RN_256_0), .o(FE_RN_257_0) );
in01f80 g749487 ( .a(n_31888), .o(n_31911) );
na02f80 g763090 ( .a(n_17411), .b(n_17448), .o(n_17590) );
in01f80 FE_RC_182_0 ( .a(n_353), .o(FE_RN_60_0) );
in01f80 fopt783111 ( .a(n_44592), .o(n_44575) );
oa22f80 g784418 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .c(n_36784), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46230) );
ao12f80 g756909 ( .a(n_23208), .b(n_23346), .c(n_23216), .o(n_23365) );
na02f80 FE_RC_2415_0 ( .a(FE_RN_953_0), .b(n_7417), .o(FE_RN_954_0) );
in01f80 FE_OCP_RBC2940_n_26276 ( .a(n_26276), .o(FE_OCP_RBN2940_n_26276) );
na02f80 g760234 ( .a(FE_OCP_RBN3613_n_20249), .b(FE_OCP_RBN3829_n_19204), .o(n_20391) );
in01f80 newInst_1029 ( .a(newNet_85), .o(newNet_1029) );
no02f80 g757896 ( .a(n_22353), .b(FE_OCPN3166_n_44267), .o(n_22420) );
no02f80 FE_RC_2710_0 ( .a(n_12945), .b(FE_RN_1140_0), .o(FE_RN_1141_0) );
no02f80 g776440 ( .a(n_4485), .b(n_3563), .o(n_4765) );
oa12f80 g749743 ( .a(FE_OCP_RBN3019_n_31117), .b(n_31324), .c(n_30920), .o(n_31325) );
in01f80 g779143 ( .a(n_1958), .o(n_1964) );
no02f80 g764480 ( .a(n_16009), .b(n_16080), .o(n_16172) );
na02f80 g750920 ( .a(n_28952), .b(n_28726), .o(n_28977) );
in01f80 newInst_2615 ( .a(newNet_776), .o(newNet_2615) );
na02f80 g775723 ( .a(n_5365), .b(n_4069), .o(n_5402) );
no02f80 g750450 ( .a(n_29552), .b(n_29575), .o(n_29645) );
in01f80 newInst_554 ( .a(newNet_553), .o(newNet_554) );
in01f80 FE_OCP_RBC1340_n_19077 ( .a(n_19077), .o(FE_OCP_RBN1340_n_19077) );
na02f80 g755433 ( .a(n_24655), .b(n_24652), .o(n_24699) );
no02f80 g752906 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .o(n_27903) );
oa12f80 g761527 ( .a(n_19546), .b(n_19545), .c(n_19544), .o(n_19848) );
no02f80 g749540 ( .a(n_31780), .b(n_31510), .o(n_31781) );
na02f80 g771777 ( .a(n_9157), .b(FE_OCP_RBN2606_FE_OCPN899_n_44593), .o(n_9327) );
in01f80 g777852 ( .a(n_3363), .o(n_3364) );
no02f80 FE_RC_3106_0 ( .a(FE_RN_1373_0), .b(FE_OCP_RBN3083_n_31819), .o(n_31903) );
in01f80 g764708 ( .a(n_15901), .o(n_15983) );
ao12f80 g772335 ( .a(n_8082), .b(n_8656), .c(n_7916), .o(n_8736) );
na02f80 g760554 ( .a(n_19843), .b(n_19867), .o(n_19942) );
ao12f80 g768978 ( .a(n_12278), .b(n_45659), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n_12706) );
no02f80 FE_RC_2189_0 ( .a(FE_RN_783_0), .b(n_21660), .o(n_21811) );
ao12f80 g774381 ( .a(n_6764), .b(n_6624), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n_7602) );
no02f80 g760694 ( .a(n_19633), .b(n_19418), .o(n_19703) );
ao22s80 g739594 ( .a(FE_OCP_RBN3338_n_44610), .b(FE_OCP_RBN3357_delay_xor_ln22_unr28_stage10_stallmux_q_0_), .c(n_44610), .d(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n_40616) );
no02f80 g767516 ( .a(n_13184), .b(n_13224), .o(n_13394) );
in01f80 g765646 ( .a(n_15038), .o(n_15039) );
oa12f80 g768296 ( .a(n_12608), .b(n_12607), .c(n_12606), .o(n_12673) );
oa22f80 FE_RC_1314_0 ( .a(n_10521), .b(n_10946), .c(n_10522), .d(n_10947), .o(n_11087) );
no02f80 g771230 ( .a(n_9657), .b(n_9405), .o(n_9702) );
in01f80 g763160 ( .a(n_17345), .o(n_17346) );
no02f80 g758014 ( .a(n_47278), .b(n_22198), .o(n_22336) );
in01f80 g748942 ( .a(n_31230), .o(n_31231) );
in01f80 FE_OCP_RBC2499_n_8835 ( .a(FE_OCP_RBN2498_n_8835), .o(FE_OCP_RBN2499_n_8835) );
na02f80 g780375 ( .a(n_856), .b(n_778), .o(n_903) );
in01f80 FE_OCP_RBC3373_n_6745 ( .a(FE_OCP_RBN2127_n_6745), .o(FE_OCP_RBN3373_n_6745) );
ao22s80 g778224 ( .a(FE_OCP_RBN2321_n_2638), .b(n_2155), .c(n_2638), .d(n_2154), .o(n_3390) );
na02f80 g773769 ( .a(n_7218), .b(n_6999), .o(n_7246) );
no02f80 g746126 ( .a(n_33918), .b(n_33917), .o(n_33919) );
in01f80 g741937 ( .a(n_38067), .o(n_38068) );
na02f80 g769634 ( .a(n_11299), .b(n_11246), .o(n_11329) );
in01f80 FE_OCP_RBC3696_n_5284 ( .a(n_5284), .o(FE_OCP_RBN3696_n_5284) );
in01f80 g759773 ( .a(n_21375), .o(n_21376) );
in01f80 newInst_2798 ( .a(newNet_582), .o(newNet_2798) );
in01f80 g771922 ( .a(n_8995), .o(n_9032) );
no02f80 g757943 ( .a(n_22029), .b(FE_OCPN1398_n_21973), .o(n_22087) );
no02f80 g751538 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_24_), .o(n_28645) );
na02f80 FE_RC_909_0 ( .a(n_11518), .b(n_45748), .o(FE_RN_268_0) );
in01f80 FE_RC_3376_0 ( .a(FE_RN_1465_0), .o(FE_RN_1464_0) );
in01f80 g743796 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_9_), .o(n_36151) );
in01f80 newInst_1341 ( .a(newNet_1340), .o(newNet_1341) );
no02f80 g748417 ( .a(n_31466), .b(n_30814), .o(n_31594) );
in01f80 g737086 ( .a(n_43017), .o(n_43018) );
in01f80 newInst_612 ( .a(newNet_598), .o(newNet_612) );
na02f80 g754389 ( .a(n_25705), .b(n_25511), .o(n_25783) );
no02f80 g738333 ( .a(n_41596), .b(n_41552), .o(n_41553) );
in01f80 newInst_2588 ( .a(newNet_2587), .o(newNet_2588) );
na02f80 g748951 ( .a(n_31131), .b(n_31105), .o(n_31194) );
in01f80 newInst_733 ( .a(newNet_732), .o(newNet_733) );
na02f80 g767557 ( .a(n_13053), .b(n_12796), .o(n_13140) );
ao12f80 g757278 ( .a(n_23224), .b(n_23223), .c(n_23222), .o(n_23278) );
na02f80 FE_RC_3560_0 ( .a(n_13436), .b(n_13388), .o(FE_RN_1546_0) );
in01f80 g752201 ( .a(n_28635), .o(n_28636) );
na02f80 g752970 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n_28256) );
no02f80 g743034 ( .a(n_37426), .b(n_37099), .o(n_37151) );
na02f80 g755469 ( .a(n_25261), .b(n_25112), .o(n_25347) );
in01f80 newInst_2738 ( .a(newNet_2737), .o(newNet_2738) );
ao12f80 g765177 ( .a(n_15340), .b(n_15296), .c(n_15256), .o(n_15526) );
in01f80 g738025 ( .a(n_42166), .o(n_42173) );
in01f80 newInst_2597 ( .a(newNet_1383), .o(newNet_2597) );
in01f80 newInst_759 ( .a(newNet_534), .o(newNet_759) );
in01f80 g763656 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .o(n_16807) );
in01f80 g763665 ( .a(n_16857), .o(n_17437) );
in01f80 g779005 ( .a(n_2192), .o(n_2193) );
no02f80 g756791 ( .a(n_23421), .b(n_23440), .o(n_23513) );
in01f80 g771971 ( .a(n_9953), .o(n_9954) );
in01f80 FE_OCP_RBC1142_n_25816 ( .a(FE_OCP_RBN1141_n_25816), .o(FE_OCP_RBN1142_n_25816) );
in01f80 newInst_1539 ( .a(newNet_1161), .o(newNet_1539) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_4_ ( .ck(newNet_3590), .d(n_15489), .o(delay_add_ln22_unr11_stage5_stallmux_q_4_) );
oa12f80 g782642 ( .a(n_37916), .b(n_37891), .c(n_37835), .o(n_44036) );
in01f80 newInst_2926 ( .a(newNet_1323), .o(newNet_2926) );
no02f80 g746736 ( .a(n_32965), .b(n_32999), .o(n_33022) );
oa22f80 g746570 ( .a(n_34810), .b(n_33993), .c(n_34666), .d(n_34643), .o(n_35245) );
oa22f80 FE_RC_1253_0 ( .a(n_23787), .b(n_24148), .c(n_23786), .d(n_24166), .o(n_24254) );
no02f80 g747623 ( .a(n_33761), .b(n_33812), .o(n_33813) );
in01f80 FE_OCPC855_n_20367 ( .a(n_20367), .o(FE_OCPN855_n_20367) );
no02f80 g780400 ( .a(n_802), .b(n_767), .o(n_789) );
in01f80 g743265 ( .a(n_36790), .o(n_36791) );
in01f80 g776953 ( .a(n_4173), .o(n_4174) );
no02f80 g757049 ( .a(n_23700), .b(n_23698), .o(n_24037) );
in01f80 FE_RC_4153_0 ( .a(n_23134), .o(FE_RN_1807_0) );
no02f80 g771949 ( .a(n_44464), .b(n_9913), .o(n_10039) );
na02f80 g779613 ( .a(n_1516), .b(n_1507), .o(n_2131) );
in01f80 g770100 ( .a(n_10797), .o(n_10802) );
no02f80 g756019 ( .a(n_25026), .b(n_25136), .o(n_25189) );
no02f80 g766158 ( .a(n_14483), .b(n_14371), .o(n_14552) );
in01f80 g747248 ( .a(n_32815), .o(n_32816) );
no02f80 g751157 ( .a(n_29932), .b(n_29768), .o(n_30091) );
in01f80 newInst_2609 ( .a(newNet_2608), .o(newNet_2609) );
in01f80 newInst_3015 ( .a(newNet_3014), .o(newNet_3015) );
in01f80 g769343 ( .a(n_11544), .o(n_11630) );
na02f80 g762279 ( .a(n_18534), .b(n_18658), .o(n_19193) );
in01f80 FE_OCP_RBC2505_n_13896 ( .a(FE_OCP_RBN2500_n_13896), .o(FE_OCP_RBN2505_n_13896) );
in01f80 fopt783514 ( .a(FE_OCP_RBN3409_n_45120), .o(n_45118) );
na02f80 g778161 ( .a(n_2801), .b(n_2193), .o(n_2802) );
in01f80 g743483 ( .a(n_36651), .o(n_36628) );
in01f80 FE_OCP_RBC3697_n_35543 ( .a(n_35543), .o(FE_OCP_RBN3697_n_35543) );
na02f80 g740865 ( .a(n_39289), .b(n_39274), .o(n_39346) );
oa22f80 g774715 ( .a(n_6346), .b(n_5403), .c(n_6345), .d(n_5404), .o(n_6405) );
in01f80 g742299 ( .a(n_37900), .o(n_37973) );
in01f80 FE_RC_2983_0 ( .a(n_9198), .o(FE_RN_1302_0) );
in01f80 g749537 ( .a(n_31815), .o(n_31816) );
no02f80 g742482 ( .a(n_37564), .b(n_37537), .o(n_37649) );
na02f80 g737320 ( .a(n_42839), .b(n_42409), .o(n_42859) );
in01f80 g764334 ( .a(n_16742), .o(n_16743) );
na02f80 g740579 ( .a(n_39662), .b(n_39661), .o(n_39693) );
na02f80 g771770 ( .a(n_8995), .b(n_44575), .o(n_9097) );
in01f80 g757413 ( .a(n_22965), .o(n_22966) );
na02f80 g751623 ( .a(n_29249), .b(n_29174), .o(n_29248) );
na02f80 FE_RC_4242_0 ( .a(n_21644), .b(FE_RN_1864_0), .o(n_21964) );
no02f80 g776836 ( .a(n_3918), .b(n_3919), .o(n_4083) );
in01f80 g769370 ( .a(n_12079), .o(n_12047) );
in01f80 g769322 ( .a(n_11894), .o(n_11973) );
no02f80 g770777 ( .a(n_9934), .b(n_9929), .o(n_10030) );
in01f80 newInst_2519 ( .a(newNet_2518), .o(newNet_2519) );
na02f80 g764210 ( .a(n_16772), .b(n_16385), .o(n_16930) );
in01f80 g743156 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_7_), .o(n_36933) );
in01f80 g756418 ( .a(n_24259), .o(n_24216) );
oa12f80 g736636 ( .a(n_299), .b(n_43115), .c(FE_OFN5_n_43918), .o(n_43237) );
oa12f80 g768434 ( .a(n_12434), .b(n_45659), .c(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .o(n_12495) );
no02f80 g775038 ( .a(n_5893), .b(n_4675), .o(n_5923) );
in01f80 g765662 ( .a(n_14986), .o(n_15012) );
in01f80 g756604 ( .a(n_23684), .o(n_23630) );
in01f80 g779525 ( .a(n_1586), .o(n_1587) );
na02f80 g779322 ( .a(n_1638), .b(n_892), .o(n_1730) );
no02f80 g778478 ( .a(n_2397), .b(n_2396), .o(n_2398) );
in01f80 g752916 ( .a(n_27951), .o(n_28105) );
no02f80 g764614 ( .a(n_15988), .b(n_15893), .o(n_16072) );
oa12f80 g750985 ( .a(n_30067), .b(n_30064), .c(n_29944), .o(n_30163) );
in01f80 g763475 ( .a(n_16908), .o(n_16909) );
in01f80 g743707 ( .a(n_36392), .o(n_36393) );
no03m80 g747962 ( .a(n_33146), .b(n_33073), .c(n_32608), .o(n_33193) );
in01f80 g737342 ( .a(n_42867), .o(n_42868) );
in01f80 newInst_1147 ( .a(newNet_1146), .o(newNet_1147) );
oa12f80 g758627 ( .a(n_21700), .b(n_21964), .c(n_21634), .o(n_21985) );
in01f80 newInst_1601 ( .a(newNet_1600), .o(newNet_1601) );
no02f80 FE_RC_2381_0 ( .a(FE_RN_926_0), .b(FE_RN_928_0), .o(FE_RN_929_0) );
in01f80 g753123 ( .a(n_27502), .o(n_27503) );
in01f80 newInst_1433 ( .a(newNet_1432), .o(newNet_1433) );
na02f80 g747224 ( .a(n_33765), .b(n_33817), .o(n_33818) );
no02f80 g736649 ( .a(n_43369), .b(n_43216), .o(n_43478) );
in01f80 FE_RC_1412_0 ( .a(n_15727), .o(FE_RN_411_0) );
na02f80 g769228 ( .a(FE_OCP_RBN3093_n_11475), .b(n_10935), .o(n_11552) );
na02f80 g766564 ( .a(n_13994), .b(n_13923), .o(n_14065) );
na02f80 FE_RC_3099_0 ( .a(n_14805), .b(FE_RN_1369_0), .o(FE_RN_1370_0) );
in01f80 g759904 ( .a(n_21751), .o(n_21693) );
in01f80 g750662 ( .a(n_30394), .o(n_30440) );
na02f80 g774462 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .o(n_6626) );
in01f80 g739091 ( .a(n_41031), .o(n_41065) );
ao22s80 FE_RC_3727_0 ( .a(FE_OCP_RBN3512_n_13960), .b(n_14287), .c(FE_OCP_RBN3514_n_13960), .d(n_14336), .o(n_14519) );
na02f80 g770148 ( .a(FE_OCP_RBN2900_n_44853), .b(n_10699), .o(n_10700) );
no02f80 g750926 ( .a(n_30185), .b(n_30254), .o(n_30255) );
no02f80 g747278 ( .a(n_45753), .b(n_33335), .o(n_33722) );
na02f80 g770905 ( .a(n_8562), .b(n_9904), .o(n_9942) );
in01f80 g737443 ( .a(n_42718), .o(n_42719) );
in01f80 g747006 ( .a(n_33010), .o(n_33011) );
no02f80 g776035 ( .a(FE_OCP_RBN2838_n_4692), .b(n_4182), .o(n_4769) );
no02f80 g752552 ( .a(n_27602), .b(n_27601), .o(n_27603) );
in01f80 g781391 ( .a(beta_8), .o(n_77) );
no02f80 g742770 ( .a(n_37298), .b(n_36952), .o(n_37340) );
in01f80 g760066 ( .a(n_20670), .o(n_20671) );
in01f80 g773511 ( .a(n_8568), .o(n_7509) );
ms00f80 cos_out_reg_22_ ( .ck(newNet_3718), .d(n_43870), .o(cos_out_22) );
in01f80 g762014 ( .a(n_18357), .o(n_18358) );
in01f80 FE_OCPC3186_FE_OCP_RBN1140_n_25816 ( .a(FE_OCPN3185_FE_OCP_RBN1140_n_25816), .o(FE_OCPN3186_FE_OCP_RBN1140_n_25816) );
in01f80 newInst_944 ( .a(newNet_943), .o(newNet_944) );
oa12f80 g775647 ( .a(n_5226), .b(n_5510), .c(n_5325), .o(n_5590) );
oa12f80 g758869 ( .a(n_21519), .b(n_22119), .c(n_21482), .o(n_22177) );
na02f80 g772440 ( .a(n_8489), .b(FE_OCPN1396_n_7881), .o(n_8508) );
in01f80 FE_OCP_RBC1333_n_20249 ( .a(FE_OCP_RBN1332_n_20249), .o(FE_OCP_RBN1333_n_20249) );
in01f80 g742220 ( .a(n_38323), .o(n_38324) );
no02f80 g777911 ( .a(n_3054), .b(n_3160), .o(n_3185) );
na02f80 g751063 ( .a(n_30431), .b(n_30029), .o(n_30900) );
na02f80 g741451 ( .a(n_38770), .b(n_38691), .o(n_38769) );
na02f80 g764459 ( .a(n_16267), .b(n_14577), .o(n_16318) );
in01f80 g754440 ( .a(n_25753), .o(n_25754) );
oa12f80 g742835 ( .a(n_37213), .b(n_37212), .c(n_37211), .o(n_37240) );
no02f80 g768649 ( .a(n_12106), .b(n_11840), .o(n_12146) );
in01f80 FE_OCP_RBC2967_n_26580 ( .a(n_26580), .o(FE_OCP_RBN2967_n_26580) );
in01f80 g752546 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .o(n_27637) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_3_ ( .ck(newNet_3378), .d(n_26536), .o(delay_add_ln22_unr17_stage7_stallmux_q_3_) );
na02f80 g742208 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38293), .o(n_38295) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_26_ ( .ck(newNet_2735), .d(n_17685), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_) );
oa22f80 FE_RC_854_0 ( .a(n_9527), .b(n_9566), .c(n_9565), .d(n_9528), .o(n_9742) );
no02f80 FE_RC_3484_0 ( .a(FE_RN_1498_0), .b(n_37299), .o(n_37380) );
no02f80 g745745 ( .a(n_34478), .b(n_34522), .o(n_34600) );
no02f80 g736973 ( .a(FE_OCPN913_n_43022), .b(n_43300), .o(n_43342) );
in01f80 g740643 ( .a(FE_OCP_RBN2896_n_39575), .o(n_39590) );
no03m80 FE_RC_3779_0 ( .a(n_27309), .b(n_27223), .c(n_27308), .o(n_27353) );
ao12f80 g768893 ( .a(n_12055), .b(n_45685), .c(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .o(n_12393) );
no02f80 g751457 ( .a(n_28492), .b(n_28550), .o(n_28572) );
in01f80 g760112 ( .a(n_20463), .o(n_20464) );
no02f80 FE_RC_35_0 ( .a(FE_RN_8_0), .b(n_6094), .o(n_6158) );
oa12f80 g764606 ( .a(n_15980), .b(n_16142), .c(n_16067), .o(n_16179) );
in01f80 newInst_3512 ( .a(newNet_3235), .o(newNet_3512) );
in01f80 FE_OCP_RBC2977_n_5555 ( .a(FE_OCP_RBN2976_n_5555), .o(FE_OCP_RBN2977_n_5555) );
in01f80 FE_OCP_RBC2520_n_8762 ( .a(FE_OCP_RBN2519_n_8762), .o(FE_OCP_RBN2520_n_8762) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_18_ ( .ck(newNet_242), .d(n_46179), .o(delay_xor_ln22_unr6_stage3_stallmux_q_18_) );
in01f80 FE_RC_2239_0 ( .a(n_37161), .o(FE_RN_818_0) );
no02f80 g778388 ( .a(n_2467), .b(FE_OCPN3761_n_2466), .o(n_2573) );
oa12f80 g752717 ( .a(n_27074), .b(n_27104), .c(n_27056), .o(n_27244) );
oa22f80 FE_RC_4268_0 ( .a(n_21227), .b(FE_OCP_RBN3855_n_21224), .c(n_21224), .d(n_21228), .o(n_21435) );
ao12f80 g782660 ( .a(FE_OFN756_n_44461), .b(n_10411), .c(n_10270), .o(n_44053) );
ao12f80 g779468 ( .a(n_1450), .b(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .o(n_1476) );
na02f80 FE_RC_2015_0 ( .a(FE_RN_665_0), .b(n_14021), .o(FE_RN_666_0) );
in01f80 g772676 ( .a(n_8215), .o(n_8289) );
na02f80 g745724 ( .a(n_35431), .b(n_35417), .o(n_35842) );
in01f80 newInst_3136 ( .a(newNet_3135), .o(newNet_3136) );
in01f80 g759098 ( .a(n_21318), .o(n_21319) );
na02f80 g774911 ( .a(n_6151), .b(n_6122), .o(n_6228) );
no02f80 g746585 ( .a(n_34810), .b(n_34802), .o(n_34885) );
oa12f80 g779113 ( .a(n_1951), .b(n_1950), .c(n_1949), .o(n_2237) );
in01f80 newInst_681 ( .a(newNet_680), .o(newNet_681) );
in01f80 g753848 ( .a(n_26424), .o(n_26458) );
na02f80 g751890 ( .a(n_28841), .b(n_28840), .o(n_28909) );
oa22f80 g780190 ( .a(n_1069), .b(n_817), .c(n_1061), .d(n_779), .o(n_1139) );
no02f80 g751955 ( .a(n_28793), .b(n_28860), .o(n_28902) );
na02f80 g749257 ( .a(n_30824), .b(FE_OCPN1490_n_30823), .o(n_30825) );
na02f80 g771517 ( .a(n_9153), .b(n_9101), .o(n_9370) );
no02f80 g764398 ( .a(n_16126), .b(n_16163), .o(n_16330) );
na02f80 g768276 ( .a(n_12621), .b(n_12618), .o(n_12622) );
in01f80 g737891 ( .a(n_42606), .o(n_42607) );
na02f80 g741916 ( .a(n_38145), .b(n_38035), .o(n_38171) );
in01f80 FE_OCP_RBC3684_FE_RN_770_0 ( .a(FE_RN_770_0), .o(FE_OCP_RBN3684_FE_RN_770_0) );
ms00f80 cos_out_reg_31_ ( .ck(newNet_3689), .d(n_43905), .o(cos_out_31) );
na02f80 g769112 ( .a(n_11674), .b(n_11629), .o(n_11856) );
no02f80 FE_RC_501_0 ( .a(FE_RN_150_0), .b(FE_RN_151_0), .o(FE_RN_152_0) );
in01f80 newInst_933 ( .a(newNet_932), .o(newNet_933) );
in01f80 g757633 ( .a(n_22774), .o(n_22751) );
in01f80 newInst_1775 ( .a(newNet_1774), .o(newNet_1775) );
in01f80 g758675 ( .a(n_21815), .o(n_21845) );
no02f80 g748350 ( .a(n_31786), .b(n_31758), .o(n_31858) );
in01f80 FE_RC_1762_0 ( .a(n_12170), .o(FE_RN_504_0) );
no02f80 g755270 ( .a(n_24941), .b(n_24974), .o(n_24942) );
in01f80 g744261 ( .a(n_35590), .o(n_35570) );
na02f80 g770141 ( .a(n_10821), .b(n_10713), .o(n_10822) );
na02f80 g753082 ( .a(n_27233), .b(n_27232), .o(n_27270) );
ao12f80 g741784 ( .a(n_38241), .b(n_38420), .c(n_38165), .o(n_38474) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_26_ ( .ck(newNet_2546), .d(n_27739), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_) );
no02f80 FE_RC_3976_0 ( .a(FE_RN_1721_0), .b(n_29518), .o(FE_RN_1722_0) );
no02f80 g740230 ( .a(n_39764), .b(n_39763), .o(n_39773) );
in01f80 newInst_2793 ( .a(newNet_2792), .o(newNet_2793) );
no02f80 g759710 ( .a(n_20417), .b(FE_OFN751_n_45003), .o(n_20508) );
in01f80 FE_OCP_RBC3428_n_12890 ( .a(n_12890), .o(FE_OCP_RBN3428_n_12890) );
no02f80 g759230 ( .a(n_21344), .b(FE_OCP_DRV_N1590_n_21343), .o(n_21456) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_2_ ( .ck(newNet_2261), .d(n_39847), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_23_ ( .ck(newNet_1840), .d(n_16924), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_) );
ao22s80 g737269 ( .a(n_42844), .b(n_42618), .c(n_42845), .d(n_42619), .o(n_42906) );
no02f80 g745367 ( .a(FE_OCP_RBN2995_n_35539), .b(n_35298), .o(n_36082) );
in01f80 FE_RC_4258_0 ( .a(n_22580), .o(FE_RN_1875_0) );
oa12f80 g738270 ( .a(n_41712), .b(n_41801), .c(n_41640), .o(n_41899) );
in01f80 FE_OCPC1478_n_28775 ( .a(FE_OCPN1477_n_28775), .o(FE_OCPN1478_n_28775) );
in01f80 g752365 ( .a(n_27784), .o(n_27757) );
na02f80 g765146 ( .a(n_15151), .b(n_15235), .o(n_15277) );
na03f80 g762171 ( .a(n_18701), .b(n_18703), .c(n_18449), .o(n_18702) );
na02f80 g761456 ( .a(n_19647), .b(n_19677), .o(n_19710) );
na02f80 g739588 ( .a(FE_OCP_RBN3338_n_44610), .b(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .o(n_40608) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_25_ ( .ck(newNet_707), .d(n_46192), .o(delay_xor_ln21_unr6_stage3_stallmux_q_25_) );
no02f80 g771861 ( .a(n_9774), .b(n_9828), .o(n_10751) );
no02f80 g738581 ( .a(n_41827), .b(n_41879), .o(n_41918) );
na02f80 g773916 ( .a(n_6935), .b(delay_add_ln22_unr5_stage3_stallmux_q_7_), .o(n_7037) );
in01f80 g742707 ( .a(n_37371), .o(n_37372) );
no02f80 g774326 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .o(n_6644) );
no02f80 g763825 ( .a(n_17354), .b(n_17104), .o(n_17961) );
in01f80 FE_OCP_RBC3411_n_33547 ( .a(n_33547), .o(FE_OCP_RBN3411_n_33547) );
na02f80 g746748 ( .a(n_33378), .b(n_33376), .o(n_33406) );
in01f80 g744944 ( .a(n_35684), .o(n_35025) );
no02f80 g775013 ( .a(n_6147), .b(n_6044), .o(n_6162) );
no02f80 g745010 ( .a(n_34830), .b(n_34794), .o(n_34903) );
in01f80 g741306 ( .a(n_38904), .o(n_38937) );
na02f80 g778321 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_29_), .o(n_2975) );
in01f80 g742687 ( .a(n_37420), .o(n_37412) );
in01f80 FE_OCP_RBC3049_n_11329 ( .a(n_11329), .o(FE_OCP_RBN3049_n_11329) );
in01f80 FE_RC_2166_0 ( .a(n_45024), .o(FE_RN_769_0) );
ao22s80 g770979 ( .a(n_9714), .b(n_9701), .c(n_9713), .d(n_9660), .o(n_9892) );
in01f80 g768716 ( .a(n_12158), .o(n_12133) );
ao12f80 g748670 ( .a(n_31297), .b(n_31399), .c(n_31352), .o(n_31421) );
in01f80 g747141 ( .a(n_34643), .o(n_33993) );
no02f80 g773130 ( .a(n_7712), .b(n_7707), .o(n_7783) );
in01f80 g748173 ( .a(n_32132), .o(n_32133) );
in01f80 newInst_3177 ( .a(newNet_3176), .o(newNet_3177) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_8_ ( .ck(newNet_1787), .d(n_16523), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_) );
no02f80 g739374 ( .a(n_40813), .b(n_40812), .o(n_41237) );
in01f80 newInst_3349 ( .a(newNet_3348), .o(newNet_3349) );
in01f80 g757203 ( .a(n_23245), .o(n_23281) );
in01f80 FE_OCP_RBC2818_n_4458 ( .a(n_4458), .o(FE_OCP_RBN2818_n_4458) );
na02f80 g776632 ( .a(n_4285), .b(n_4071), .o(n_4389) );
na02f80 g746757 ( .a(n_34169), .b(n_34168), .o(n_34170) );
no02f80 FE_RC_2950_0 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(n_35063), .o(FE_RN_1288_0) );
in01f80 FE_OCP_RBC3381_n_1732 ( .a(n_1732), .o(FE_OCP_RBN3381_n_1732) );
oa22f80 g754881 ( .a(n_25542), .b(n_24857), .c(FE_OCPN1026_n_25481), .d(n_24872), .o(n_25775) );
no02f80 g750440 ( .a(n_29607), .b(n_29606), .o(n_29608) );
na02f80 g741157 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39181), .o(n_39251) );
na03f80 FE_RC_3930_0 ( .a(n_32632), .b(n_32687), .c(n_32636), .o(n_32754) );
in01f80 g765390 ( .a(n_15023), .o(n_15055) );
in01f80 g761599 ( .a(n_19980), .o(n_20086) );
na02f80 g741933 ( .a(n_38141), .b(n_44029), .o(n_38187) );
no02f80 g758189 ( .a(n_22434), .b(n_22213), .o(n_22500) );
na02f80 g744224 ( .a(n_36182), .b(n_36134), .o(n_36287) );
no02f80 g740097 ( .a(n_40220), .b(n_39921), .o(n_40326) );
oa22f80 g784346 ( .a(FE_OFN86_n_46137), .b(n_6005), .c(FE_OCP_RBN3076_FE_OFN807_n_46195), .d(n_6047), .o(n_46152) );
no02f80 g767089 ( .a(n_13734), .b(n_13733), .o(n_13735) );
oa22f80 FE_RC_1632_0 ( .a(n_16950), .b(n_17237), .c(n_16995), .d(n_17238), .o(n_17459) );
na02f80 FE_RC_3082_0 ( .a(FE_OCP_RBN1700_n_19353), .b(n_19461), .o(FE_RN_1359_0) );
in01f80 g773167 ( .a(n_7921), .o(n_7988) );
ao12f80 g754748 ( .a(n_25334), .b(n_25366), .c(n_25333), .o(n_27018) );
na02f80 g757986 ( .a(n_22153), .b(n_22129), .o(n_22270) );
in01f80 g737627 ( .a(n_42661), .o(n_42662) );
na02f80 g776942 ( .a(n_3583), .b(n_3509), .o(n_3607) );
na02f80 g763215 ( .a(n_16954), .b(n_17008), .o(n_17199) );
na02f80 FE_RC_653_0 ( .a(FE_RN_209_0), .b(n_6933), .o(n_7002) );
no02f80 g759284 ( .a(n_20920), .b(n_20855), .o(n_20975) );
oa12f80 g784669 ( .a(n_5592), .b(n_5506), .c(n_5559), .o(n_46999) );
in01f80 newInst_1031 ( .a(newNet_1030), .o(newNet_1031) );
in01f80 newInst_355 ( .a(newNet_354), .o(newNet_355) );
in01f80 g754020 ( .a(n_26206), .o(n_26207) );
no02f80 g766866 ( .a(FE_OCP_RBN2324_n_13616), .b(FE_OCP_RBN2246_n_13017), .o(n_13644) );
oa12f80 g758973 ( .a(n_21996), .b(n_22011), .c(n_21995), .o(n_22031) );
oa12f80 g777887 ( .a(n_2271), .b(n_3147), .c(n_2313), .o(n_3204) );
na02f80 g746164 ( .a(n_33648), .b(n_33196), .o(n_33665) );
in01f80 g737532 ( .a(n_42550), .o(n_42551) );
in01f80 g763106 ( .a(n_17548), .o(n_17549) );
no02f80 g748273 ( .a(FE_OCP_RBN3735_n_31819), .b(n_30711), .o(n_32049) );
in01f80 newInst_62 ( .a(newNet_61), .o(newNet_62) );
na02f80 g770593 ( .a(FE_OCP_RBN3666_n_10106), .b(n_9146), .o(n_10329) );
no02f80 g771968 ( .a(FE_OCP_RBN3644_n_44490), .b(n_8688), .o(n_9774) );
in01f80 g777370 ( .a(n_3997), .o(n_3998) );
in01f80 g741672 ( .a(FE_OCP_RBN2397_n_38586), .o(n_38608) );
oa12f80 g749401 ( .a(n_31343), .b(n_31981), .c(n_31279), .o(n_32006) );
in01f80 newInst_3101 ( .a(newNet_3100), .o(newNet_3101) );
na02f80 g764731 ( .a(n_15796), .b(FE_OCP_RBN2941_FE_RN_473_0), .o(n_15897) );
no02f80 g744095 ( .a(n_44223), .b(n_35060), .o(n_36531) );
no02f80 g744317 ( .a(n_35505), .b(n_35504), .o(n_35553) );
na02f80 g752821 ( .a(n_27310), .b(n_27230), .o(n_27356) );
in01f80 g775403 ( .a(n_5586), .o(n_5649) );
no02f80 g768059 ( .a(n_12914), .b(n_12257), .o(n_13035) );
no02f80 g738170 ( .a(n_42027), .b(n_42014), .o(n_42015) );
no02f80 g778346 ( .a(n_2599), .b(FE_OCP_RBN2274_n_2457), .o(n_2600) );
na02f80 g779245 ( .a(n_1766), .b(n_1038), .o(n_1844) );
na02f80 g771185 ( .a(n_9161), .b(n_9144), .o(n_9360) );
in01f80 newInst_2663 ( .a(newNet_2662), .o(newNet_2663) );
in01f80 g763450 ( .a(n_17317), .o(n_17318) );
na02f80 g740827 ( .a(n_39374), .b(n_39321), .o(n_39405) );
in01f80 newInst_331 ( .a(newNet_330), .o(newNet_331) );
na02f80 g779097 ( .a(n_1987), .b(n_1981), .o(n_1982) );
na02f80 g776637 ( .a(n_4081), .b(n_4046), .o(n_4286) );
no02f80 g758223 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .o(n_22845) );
oa12f80 g770097 ( .a(n_10943), .b(n_10951), .c(n_10942), .o(n_10981) );
in01f80 g778713 ( .a(n_2452), .o(n_2404) );
in01f80 g768724 ( .a(n_12162), .o(n_12132) );
in01f80 newInst_1070 ( .a(newNet_363), .o(newNet_1070) );
in01f80 g739720 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .o(n_40522) );
na02f80 FE_RC_2372_0 ( .a(n_42358), .b(n_42562), .o(FE_RN_921_0) );
no02f80 g744578 ( .a(n_35383), .b(n_35382), .o(n_35393) );
in01f80 FE_RC_3975_0 ( .a(FE_RN_1722_0), .o(n_29585) );
in01f80 newInst_3548 ( .a(newNet_3547), .o(newNet_3548) );
no02f80 g759303 ( .a(n_20805), .b(n_45024), .o(n_20865) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_10_ ( .ck(newNet_423), .d(n_32567), .o(delay_xor_ln22_unr21_stage8_stallmux_q_10_) );
ao12f80 g774199 ( .a(n_6873), .b(n_6872), .c(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .o(n_6988) );
na02f80 g754325 ( .a(n_25813), .b(n_25479), .o(n_25855) );
oa12f80 g747209 ( .a(n_32597), .b(n_32643), .c(FE_OCP_RBN3370_n_32436), .o(n_32698) );
no02f80 g772025 ( .a(n_8711), .b(FE_OCP_RBN2492_n_8508), .o(n_8751) );
in01f80 g769881 ( .a(n_11259), .o(n_11260) );
no02f80 g755290 ( .a(n_25638), .b(n_25637), .o(n_25639) );
no02f80 g736741 ( .a(n_43152), .b(n_43085), .o(n_43091) );
na02f80 g764318 ( .a(n_16373), .b(n_16283), .o(n_16397) );
ao22s80 FE_RC_976_0 ( .a(n_27503), .b(n_44265), .c(n_27620), .d(n_27502), .o(n_27736) );
in01f80 newInst_2367 ( .a(newNet_809), .o(newNet_2367) );
no02f80 g779784 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n_1422) );
na02f80 g768500 ( .a(n_12299), .b(n_12335), .o(n_12551) );
in01f80 g751574 ( .a(n_28491), .o(n_28501) );
oa12f80 g745983 ( .a(n_35244), .b(n_35243), .c(n_35242), .o(n_35763) );
na02f80 g763898 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .o(n_17302) );
na02f80 g767407 ( .a(n_13545), .b(n_13544), .o(n_13546) );
no02f80 g781106 ( .a(n_244), .b(n_156), .o(n_239) );
in01f80 g751450 ( .a(n_28802), .o(n_28803) );
na02f80 g768455 ( .a(n_12378), .b(n_12377), .o(n_12379) );
oa12f80 g759336 ( .a(n_21889), .b(n_21888), .c(n_21887), .o(n_21932) );
na02f80 FE_RC_2769_0 ( .a(n_2626), .b(FE_RN_1179_0), .o(n_2778) );
in01f80 FE_RC_3825_0 ( .a(FE_RN_1668_0), .o(n_23467) );
no02f80 g743985 ( .a(n_35574), .b(n_35516), .o(n_35599) );
no02f80 g779172 ( .a(n_1874), .b(n_1873), .o(n_1875) );
in01f80 g754559 ( .a(n_26899), .o(n_26900) );
oa22f80 FE_RC_1048_0 ( .a(n_39226), .b(n_39467), .c(n_39227), .d(n_39466), .o(n_39551) );
in01f80 newInst_3672 ( .a(newNet_3671), .o(newNet_3672) );
in01f80 g753607 ( .a(n_26721), .o(n_26722) );
na02f80 g742715 ( .a(n_37408), .b(n_37210), .o(n_37497) );
in01f80 newInst_1185 ( .a(newNet_1184), .o(newNet_1185) );
ao12f80 g780057 ( .a(n_818), .b(n_1225), .c(n_842), .o(n_1232) );
no02f80 g771297 ( .a(n_9214), .b(n_9366), .o(n_9413) );
ao12f80 g742756 ( .a(n_37231), .b(n_37291), .c(n_37186), .o(n_37299) );
ao22s80 FE_RC_608_0 ( .a(n_38153), .b(n_38418), .c(n_38154), .d(n_38419), .o(n_38515) );
no02f80 g759558 ( .a(n_21724), .b(n_21781), .o(n_21782) );
na02f80 g740103 ( .a(n_40182), .b(n_40013), .o(n_40285) );
ao22s80 g780306 ( .a(n_922), .b(n_1148), .c(n_903), .d(n_770), .o(n_954) );
in01f80 newInst_2050 ( .a(newNet_2049), .o(newNet_2050) );
in01f80 FE_OFC760_n_45813 ( .a(FE_OFN757_n_45813), .o(FE_OFN760_n_45813) );
na02f80 g762387 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18065), .o(n_18659) );
in01f80 g743494 ( .a(n_37625), .o(n_36686) );
na02f80 g778651 ( .a(n_2455), .b(n_2012), .o(n_2514) );
na02f80 g736797 ( .a(n_43111), .b(n_43062), .o(n_43145) );
no02f80 g740261 ( .a(n_40060), .b(n_40059), .o(n_40102) );
in01f80 g739726 ( .a(n_40543), .o(n_40550) );
in01f80 fopt783151 ( .a(n_1282), .o(n_44652) );
in01f80 g779307 ( .a(n_2442), .o(n_2461) );
no02f80 g739007 ( .a(n_41156), .b(n_41126), .o(n_41157) );
ao22s80 FE_RC_1294_0 ( .a(n_38778), .b(n_38606), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .d(n_38605), .o(n_38669) );
na02f80 g752032 ( .a(n_28071), .b(n_28002), .o(n_28072) );
in01f80 newInst_1323 ( .a(newNet_1202), .o(newNet_1323) );
in01f80 g751161 ( .a(n_30096), .o(n_30029) );
no02f80 g774084 ( .a(n_6835), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n_6803) );
no02f80 g777264 ( .a(n_3576), .b(FE_OCP_RBN2537_n_3645), .o(n_3599) );
in01f80 g769773 ( .a(n_11198), .o(n_11199) );
in01f80 FE_OCP_RBC2619_n_44561 ( .a(FE_OCP_RBN2617_n_44561), .o(FE_OCP_RBN2619_n_44561) );
ao12f80 g752482 ( .a(FE_OCPN1750_n_27223), .b(n_27661), .c(n_27144), .o(n_27723) );
na02f80 FE_RC_4081_0 ( .a(FE_RN_1779_0), .b(FE_RN_1780_0), .o(FE_RN_1781_0) );
in01f80 newInst_2422 ( .a(newNet_2421), .o(newNet_2422) );
na02f80 g746122 ( .a(n_33695), .b(n_33179), .o(n_33718) );
na02f80 g756918 ( .a(n_23833), .b(n_23864), .o(n_23936) );
na02f80 g752815 ( .a(n_27764), .b(n_27812), .o(n_27851) );
oa12f80 g765367 ( .a(n_15784), .b(n_15874), .c(n_15711), .o(n_16304) );
in01f80 g766339 ( .a(n_14365), .o(n_14398) );
na02f80 g780241 ( .a(n_1003), .b(n_1002), .o(n_1041) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_1_ ( .ck(newNet_3421), .d(n_26439), .o(delay_add_ln22_unr17_stage7_stallmux_q_1_) );
no02f80 g761789 ( .a(n_19197), .b(n_19196), .o(n_19198) );
na02f80 g781065 ( .a(sin_out_27), .b(FE_OFN4_n_43918), .o(n_293) );
in01f80 g763446 ( .a(n_17321), .o(n_17322) );
no02f80 FE_RC_220_0 ( .a(FE_RN_72_0), .b(FE_OCP_RBN1103_n_45224), .o(FE_RN_74_0) );
in01f80 g742657 ( .a(n_37505), .o(n_37499) );
na02f80 g757782 ( .a(n_23028), .b(n_23087), .o(n_23088) );
no02f80 g748310 ( .a(n_31554), .b(n_31735), .o(n_31768) );
ao12f80 g757070 ( .a(n_23302), .b(n_23301), .c(n_23300), .o(n_23359) );
oa22f80 FE_RC_981_0 ( .a(n_27484), .b(n_27688), .c(n_44360), .d(n_27485), .o(n_27781) );
no02f80 g756455 ( .a(n_23970), .b(n_23969), .o(n_23997) );
oa22f80 g745789 ( .a(n_44102), .b(n_33895), .c(n_44104), .d(FE_OCP_RBN2283_n_33846), .o(n_34334) );
in01f80 FE_RC_2737_0 ( .a(n_8232), .o(FE_RN_1160_0) );
no02f80 g761485 ( .a(n_19649), .b(n_19650), .o(n_19676) );
oa12f80 g780341 ( .a(n_718), .b(n_739), .c(n_717), .o(n_740) );
in01f80 FE_OCP_RBC2929_n_5221 ( .a(n_5221), .o(FE_OCP_RBN2929_n_5221) );
in01f80 g759058 ( .a(n_21495), .o(n_21531) );
ao12f80 g739113 ( .a(n_40782), .b(n_41030), .c(n_40803), .o(n_41083) );
oa12f80 g738018 ( .a(n_42164), .b(n_42163), .c(n_42162), .o(n_42172) );
no02f80 g767584 ( .a(n_13423), .b(n_13470), .o(n_13471) );
oa22f80 FE_RC_1157_0 ( .a(n_32664), .b(FE_OCP_RBN2131_n_32649), .c(n_32663), .d(n_32649), .o(n_32773) );
in01f80 g773941 ( .a(n_7255), .o(n_7256) );
no02f80 g778669 ( .a(n_2289), .b(n_2858), .o(n_2341) );
in01f80 g756333 ( .a(n_24054), .o(n_24055) );
no02f80 g753868 ( .a(n_26306), .b(n_26252), .o(n_26334) );
no02f80 g763020 ( .a(n_17905), .b(n_17266), .o(n_17962) );
in01f80 newInst_578 ( .a(newNet_577), .o(newNet_578) );
na02f80 g756286 ( .a(n_24608), .b(n_23992), .o(n_24737) );
no02f80 g753396 ( .a(n_26989), .b(n_26918), .o(n_27011) );
no02f80 g763121 ( .a(n_17146), .b(n_17045), .o(n_17147) );
ao12f80 g752293 ( .a(n_27918), .b(n_44723), .c(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .o(n_27839) );
in01f80 newInst_2575 ( .a(newNet_2574), .o(newNet_2575) );
in01f80 FE_OCP_RBC3677_n_21051 ( .a(n_21051), .o(FE_OCP_RBN3677_n_21051) );
na02f80 g768687 ( .a(n_12137), .b(delay_add_ln22_unr8_stage4_stallmux_q_5_), .o(n_12251) );
na02f80 g749034 ( .a(n_30918), .b(FE_OCP_DRV_N1584_n_30917), .o(n_31011) );
in01f80 newInst_2842 ( .a(newNet_2841), .o(newNet_2842) );
no02f80 g764669 ( .a(n_15854), .b(n_15455), .o(n_15989) );
na02f80 g753933 ( .a(n_26228), .b(n_25694), .o(n_26263) );
no02f80 g750138 ( .a(n_29813), .b(n_29812), .o(n_29832) );
no02f80 g777990 ( .a(n_3022), .b(n_2635), .o(n_3072) );
in01f80 g763486 ( .a(n_17118), .o(n_17172) );
in01f80 FE_OCPC868_n_16086 ( .a(n_16086), .o(FE_OCPN868_n_16086) );
no02f80 g742212 ( .a(n_44887), .b(n_37849), .o(n_38249) );
na02f80 g753275 ( .a(n_27167), .b(FE_OCP_RBN2909_n_26173), .o(n_27211) );
no02f80 g742211 ( .a(n_37850), .b(n_37849), .o(n_37851) );
in01f80 g739037 ( .a(n_41158), .o(n_41192) );
ao12f80 g784073 ( .a(n_45812), .b(n_970), .c(n_1002), .o(n_45819) );
oa12f80 g741805 ( .a(n_38188), .b(n_38288), .c(n_38169), .o(n_38344) );
in01f80 FE_OCP_RBC3142_n_32395 ( .a(n_32395), .o(FE_OCP_RBN3142_n_32395) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_5_ ( .ck(newNet_1176), .d(n_4526), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_) );
oa12f80 g764942 ( .a(n_15675), .b(n_15674), .c(n_15673), .o(n_15751) );
no02f80 g752946 ( .a(n_27050), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27787) );
in01f80 FE_OCPC1046_n_13570 ( .a(FE_OCPN1045_n_13570), .o(FE_OCPN1046_n_13570) );
ao12f80 g748693 ( .a(n_32561), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n_33192) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_11_ ( .ck(newNet_3261), .d(n_36421), .o(delay_add_ln22_unr23_stage9_stallmux_q_11_) );
na02f80 g780575 ( .a(n_745), .b(n_906), .o(n_976) );
no02f80 g760401 ( .a(n_20096), .b(n_18712), .o(n_20191) );
oa12f80 g736263 ( .a(n_302), .b(n_43901), .c(FE_OFN4_n_43918), .o(n_43915) );
na02f80 g770991 ( .a(n_9743), .b(n_9804), .o(n_9849) );
oa22f80 FE_RC_3433_0 ( .a(n_22381), .b(n_22518), .c(n_22538), .d(n_22382), .o(n_22640) );
in01f80 g763643 ( .a(FE_OCP_RBN1209_n_16814), .o(n_16977) );
na02f80 g781042 ( .a(cos_out_12), .b(FE_OFN2_n_43918), .o(n_348) );
na02f80 g774796 ( .a(n_6261), .b(n_6205), .o(n_6298) );
in01f80 g770377 ( .a(n_10541), .o(n_10511) );
no02f80 g778327 ( .a(n_47024), .b(n_1095), .o(n_2988) );
ao12f80 g747085 ( .a(n_32798), .b(n_32799), .c(n_32797), .o(n_34058) );
oa12f80 g770787 ( .a(n_9422), .b(n_9855), .c(n_9420), .o(n_9860) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_10_ ( .ck(newNet_852), .d(n_1322), .o(delay_xor_ln21_unr3_stage2_stallmux_q_10_) );
in01f80 FE_OCP_RBC2909_n_26173 ( .a(n_26173), .o(FE_OCP_RBN2909_n_26173) );
in01f80 g737100 ( .a(n_43120), .o(n_43242) );
no02f80 g756413 ( .a(n_23742), .b(n_23719), .o(n_23720) );
na02f80 g749723 ( .a(n_31174), .b(n_186), .o(n_31175) );
in01f80 FE_OCPC1466_n_13014 ( .a(FE_OCPN1465_n_13014), .o(FE_OCPN1466_n_13014) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_27_ ( .ck(newNet_1592), .d(n_27588), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_) );
na02f80 g749019 ( .a(n_30834), .b(n_30743), .o(n_30919) );
oa22f80 g743605 ( .a(n_36437), .b(n_36364), .c(n_36438), .d(n_36363), .o(n_36487) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_3_ ( .ck(newNet_217), .d(n_46145), .o(delay_xor_ln22_unr6_stage3_stallmux_q_3_) );
in01f80 g741201 ( .a(n_39098), .o(n_39099) );
na02f80 g771091 ( .a(n_9841), .b(n_9707), .o(n_9922) );
no02f80 g744060 ( .a(n_44222), .b(n_34861), .o(n_35910) );
no02f80 g741897 ( .a(n_38356), .b(n_38355), .o(n_38357) );
in01f80 newInst_3682 ( .a(newNet_3681), .o(newNet_3682) );
no02f80 g777395 ( .a(n_3519), .b(n_3573), .o(n_3629) );
in01f80 g741048 ( .a(n_39457), .o(n_39458) );
ao12f80 g738152 ( .a(n_42015), .b(n_42027), .c(n_42014), .o(n_42115) );
no02f80 g737909 ( .a(n_42202), .b(n_41922), .o(n_42306) );
na02f80 g744046 ( .a(FE_OCPN3751_n_44222), .b(n_34660), .o(n_36265) );
na02f80 g736896 ( .a(n_43485), .b(n_43206), .o(n_43585) );
na02f80 g764678 ( .a(FE_OCP_RBN2800_n_15706), .b(n_14419), .o(n_15775) );
in01f80 newInst_1360 ( .a(newNet_1359), .o(newNet_1360) );
na02f80 g749873 ( .a(FE_OCP_RBN3010_n_31117), .b(n_31275), .o(n_31282) );
no03m80 FE_RC_3705_0 ( .a(n_5797), .b(n_5601), .c(n_5672), .o(n_5905) );
in01f80 FE_OCP_RBC3450_n_37945 ( .a(FE_OCP_RBN3446_n_37945), .o(FE_OCP_RBN3450_n_37945) );
in01f80 FE_RC_3210_0 ( .a(FE_RN_1427_0), .o(FE_RN_1426_0) );
in01f80 newInst_2820 ( .a(newNet_2202), .o(newNet_2820) );
in01f80 newInst_2683 ( .a(newNet_2682), .o(newNet_2683) );
in01f80 FE_OCPC1426_n_18099 ( .a(FE_OCPN1425_n_18099), .o(FE_OCPN1426_n_18099) );
no02f80 g762886 ( .a(n_17771), .b(n_17746), .o(n_17747) );
in01f80 g776964 ( .a(n_3955), .o(n_3877) );
na02f80 g769762 ( .a(FE_OCP_RBN2996_n_11004), .b(n_44498), .o(n_11054) );
in01f80 FE_OCP_RBC3552_n_44575 ( .a(FE_OCP_RBN3545_n_44575), .o(FE_OCP_RBN3552_n_44575) );
na02f80 g751619 ( .a(n_28447), .b(n_27642), .o(n_28484) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_8_ ( .ck(newNet_942), .d(n_22826), .o(delay_xor_ln21_unr15_stage6_stallmux_q_8_) );
in01f80 g749419 ( .a(n_30582), .o(n_30601) );
in01f80 FE_OCPC3177_n_21901 ( .a(n_21901), .o(FE_OCPN3177_n_21901) );
in01f80 g749599 ( .a(n_31773), .o(n_30522) );
in01f80 newInst_384 ( .a(newNet_383), .o(newNet_384) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_8_ ( .ck(newNet_2506), .d(n_26968), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_) );
in01f80 g773066 ( .a(n_7951), .o(n_7952) );
in01f80 g746510 ( .a(n_34913), .o(n_34914) );
in01f80 FE_OCP_RBC2284_n_33846 ( .a(n_33846), .o(FE_OCP_RBN2284_n_33846) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_1_ ( .ck(newNet_3227), .d(n_35409), .o(delay_add_ln22_unr23_stage9_stallmux_q_1_) );
ao12f80 g751431 ( .a(n_28447), .b(n_28543), .c(n_28606), .o(n_28607) );
in01f80 g769365 ( .a(n_11968), .o(n_12076) );
na02f80 g779027 ( .a(n_45717), .b(n_1597), .o(n_2077) );
in01f80 FE_OCP_RBC1725_FE_RN_422_0 ( .a(FE_RN_422_0), .o(FE_OCP_RBN1725_FE_RN_422_0) );
no02f80 g772656 ( .a(n_8164), .b(n_7817), .o(n_8205) );
ao22s80 FE_RC_426_0 ( .a(n_15377), .b(n_15660), .c(n_15376), .d(n_15629), .o(n_15817) );
no02f80 g747615 ( .a(n_34071), .b(n_34070), .o(n_34072) );
na02f80 g739443 ( .a(n_44769), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .o(n_40805) );
na02f80 g770619 ( .a(n_10410), .b(n_10409), .o(n_10454) );
ao12f80 g746563 ( .a(n_34801), .b(n_34810), .c(n_34155), .o(n_35372) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_10_ ( .ck(newNet_931), .d(n_27819), .o(delay_xor_ln21_unr18_stage7_stallmux_q_10_) );
na02f80 g748766 ( .a(n_31354), .b(n_31353), .o(n_31355) );
in01f80 newInst_1983 ( .a(newNet_1572), .o(newNet_1983) );
no02f80 g753592 ( .a(n_26697), .b(n_26519), .o(n_26724) );
oa12f80 g738254 ( .a(n_41895), .b(n_41894), .c(n_41893), .o(n_42358) );
in01f80 g774227 ( .a(n_6852), .o(n_6853) );
in01f80 g754533 ( .a(n_26907), .o(n_26350) );
no02f80 g745330 ( .a(n_35850), .b(n_36082), .o(n_36215) );
na02f80 g761973 ( .a(n_19406), .b(n_18840), .o(n_19049) );
ao12f80 g777758 ( .a(n_3411), .b(n_3410), .c(n_3409), .o(n_3500) );
in01f80 g769691 ( .a(n_11317), .o(n_11340) );
in01f80 g740253 ( .a(n_40311), .o(n_40312) );
oa22f80 g784337 ( .a(FE_OFN775_n_46137), .b(n_5286), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5379), .o(n_46141) );
no02f80 g771665 ( .a(n_9129), .b(n_9169), .o(n_9241) );
in01f80 newInst_1535 ( .a(newNet_1534), .o(newNet_1535) );
oa12f80 g767467 ( .a(n_13427), .b(n_13426), .c(n_13425), .o(n_13501) );
ao12f80 g741847 ( .a(n_38263), .b(n_38262), .c(n_38261), .o(n_38829) );
na02f80 g778979 ( .a(n_2224), .b(n_1946), .o(n_2260) );
in01f80 g762222 ( .a(n_18164), .o(n_18165) );
no02f80 FE_RC_3496_0 ( .a(FE_RN_1507_0), .b(n_31518), .o(FE_RN_1508_0) );
no02f80 g752474 ( .a(n_28378), .b(n_28351), .o(n_28352) );
in01f80 g766618 ( .a(n_15631), .o(n_14391) );
no02f80 g754818 ( .a(n_25280), .b(n_25279), .o(n_25281) );
in01f80 g753623 ( .a(n_46934), .o(n_26747) );
no02f80 g744126 ( .a(n_35553), .b(n_35533), .o(n_35534) );
no02f80 g764957 ( .a(n_15430), .b(n_15500), .o(n_15545) );
ao22s80 FE_RC_3356_0 ( .a(n_26785), .b(n_26747), .c(n_46934), .d(n_26758), .o(n_26844) );
in01f80 FE_OCPC3779_n_36126 ( .a(FE_OCPN3778_n_36126), .o(FE_OCPN3779_n_36126) );
oa12f80 g754367 ( .a(n_25454), .b(n_25727), .c(n_25425), .o(n_25845) );
in01f80 FE_OCP_RBC3711_n_46337 ( .a(FE_OCP_RBN3039_n_46337), .o(FE_OCP_RBN3711_n_46337) );
in01f80 fopt782795 ( .a(n_32290), .o(n_44216) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_19_ ( .ck(newNet_1751), .d(n_22398), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_21_ ( .ck(newNet_1229), .d(n_5992), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_) );
in01f80 g760282 ( .a(n_20299), .o(n_20340) );
na02f80 g738051 ( .a(n_42135), .b(n_42121), .o(n_42147) );
oa22f80 FE_RC_211_0 ( .a(n_14244), .b(n_14412), .c(n_14285), .d(n_14413), .o(n_14554) );
in01f80 newInst_344 ( .a(newNet_343), .o(newNet_344) );
no02f80 g753548 ( .a(n_26695), .b(n_26614), .o(n_26759) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_1_ ( .ck(newNet_3536), .d(n_21027), .o(delay_add_ln22_unr14_stage6_stallmux_q_1_) );
oa12f80 g772468 ( .a(n_8263), .b(n_8403), .c(n_8313), .o(n_8460) );
na02f80 g748068 ( .a(n_31971), .b(n_31933), .o(n_32026) );
no02f80 g781320 ( .a(beta_31), .b(beta_5), .o(n_65) );
na02f80 g775268 ( .a(n_5713), .b(n_5669), .o(n_5818) );
oa22f80 FE_RC_139_0 ( .a(n_12830), .b(n_12533), .c(n_12534), .d(FE_OCP_RBN2197_n_12830), .o(n_12981) );
na02f80 g750332 ( .a(n_30687), .b(n_30100), .o(n_30786) );
in01f80 g749735 ( .a(n_31391), .o(n_31392) );
na02f80 g755445 ( .a(n_24820), .b(n_24632), .o(n_24853) );
in01f80 FE_OCP_RBC3479_n_3006 ( .a(n_3006), .o(FE_OCP_RBN3479_n_3006) );
na02f80 g778955 ( .a(n_2197), .b(n_1101), .o(n_2265) );
no02f80 g778736 ( .a(n_45903), .b(n_2702), .o(n_2211) );
in01f80 newInst_2894 ( .a(newNet_2893), .o(newNet_2894) );
no02f80 g751900 ( .a(n_28986), .b(n_28943), .o(n_29431) );
in01f80 g758025 ( .a(n_22080), .o(n_22106) );
no03m80 FE_RC_2508_0 ( .a(FE_RN_1019_0), .b(n_17884), .c(n_17885), .o(n_17914) );
oa22f80 g754477 ( .a(n_26907), .b(n_26856), .c(n_26350), .d(n_26896), .o(n_26935) );
oa12f80 g748851 ( .a(n_31055), .b(n_31054), .c(n_31053), .o(n_31110) );
ao12f80 g751021 ( .a(n_29944), .b(n_30000), .c(n_29999), .o(n_30034) );
in01f80 g743115 ( .a(n_37205), .o(n_37044) );
no02f80 FE_RC_4063_0 ( .a(n_35740), .b(n_35739), .o(FE_RN_1768_0) );
no02f80 g775128 ( .a(n_5813), .b(n_4556), .o(n_5831) );
no02f80 FE_RC_794_0 ( .a(FE_RN_240_0), .b(FE_RN_241_0), .o(FE_RN_242_0) );
ao12f80 g742934 ( .a(n_37002), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n_37063) );
na02f80 g764620 ( .a(n_15898), .b(FE_OCPN3775_n_14730), .o(n_15997) );
in01f80 g751942 ( .a(n_28147), .o(n_28148) );
na02f80 g770039 ( .a(FE_OCP_RBN3692_n_10852), .b(FE_OCP_RBN3643_n_44490), .o(n_10888) );
oa12f80 g743855 ( .a(n_37025), .b(n_46250), .c(n_46229), .o(n_37166) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_12_ ( .ck(newNet_923), .d(n_27862), .o(delay_xor_ln21_unr18_stage7_stallmux_q_12_) );
in01f80 g755421 ( .a(n_25440), .o(n_25441) );
ao22s80 FE_RC_3327_0 ( .a(FE_OCP_RBN3206_n_44365), .b(FE_OCP_RBN1677_n_44847), .c(n_44847), .d(FE_OCP_RBN3209_n_44365), .o(n_16829) );
in01f80 newInst_3160 ( .a(newNet_3159), .o(newNet_3160) );
oa12f80 g762068 ( .a(n_18178), .b(n_18177), .c(n_18176), .o(n_18224) );
in01f80 g743010 ( .a(n_36960), .o(n_36961) );
oa12f80 g752576 ( .a(n_28279), .b(n_28298), .c(n_28278), .o(n_28810) );
in01f80 g743733 ( .a(n_36248), .o(n_36279) );
in01f80 FE_OCP_RBC2563_n_34905 ( .a(n_34905), .o(FE_OCP_RBN2563_n_34905) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_29_ ( .ck(newNet_1818), .d(n_17103), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_) );
in01f80 g779446 ( .a(n_1649), .o(n_1650) );
in01f80 g747101 ( .a(n_32954), .o(n_32955) );
in01f80 FE_OCPC907_n_23227 ( .a(n_23227), .o(FE_OCPN907_n_23227) );
no02f80 g776434 ( .a(n_4265), .b(n_4182), .o(n_4549) );
oa12f80 g784621 ( .a(n_39472), .b(n_39431), .c(n_39391), .o(n_46950) );
in01f80 g770942 ( .a(n_9899), .o(n_9900) );
oa22f80 g758379 ( .a(n_22528), .b(n_21864), .c(n_22527), .d(n_21863), .o(n_22588) );
in01f80 g779165 ( .a(n_2218), .o(n_2622) );
na02f80 g761002 ( .a(n_19274), .b(n_18915), .o(n_19275) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_10_ ( .ck(newNet_1881), .d(n_16550), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_) );
ao12f80 g752832 ( .a(n_28326), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(n_28756) );
no02f80 g771448 ( .a(n_9317), .b(n_9341), .o(n_9404) );
na02f80 g753673 ( .a(n_26553), .b(n_23509), .o(n_26620) );
in01f80 g751631 ( .a(FE_OCPN1009_n_28439), .o(n_28440) );
in01f80 g745218 ( .a(n_35648), .o(n_34593) );
in01f80 FE_OCP_DRV_C3740_n_29576 ( .a(n_29576), .o(FE_OCP_DRV_N3740_n_29576) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_7_ ( .ck(newNet_690), .d(n_46163), .o(delay_xor_ln21_unr6_stage3_stallmux_q_7_) );
in01f80 newInst_14 ( .a(tau_clk), .o(newNet_14) );
na02f80 g780924 ( .a(n_457), .b(n_516), .o(n_530) );
ao12f80 g770300 ( .a(FE_OCP_RBN2794_n_10106), .b(n_10406), .c(n_10484), .o(n_10507) );
no02f80 g760583 ( .a(n_19886), .b(FE_OFN816_n_19885), .o(n_19919) );
na02f80 g745372 ( .a(FE_OCP_RBN2987_n_35539), .b(n_35800), .o(n_35891) );
ao22s80 FE_RC_4127_0 ( .a(n_30770), .b(n_30777), .c(n_30769), .d(n_30776), .o(n_30918) );
in01f80 newInst_1270 ( .a(newNet_1269), .o(newNet_1270) );
in01f80 g777678 ( .a(n_4905), .o(n_3524) );
no02f80 g743283 ( .a(n_36725), .b(n_36743), .o(n_36761) );
in01f80 newInst_2409 ( .a(newNet_2408), .o(newNet_2409) );
na02f80 g761194 ( .a(n_19991), .b(n_19959), .o(n_21098) );
na02f80 g746991 ( .a(n_34075), .b(n_33667), .o(n_34081) );
in01f80 g762400 ( .a(n_18444), .o(n_18445) );
ao12f80 g762997 ( .a(n_17370), .b(n_17905), .c(n_17299), .o(n_17987) );
in01f80 g761272 ( .a(n_19956), .o(n_19957) );
na02f80 g775986 ( .a(n_5036), .b(n_5048), .o(n_5127) );
ao12f80 g753536 ( .a(n_26586), .b(n_26705), .c(n_26532), .o(n_26788) );
no02f80 g738615 ( .a(n_41361), .b(n_41368), .o(n_41390) );
no02f80 g753187 ( .a(n_27204), .b(FE_OCPN3186_FE_OCP_RBN1140_n_25816), .o(n_27346) );
in01f80 g755605 ( .a(n_24510), .o(n_24528) );
na02f80 FE_RC_3945_0 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_8_), .b(n_28273), .o(FE_RN_1706_0) );
na02f80 g762355 ( .a(n_45120), .b(n_18448), .o(n_18495) );
no02f80 g751192 ( .a(n_29818), .b(n_29311), .o(n_29886) );
na02f80 g739965 ( .a(n_39929), .b(n_39796), .o(n_39961) );
na02f80 g755398 ( .a(n_24765), .b(n_24764), .o(n_24784) );
oa22f80 FE_RC_1718_0 ( .a(n_24059), .b(n_27686), .c(n_27845), .d(n_27662), .o(n_27725) );
na02f80 g765204 ( .a(n_15302), .b(n_15299), .o(n_15341) );
in01f80 newInst_2321 ( .a(newNet_2320), .o(newNet_2321) );
in01f80 newInst_583 ( .a(newNet_276), .o(newNet_583) );
ao12f80 g755314 ( .a(n_24880), .b(n_24879), .c(n_24878), .o(n_26528) );
na02f80 g743926 ( .a(n_35750), .b(n_44221), .o(n_35868) );
in01f80 newInst_2296 ( .a(newNet_2295), .o(newNet_2296) );
ao12f80 g749267 ( .a(n_31527), .b(n_32063), .c(n_31571), .o(n_32152) );
in01f80 FE_OCP_RBC2548_n_44944 ( .a(n_44944), .o(FE_OCP_RBN2548_n_44944) );
oa22f80 g768520 ( .a(n_12267), .b(n_11939), .c(n_12333), .d(n_11938), .o(n_12350) );
in01f80 newInst_1739 ( .a(newNet_1738), .o(newNet_1739) );
in01f80 g760316 ( .a(n_20325), .o(n_21901) );
in01f80 newInst_39 ( .a(newNet_38), .o(newNet_39) );
no02f80 g778154 ( .a(n_2783), .b(n_2536), .o(n_2891) );
no02f80 g773216 ( .a(n_7743), .b(n_7945), .o(n_7962) );
in01f80 newInst_2858 ( .a(newNet_2127), .o(newNet_2858) );
ao22s80 g760808 ( .a(n_19393), .b(n_18591), .c(n_19479), .d(n_18592), .o(n_19538) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_29_ ( .ck(newNet_3502), .d(n_22902), .o(delay_add_ln22_unr14_stage6_stallmux_q_29_) );
in01f80 newInst_1337 ( .a(newNet_1336), .o(newNet_1337) );
no02f80 g743751 ( .a(n_37305), .b(n_37304), .o(n_37306) );
na02f80 g772829 ( .a(n_7985), .b(n_7907), .o(n_8095) );
in01f80 g754308 ( .a(n_25954), .o(n_25955) );
na02f80 g753674 ( .a(n_26524), .b(n_26363), .o(n_26630) );
in01f80 FE_OCP_RBC3422_n_12879 ( .a(n_12879), .o(FE_OCP_RBN3422_n_12879) );
oa12f80 g768812 ( .a(n_11648), .b(n_11929), .c(n_11631), .o(n_12030) );
oa12f80 g744007 ( .a(n_35523), .b(n_35537), .c(n_35522), .o(n_35557) );
na02f80 g780881 ( .a(n_420), .b(n_439), .o(n_488) );
in01f80 g754738 ( .a(n_26381), .o(n_26382) );
na02f80 g770557 ( .a(n_10326), .b(n_44463), .o(n_10362) );
in01f80 g763858 ( .a(n_17602), .o(n_17603) );
in01f80 newInst_3027 ( .a(newNet_3026), .o(newNet_3027) );
na02f80 g775975 ( .a(n_5216), .b(n_5154), .o(n_5520) );
in01f80 g773464 ( .a(n_7511), .o(n_7512) );
oa22f80 g784339 ( .a(FE_OFN775_n_46137), .b(n_5489), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5527), .o(n_46145) );
na02f80 FE_RC_2862_0 ( .a(n_13469), .b(n_14233), .o(FE_RN_1233_0) );
na02f80 g747254 ( .a(n_32773), .b(delay_add_ln22_unr20_stage8_stallmux_q_2_), .o(n_32786) );
na02f80 g766792 ( .a(FE_OCP_RBN3481_n_13667), .b(FE_OCP_RBN2244_n_13017), .o(n_13706) );
in01f80 newInst_810 ( .a(newNet_228), .o(newNet_810) );
no02f80 g736434 ( .a(n_43768), .b(n_43435), .o(n_43800) );
no02f80 g754542 ( .a(n_26633), .b(n_26572), .o(n_26711) );
in01f80 g768492 ( .a(n_12353), .o(n_12354) );
no02f80 g756323 ( .a(n_24587), .b(n_24543), .o(n_24544) );
in01f80 newInst_2745 ( .a(newNet_2744), .o(newNet_2745) );
oa12f80 g784680 ( .a(n_3949), .b(n_3948), .c(n_3920), .o(n_47010) );
na02f80 g779132 ( .a(n_1922), .b(n_1784), .o(n_1987) );
na02f80 g750504 ( .a(n_29518), .b(FE_OFN788_n_25834), .o(n_29603) );
ao12f80 g745090 ( .a(n_34437), .b(n_34661), .c(n_34267), .o(n_34795) );
na02f80 FE_RC_2659_0 ( .a(n_8213), .b(FE_RN_1111_0), .o(n_8243) );
na02f80 g753284 ( .a(n_27110), .b(n_26398), .o(n_27376) );
in01f80 g742243 ( .a(n_38179), .o(n_38180) );
na02f80 FE_RC_2460_0 ( .a(FE_RN_986_0), .b(n_14139), .o(n_14217) );
in01f80 g745437 ( .a(n_35796), .o(n_35797) );
na02f80 g777773 ( .a(n_3347), .b(n_2913), .o(n_3368) );
na02f80 g764642 ( .a(n_15775), .b(n_15743), .o(n_15915) );
in01f80 g743411 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .o(n_36591) );
in01f80 g742535 ( .a(n_37760), .o(n_37622) );
na02f80 g767817 ( .a(n_12753), .b(n_12799), .o(n_12849) );
ao12f80 g754877 ( .a(n_25186), .b(n_25185), .c(n_25184), .o(n_26850) );
in01f80 g774253 ( .a(n_6818), .o(n_6819) );
in01f80 fopt783922 ( .a(n_33492), .o(n_45627) );
in01f80 g773172 ( .a(n_7858), .o(n_7841) );
in01f80 g769784 ( .a(n_11238), .o(n_11239) );
oa12f80 g755782 ( .a(n_25061), .b(n_25060), .c(n_25059), .o(n_26162) );
oa22f80 FE_RC_1454_0 ( .a(n_22801), .b(n_22640), .c(n_22833), .d(n_22617), .o(n_22716) );
oa12f80 g779409 ( .a(n_1781), .b(n_1493), .c(FE_OCPN946_n_1780), .o(n_1782) );
na02f80 g764490 ( .a(n_16122), .b(n_14524), .o(n_16157) );
in01f80 newInst_2041 ( .a(newNet_2040), .o(newNet_2041) );
no02f80 g758230 ( .a(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .o(n_22729) );
na02f80 g780466 ( .a(n_1109), .b(n_1108), .o(n_1110) );
in01f80 g739473 ( .a(n_40753), .o(n_40754) );
in01f80 g738664 ( .a(n_41393), .o(n_41387) );
in01f80 newInst_2147 ( .a(newNet_2146), .o(newNet_2147) );
in01f80 g763172 ( .a(n_17459), .o(n_17441) );
no02f80 g742051 ( .a(FE_OCP_RBN2257_n_37844), .b(n_37544), .o(n_37946) );
in01f80 g770825 ( .a(n_10174), .o(n_10175) );
na03f80 g738202 ( .a(n_41941), .b(n_41924), .c(n_41785), .o(n_41976) );
no02f80 g752339 ( .a(n_44761), .b(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .o(n_27936) );
no02f80 g748255 ( .a(n_30465), .b(n_31783), .o(n_31868) );
ao22s80 g771036 ( .a(n_9511), .b(n_9413), .c(n_9510), .d(n_9414), .o(n_9682) );
na02f80 g740720 ( .a(n_39450), .b(n_39190), .o(n_39418) );
in01f80 g773428 ( .a(n_7555), .o(n_7556) );
ao22s80 g779312 ( .a(FE_OCP_RBN2160_n_1675), .b(n_1474), .c(n_1675), .d(n_1475), .o(n_1727) );
in01f80 g755093 ( .a(n_25147), .o(n_25209) );
no02f80 FE_RC_2258_0 ( .a(n_27899), .b(FE_RN_834_0), .o(FE_RN_835_0) );
in01f80 g751973 ( .a(n_28943), .o(n_28898) );
na02f80 g768601 ( .a(n_12232), .b(delay_add_ln22_unr8_stage4_stallmux_q_7_), .o(n_12313) );
no02f80 g748687 ( .a(n_31207), .b(n_31206), .o(n_31269) );
no02f80 g763580 ( .a(n_16893), .b(n_16936), .o(n_16937) );
in01f80 fopt783669 ( .a(n_5031), .o(n_45319) );
na02f80 g784606 ( .a(n_26727), .b(n_26620), .o(n_46934) );
in01f80 newInst_3261 ( .a(newNet_3260), .o(newNet_3261) );
no02f80 g762035 ( .a(n_18593), .b(n_18541), .o(n_18591) );
no02f80 FE_RC_1363_0 ( .a(FE_RN_405_0), .b(FE_RN_406_0), .o(FE_RN_407_0) );
ao12f80 g737948 ( .a(FE_OCPN936_n_42192), .b(n_42212), .c(n_42191), .o(n_42497) );
no02f80 FE_RC_2515_0 ( .a(n_27131), .b(n_31107), .o(FE_RN_1023_0) );
na02f80 g766501 ( .a(n_14065), .b(n_14064), .o(n_14066) );
no02f80 g737503 ( .a(n_42649), .b(n_42664), .o(n_43037) );
no02f80 g772232 ( .a(n_8734), .b(n_8144), .o(n_8852) );
no02f80 g756164 ( .a(n_24163), .b(n_23764), .o(n_24203) );
na02f80 FE_RC_3051_0 ( .a(n_35312), .b(n_35379), .o(FE_RN_1337_0) );
in01f80 FE_OCPC978_n_21973 ( .a(n_21973), .o(FE_OCPN978_n_21973) );
no02f80 FE_RC_4227_0 ( .a(FE_RN_1852_0), .b(FE_RN_1855_0), .o(n_30405) );
no02f80 g744039 ( .a(n_44221), .b(n_35667), .o(n_35755) );
in01f80 FE_RC_4248_0 ( .a(FE_OCPN1771_n_26801), .o(FE_RN_1869_0) );
in01f80 g750944 ( .a(n_29030), .o(n_29053) );
no02f80 g764874 ( .a(n_16137), .b(n_16138), .o(n_16139) );
in01f80 g737901 ( .a(n_42225), .o(n_42226) );
in01f80 g747461 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n_33155) );
ao12f80 g745954 ( .a(n_34062), .b(n_34061), .c(n_34060), .o(n_35315) );
in01f80 newInst_1130 ( .a(newNet_1129), .o(newNet_1130) );
in01f80 newInst_815 ( .a(newNet_393), .o(newNet_815) );
ao12f80 g757459 ( .a(n_23227), .b(n_44084), .c(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .o(n_23011) );
na02f80 g738533 ( .a(n_41425), .b(n_41174), .o(n_41450) );
na02f80 g766224 ( .a(n_14372), .b(FE_OCP_RBN1147_n_13098), .o(n_14510) );
no02f80 g739909 ( .a(n_40374), .b(n_40154), .o(n_40375) );
na02f80 g751843 ( .a(n_29124), .b(n_29123), .o(n_29125) );
in01f80 FE_OCP_DRV_C1578_n_33904 ( .a(FE_OCP_DRV_N1577_n_33904), .o(FE_OCP_DRV_N1578_n_33904) );
no02f80 g760777 ( .a(n_19536), .b(n_19511), .o(n_19596) );
no02f80 g749802 ( .a(n_31510), .b(n_31509), .o(n_31534) );
na02f80 g764253 ( .a(n_16402), .b(n_16374), .o(n_16440) );
ao12f80 g758155 ( .a(n_22846), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n_23148) );
no02f80 FE_RC_1728_0 ( .a(n_23371), .b(n_23361), .o(FE_RN_479_0) );
na02f80 g772949 ( .a(n_7834), .b(n_7701), .o(n_7887) );
in01f80 FE_OCP_RBC1154_n_18375 ( .a(n_18375), .o(FE_OCP_RBN1154_n_18375) );
no02f80 g768264 ( .a(n_12623), .b(n_12279), .o(n_12663) );
na02f80 g761355 ( .a(n_19054), .b(FE_OCP_DRV_N1550_n_19053), .o(n_19072) );
na02f80 g778382 ( .a(n_2502), .b(n_2898), .o(n_2507) );
oa12f80 g777739 ( .a(n_3317), .b(n_3318), .c(n_3319), .o(n_3343) );
no02f80 g766754 ( .a(n_14085), .b(n_13902), .o(n_14139) );
no02f80 g762314 ( .a(n_18047), .b(n_18004), .o(n_18093) );
in01f80 FE_RC_2062_0 ( .a(n_35012), .o(FE_RN_699_0) );
oa12f80 g738427 ( .a(n_41729), .b(n_41537), .c(n_41615), .o(n_41770) );
in01f80 g744997 ( .a(n_35659), .o(n_34989) );
ao12f80 g757470 ( .a(n_23358), .b(n_23357), .c(n_23356), .o(n_23901) );
na02f80 g738415 ( .a(n_41635), .b(n_41634), .o(n_41636) );
in01f80 g755770 ( .a(n_24432), .o(n_24433) );
in01f80 g736905 ( .a(n_43577), .o(n_43578) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_20_ ( .ck(newNet_1744), .d(n_22521), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_20_) );
in01f80 newInst_1128 ( .a(newNet_1127), .o(newNet_1128) );
na02f80 g763374 ( .a(n_16986), .b(n_16948), .o(n_17081) );
in01f80 newInst_1525 ( .a(newNet_504), .o(newNet_1525) );
na02f80 g740908 ( .a(n_39309), .b(n_39341), .o(n_39460) );
no02f80 g770112 ( .a(n_10769), .b(n_10290), .o(n_10808) );
oa12f80 g777791 ( .a(n_3245), .b(n_3287), .c(n_3286), .o(n_3296) );
no02f80 g749890 ( .a(n_29871), .b(n_29847), .o(n_31490) );
no02f80 FE_RC_2220_0 ( .a(n_32949), .b(n_32914), .o(FE_RN_803_0) );
no02f80 FE_RC_1830_0 ( .a(FE_RN_547_0), .b(FE_RN_549_0), .o(n_16972) );
na02f80 g780823 ( .a(n_409), .b(n_408), .o(n_410) );
oa12f80 g743530 ( .a(n_36008), .b(n_36474), .c(n_47265), .o(n_36506) );
in01f80 g776400 ( .a(n_4396), .o(n_4466) );
in01f80 FE_OCP_RBC1837_FE_RN_1542_0 ( .a(FE_RN_1542_0), .o(FE_OCP_RBN1837_FE_RN_1542_0) );
in01f80 g745619 ( .a(n_34564), .o(n_34537) );
oa22f80 FE_RC_947_0 ( .a(n_20231), .b(n_22874), .c(n_20252), .d(n_44327), .o(n_22947) );
in01f80 newInst_1769 ( .a(newNet_1768), .o(newNet_1769) );
in01f80 g760967 ( .a(n_19280), .o(n_19281) );
na02f80 g772219 ( .a(n_8622), .b(n_8668), .o(n_8765) );
in01f80 FE_OCP_RBC1698_n_19353 ( .a(n_19353), .o(FE_OCP_RBN1698_n_19353) );
na02f80 g768002 ( .a(n_12616), .b(n_12666), .o(n_12667) );
in01f80 g768101 ( .a(n_12816), .o(n_12817) );
ao12f80 g769071 ( .a(n_11972), .b(n_12016), .c(n_11794), .o(n_12051) );
na02f80 g768598 ( .a(n_12261), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_), .o(n_12309) );
na02f80 g751591 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .o(n_28543) );
no02f80 g761641 ( .a(n_18683), .b(n_18652), .o(n_18797) );
no02f80 g746084 ( .a(n_35163), .b(n_35162), .o(n_35164) );
in01f80 FE_OCP_RBC2662_n_20333 ( .a(n_20333), .o(FE_OCP_RBN2662_n_20333) );
in01f80 g763694 ( .a(n_16759), .o(n_16832) );
no02f80 g761550 ( .a(n_19542), .b(n_19541), .o(n_19543) );
na02f80 g753891 ( .a(n_26297), .b(FE_OCPN1528_n_26296), .o(n_26325) );
in01f80 newInst_616 ( .a(newNet_615), .o(newNet_616) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_3_ ( .ck(newNet_2061), .d(n_4793), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_) );
na02f80 FE_RC_3928_0 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .b(FE_OCP_RBN3331_n_44962), .o(FE_RN_1699_0) );
ao12f80 g756823 ( .a(n_23245), .b(n_23420), .c(n_23289), .o(n_23458) );
no02f80 g757302 ( .a(n_23468), .b(n_22978), .o(n_23495) );
in01f80 newInst_3 ( .a(tau_clk), .o(newNet_3) );
in01f80 g757688 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .o(n_22630) );
in01f80 newInst_2540 ( .a(newNet_2539), .o(newNet_2540) );
no02f80 g757007 ( .a(n_23251), .b(n_23250), .o(n_23408) );
no02f80 g755575 ( .a(n_24626), .b(n_24368), .o(n_24574) );
na02f80 g769601 ( .a(n_11320), .b(FE_OCP_RBN2845_n_10326), .o(n_11318) );
oa22f80 g740955 ( .a(n_39065), .b(n_38895), .c(n_38971), .d(n_38896), .o(n_39112) );
oa12f80 g757582 ( .a(n_22888), .b(n_23243), .c(n_23295), .o(n_23343) );
no02f80 g740196 ( .a(FE_OCP_RBN3722_n_39913), .b(n_40177), .o(n_40214) );
no02f80 g769249 ( .a(n_11475), .b(FE_OCP_RBN2891_n_10568), .o(n_11497) );
in01f80 g752596 ( .a(n_27630), .o(n_27631) );
in01f80 g771117 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n_11879) );
in01f80 newInst_3180 ( .a(newNet_3179), .o(newNet_3180) );
na02f80 g738948 ( .a(n_41159), .b(n_40911), .o(n_41195) );
in01f80 g737331 ( .a(n_43181), .o(n_42883) );
in01f80 newInst_1895 ( .a(newNet_1894), .o(newNet_1895) );
in01f80 newInst_1119 ( .a(newNet_1118), .o(newNet_1119) );
na03f80 g748721 ( .a(n_32426), .b(n_32556), .c(n_32555), .o(n_32557) );
no02f80 g776081 ( .a(n_4928), .b(n_4292), .o(n_5080) );
in01f80 g758266 ( .a(n_22643), .o(n_22644) );
in01f80 g740732 ( .a(n_40009), .o(n_39580) );
na02f80 g740688 ( .a(n_39969), .b(n_39538), .o(n_39539) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_28_ ( .ck(newNet_309), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_28_) );
no02f80 g750644 ( .a(n_29376), .b(FE_OCPUNCON1802_n_29375), .o(n_29443) );
na02f80 g764362 ( .a(n_16205), .b(n_16206), .o(n_16207) );
in01f80 g745253 ( .a(n_35681), .o(n_35682) );
in01f80 g773149 ( .a(n_7909), .o(n_7910) );
in01f80 g737631 ( .a(n_42698), .o(n_42699) );
oa22f80 FE_RC_1459_0 ( .a(n_22801), .b(n_22684), .c(n_22833), .d(n_22637), .o(n_22758) );
in01f80 FE_OCP_RBC3099_n_32001 ( .a(n_32001), .o(FE_OCP_RBN3099_n_32001) );
in01f80 newInst_3291 ( .a(newNet_3290), .o(newNet_3291) );
in01f80 newInst_36 ( .a(newNet_35), .o(newNet_36) );
no02f80 g763311 ( .a(n_16910), .b(n_16868), .o(n_17005) );
in01f80 FE_RC_363_0 ( .a(n_176), .o(FE_RN_109_0) );
oa12f80 g760347 ( .a(n_20811), .b(n_20835), .c(n_20810), .o(n_20894) );
no02f80 g753688 ( .a(n_26523), .b(n_25014), .o(n_26766) );
na02f80 g742639 ( .a(n_37465), .b(n_37464), .o(n_37466) );
in01f80 newInst_3691 ( .a(newNet_3690), .o(newNet_3691) );
oa12f80 g773723 ( .a(n_7243), .b(n_7264), .c(n_7242), .o(n_7801) );
no02f80 g779559 ( .a(n_1456), .b(n_1408), .o(n_1501) );
na02f80 g755749 ( .a(n_25219), .b(n_25161), .o(n_25343) );
no02f80 g748795 ( .a(n_32409), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n_32493) );
na02f80 g746135 ( .a(n_35653), .b(n_35125), .o(n_35189) );
na02f80 g775457 ( .a(n_46999), .b(FE_OCP_RBN2767_n_4376), .o(n_5824) );
no02f80 g745538 ( .a(n_34535), .b(n_34484), .o(n_34536) );
in01f80 g752932 ( .a(n_28076), .o(n_28154) );
in01f80 g737482 ( .a(n_42600), .o(n_42637) );
in01f80 g752383 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .o(n_28606) );
na02f80 g777142 ( .a(n_3629), .b(n_3679), .o(n_3837) );
na02f80 g765824 ( .a(n_14918), .b(n_14843), .o(n_14974) );
in01f80 FE_OCPC1519_n_31403 ( .a(n_31403), .o(FE_OCPN1519_n_31403) );
in01f80 g771098 ( .a(n_9666), .o(n_9667) );
oa12f80 g770525 ( .a(n_10174), .b(n_10498), .c(n_10257), .o(n_10572) );
in01f80 g737297 ( .a(n_42924), .o(n_42925) );
na02f80 g740655 ( .a(n_39597), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39637) );
no02f80 g750736 ( .a(n_29218), .b(n_28725), .o(n_29236) );
no02f80 g748014 ( .a(n_31975), .b(n_31837), .o(n_32060) );
in01f80 g742994 ( .a(n_36964), .o(n_36965) );
no02f80 g746925 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_), .o(n_32962) );
no02f80 g761811 ( .a(n_18379), .b(n_18244), .o(n_18380) );
in01f80 FE_OCP_RBC3525_n_29624 ( .a(n_29624), .o(FE_OCP_RBN3525_n_29624) );
in01f80 g742960 ( .a(n_37056), .o(n_37057) );
in01f80 newInst_2433 ( .a(newNet_2432), .o(newNet_2433) );
no02f80 g771820 ( .a(n_9547), .b(n_9433), .o(n_9548) );
in01f80 g778705 ( .a(n_2383), .o(n_2384) );
na02f80 g747873 ( .a(FE_OCP_RBN1212_n_32142), .b(n_31861), .o(n_32216) );
no02f80 g743945 ( .a(n_35984), .b(n_47266), .o(n_36099) );
ao12f80 g763047 ( .a(n_17904), .b(n_17903), .c(n_17902), .o(n_18494) );
in01f80 newInst_698 ( .a(newNet_697), .o(newNet_698) );
in01f80 g771335 ( .a(n_9374), .o(n_9375) );
no03m80 g746716 ( .a(n_34211), .b(n_34234), .c(n_33792), .o(n_34330) );
oa12f80 g742265 ( .a(n_37820), .b(n_37819), .c(n_37818), .o(n_38731) );
ao12f80 g752665 ( .a(n_28137), .b(n_28136), .c(n_28135), .o(n_28856) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_7_ ( .ck(newNet_1942), .d(n_10490), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_7_) );
no02f80 FE_RC_2044_0 ( .a(FE_RN_684_0), .b(FE_RN_685_0), .o(FE_RN_686_0) );
na02f80 g743134 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .o(n_37145) );
no02f80 g740416 ( .a(n_39942), .b(n_39496), .o(n_40130) );
in01f80 g763192 ( .a(n_17399), .o(n_17400) );
in01f80 g748191 ( .a(n_31506), .o(n_31524) );
in01f80 newInst_2749 ( .a(newNet_580), .o(newNet_2749) );
oa12f80 g778444 ( .a(n_2882), .b(n_2878), .c(n_3029), .o(n_3525) );
na02f80 g736571 ( .a(n_43682), .b(n_43424), .o(n_43684) );
no02f80 g744143 ( .a(n_35821), .b(n_35820), .o(n_35859) );
in01f80 newInst_411 ( .a(newNet_410), .o(newNet_411) );
na02f80 FE_RC_1312_0 ( .a(FE_RN_384_0), .b(FE_RN_385_0), .o(FE_RN_386_0) );
in01f80 FE_OCP_RBC2414_n_2922 ( .a(n_2922), .o(FE_OCP_RBN2414_n_2922) );
in01f80 newInst_2963 ( .a(newNet_2962), .o(newNet_2963) );
no02f80 g765317 ( .a(n_15156), .b(FE_OCP_RBN3509_n_13860), .o(n_15270) );
na02f80 g741053 ( .a(n_39422), .b(n_39487), .o(n_39504) );
in01f80 FE_OFC780_n_17093 ( .a(FE_OFN777_n_17093), .o(FE_OFN780_n_17093) );
na02f80 g779148 ( .a(n_1921), .b(n_1785), .o(n_1922) );
in01f80 newInst_3124 ( .a(newNet_127), .o(newNet_3124) );
na02f80 g777865 ( .a(n_3263), .b(n_3277), .o(n_3362) );
na02f80 g743046 ( .a(n_37145), .b(n_37037), .o(n_37176) );
in01f80 g739887 ( .a(n_40345), .o(n_40346) );
in01f80 g736389 ( .a(n_43840), .o(n_43841) );
na02f80 g737439 ( .a(n_42717), .b(n_42426), .o(n_42749) );
oa22f80 FE_RC_1693_0 ( .a(n_25586), .b(FE_OCP_RBN2765_n_25895), .c(n_25585), .d(n_25895), .o(n_25986) );
na02f80 g764265 ( .a(n_16394), .b(n_16436), .o(n_16437) );
in01f80 g758677 ( .a(n_21813), .o(n_21814) );
in01f80 FE_OCP_RBC3096_n_43489 ( .a(n_43489), .o(FE_OCP_RBN3096_n_43489) );
in01f80 newInst_1069 ( .a(newNet_1068), .o(newNet_1069) );
na02f80 g743564 ( .a(n_36446), .b(n_36246), .o(n_36490) );
in01f80 newInst_2413 ( .a(newNet_2412), .o(newNet_2413) );
na02f80 g739294 ( .a(n_40876), .b(n_40875), .o(n_40877) );
no02f80 g744271 ( .a(n_44174), .b(n_34870), .o(n_35616) );
no03m80 g779435 ( .a(n_1512), .b(n_1443), .c(n_1508), .o(n_1597) );
na02f80 FE_RC_2964_0 ( .a(n_10760), .b(FE_RN_1294_0), .o(n_10827) );
no02f80 g774829 ( .a(n_6228), .b(FE_OCP_RBN2975_n_5531), .o(n_6287) );
no02f80 g766992 ( .a(n_13767), .b(n_13766), .o(n_13768) );
in01f80 g742498 ( .a(n_37662), .o(n_37796) );
na02f80 g775961 ( .a(n_5181), .b(n_4507), .o(n_5234) );
na02f80 g754337 ( .a(n_26646), .b(n_26312), .o(n_26688) );
no02f80 g743526 ( .a(n_36462), .b(n_36000), .o(n_36508) );
no03m80 g743272 ( .a(n_38021), .b(n_37858), .c(n_37920), .o(n_38022) );
no02f80 g775866 ( .a(FE_OCP_RBN2727_n_4219), .b(n_4923), .o(n_5050) );
no02f80 g754959 ( .a(n_25156), .b(n_25182), .o(n_25214) );
in01f80 g771594 ( .a(n_10385), .o(n_10386) );
in01f80 FE_RC_3662_0 ( .a(FE_OCPN856_n_20367), .o(FE_RN_1608_0) );
oa12f80 g778294 ( .a(n_2555), .b(n_2554), .c(FE_OCP_RBN2267_n_2430), .o(n_4280) );
oa12f80 g780795 ( .a(n_472), .b(n_469), .c(n_462), .o(n_496) );
no04s80 FE_RC_1195_0 ( .a(n_32962), .b(n_33023), .c(n_32961), .d(n_32976), .o(n_33024) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_15_ ( .ck(newNet_1538), .d(n_32093), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_) );
oa12f80 g753804 ( .a(n_26427), .b(n_26426), .c(n_26425), .o(n_26491) );
in01f80 FE_OCP_RBC3451_n_37945 ( .a(FE_OCP_RBN3447_n_37945), .o(FE_OCP_RBN3451_n_37945) );
na02f80 FE_RC_2632_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .b(FE_OCP_RBN2117_n_45224), .o(FE_RN_1096_0) );
na02f80 g765527 ( .a(n_15599), .b(n_15712), .o(n_15922) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_29_ ( .ck(newNet_1295), .d(n_44624), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
oa12f80 g758004 ( .a(n_22725), .b(n_22917), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n_22922) );
no02f80 FE_RC_1948_0 ( .a(n_25786), .b(FE_RN_623_0), .o(FE_RN_624_0) );
na02f80 g780930 ( .a(n_357), .b(n_372), .o(n_373) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_11_ ( .ck(newNet_1547), .d(n_32005), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_) );
ao12f80 g752607 ( .a(n_28246), .b(n_28245), .c(n_28244), .o(n_28860) );
oa22f80 g779243 ( .a(n_1725), .b(n_1564), .c(n_1786), .d(n_1563), .o(n_1837) );
in01f80 FE_RC_2957_0 ( .a(n_11370), .o(FE_RN_1291_0) );
na02f80 g744509 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n_36727) );
no02f80 g770817 ( .a(n_9908), .b(n_9928), .o(n_9934) );
in01f80 FE_OFC221_n_35655 ( .a(FE_OFN220_n_35655), .o(FE_OFN221_n_35655) );
no02f80 g738077 ( .a(n_42075), .b(n_42098), .o(n_42128) );
no02f80 g741168 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39232), .o(n_39244) );
no02f80 g766593 ( .a(n_13988), .b(n_14019), .o(n_14020) );
in01f80 newInst_3460 ( .a(newNet_3459), .o(newNet_3460) );
na02f80 g750781 ( .a(n_29258), .b(FE_OCP_RBN1143_n_29292), .o(n_29259) );
in01f80 FE_OCPC3757_n_13889 ( .a(FE_OCPN3756_n_13889), .o(FE_OCPN3757_n_13889) );
no02f80 g780908 ( .a(n_403), .b(n_437), .o(n_478) );
oa22f80 g779223 ( .a(n_1812), .b(n_1610), .c(n_1807), .d(n_1609), .o(n_1898) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_25_ ( .ck(newNet_225), .d(n_46193), .o(delay_xor_ln22_unr6_stage3_stallmux_q_25_) );
na02f80 g752232 ( .a(n_27871), .b(FE_OCP_RBN3308_n_44722), .o(n_27872) );
in01f80 FE_RC_2109_0 ( .a(n_31014), .o(FE_RN_730_0) );
in01f80 g752598 ( .a(n_27628), .o(n_27629) );
na02f80 g780802 ( .a(n_386), .b(n_382), .o(n_383) );
in01f80 g773189 ( .a(n_7627), .o(n_7641) );
no02f80 g778344 ( .a(n_2607), .b(n_2606), .o(n_2636) );
in01f80 g738280 ( .a(n_41947), .o(n_42478) );
in01f80 g773215 ( .a(n_7962), .o(n_8031) );
no02f80 g780765 ( .a(n_505), .b(n_391), .o(n_506) );
in01f80 newInst_485 ( .a(newNet_132), .o(newNet_485) );
in01f80 g767907 ( .a(n_12690), .o(n_12691) );
in01f80 g741088 ( .a(n_39002), .o(n_39107) );
in01f80 g760611 ( .a(n_19862), .o(n_19888) );
na02f80 g768637 ( .a(n_12254), .b(n_12209), .o(n_12255) );
no02f80 g766716 ( .a(n_13775), .b(n_13808), .o(n_13918) );
in01f80 FE_OFC820_n_4333 ( .a(FE_OFN835_n_4333), .o(FE_OFN820_n_4333) );
oa12f80 g768943 ( .a(n_11525), .b(n_11775), .c(n_11607), .o(n_11835) );
na02f80 g764267 ( .a(n_16452), .b(n_16455), .o(n_16513) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_26_ ( .ck(newNet_1389), .d(n_36698), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_) );
no02f80 g766394 ( .a(n_14131), .b(n_14129), .o(n_14185) );
no02f80 g764879 ( .a(n_15687), .b(n_15686), .o(n_15725) );
no02f80 g776848 ( .a(n_4176), .b(n_4222), .o(n_4254) );
na02f80 FE_RC_1325_0 ( .a(FE_RN_392_0), .b(n_9869), .o(n_10181) );
no02f80 g777384 ( .a(n_3507), .b(n_3363), .o(n_3508) );
in01f80 FE_OCP_RBC3594_n_44561 ( .a(FE_OCP_RBN2616_n_44561), .o(FE_OCP_RBN3594_n_44561) );
oa22f80 g738841 ( .a(n_41258), .b(n_40953), .c(n_41259), .d(n_40952), .o(n_41313) );
ao22s80 FE_RC_421_0 ( .a(n_14758), .b(FE_OCP_RBN2652_n_14684), .c(FE_OCP_RBN2507_n_13896), .d(n_14684), .o(n_14785) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_12_ ( .ck(newNet_1766), .d(n_22031), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_) );
no02f80 g776939 ( .a(n_3973), .b(n_47022), .o(n_4019) );
in01f80 g752481 ( .a(n_27723), .o(n_27724) );
na02f80 g773689 ( .a(n_7275), .b(n_7106), .o(n_7346) );
no02f80 g769199 ( .a(n_11896), .b(n_11895), .o(n_12513) );
in01f80 newInst_3551 ( .a(newNet_3550), .o(newNet_3551) );
no02f80 g746347 ( .a(n_33607), .b(n_33606), .o(n_33608) );
oa22f80 g773808 ( .a(n_7072), .b(n_7034), .c(n_7101), .d(n_7035), .o(n_7156) );
no02f80 g772931 ( .a(n_7875), .b(n_7874), .o(n_7936) );
in01f80 g741529 ( .a(n_38740), .o(n_38741) );
in01f80 FE_RC_3072_0 ( .a(FE_RN_1352_0), .o(n_26519) );
no02f80 g769341 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .o(n_11631) );
in01f80 g748297 ( .a(n_31706), .o(n_31738) );
in01f80 g775564 ( .a(n_5608), .o(n_5641) );
in01f80 newInst_2309 ( .a(newNet_2308), .o(newNet_2309) );
in01f80 g767442 ( .a(n_13175), .o(n_13176) );
no02f80 g748932 ( .a(n_31082), .b(n_31108), .o(n_31109) );
oa12f80 g741771 ( .a(n_38403), .b(n_38425), .c(n_38402), .o(n_38572) );
ao12f80 g779473 ( .a(n_1881), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .o(n_2088) );
in01f80 newInst_1885 ( .a(newNet_1884), .o(newNet_1885) );
no02f80 g780460 ( .a(FE_OFN795_n_45813), .b(n_745), .o(n_846) );
in01f80 g766054 ( .a(n_14613), .o(n_14614) );
na02f80 g776600 ( .a(n_4241), .b(n_4133), .o(n_4391) );
na02f80 g759290 ( .a(FE_OCP_RBN1375_n_20889), .b(n_45091), .o(n_20948) );
na02f80 g736766 ( .a(n_43257), .b(n_43320), .o(n_43353) );
no02f80 FE_RC_2425_0 ( .a(FE_RN_959_0), .b(FE_RN_961_0), .o(FE_RN_962_0) );
in01f80 newInst_2708 ( .a(newNet_2707), .o(newNet_2708) );
na02f80 g758122 ( .a(n_44267), .b(n_21312), .o(n_22259) );
in01f80 g751607 ( .a(n_28815), .o(n_28816) );
no02f80 g775830 ( .a(n_5163), .b(n_4182), .o(n_5198) );
in01f80 fopt782962 ( .a(n_24990), .o(n_44423) );
in01f80 g743756 ( .a(n_36273), .o(n_36274) );
in01f80 g760520 ( .a(n_20020), .o(n_20021) );
in01f80 g749552 ( .a(n_30428), .o(n_31804) );
in01f80 g766359 ( .a(n_14362), .o(n_14363) );
in01f80 g745055 ( .a(n_34828), .o(n_34827) );
in01f80 FE_RC_1554_0 ( .a(n_8492), .o(FE_RN_439_0) );
in01f80 FE_OCP_RBC1688_n_18986 ( .a(FE_OCP_RBN1686_n_18986), .o(FE_OCP_RBN1688_n_18986) );
in01f80 g776573 ( .a(n_4449), .o(n_4450) );
no02f80 FE_RC_2270_0 ( .a(FE_RN_844_0), .b(n_25715), .o(n_25743) );
in01f80 g767002 ( .a(n_14211), .o(n_14338) );
na02f80 g763675 ( .a(n_16829), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n_16828) );
na02f80 g737882 ( .a(n_42201), .b(n_42309), .o(n_42362) );
in01f80 newInst_861 ( .a(newNet_780), .o(newNet_861) );
na02f80 g755345 ( .a(n_25410), .b(n_24997), .o(n_25409) );
na02f80 g740787 ( .a(n_39462), .b(n_39323), .o(n_39492) );
oa12f80 g736372 ( .a(n_349), .b(n_43771), .c(FE_OFN3_n_43918), .o(n_43805) );
na02f80 g773079 ( .a(n_7716), .b(n_7827), .o(n_8281) );
in01f80 g774960 ( .a(n_6149), .o(n_6150) );
no02f80 g749528 ( .a(n_30573), .b(n_30572), .o(n_30574) );
na02f80 g758940 ( .a(n_21606), .b(n_21644), .o(n_21645) );
no02f80 g754731 ( .a(n_26541), .b(n_26634), .o(n_26712) );
na02f80 g746002 ( .a(n_35243), .b(n_35242), .o(n_35244) );
in01f80 g779796 ( .a(n_1682), .o(n_1409) );
oa12f80 g751017 ( .a(n_29932), .b(n_30089), .c(n_30030), .o(n_30067) );
no02f80 g749740 ( .a(n_31225), .b(FE_OCP_RBN3012_n_31117), .o(n_31291) );
oa12f80 g739712 ( .a(n_40335), .b(n_40505), .c(n_40192), .o(n_40515) );
in01f80 newInst_3527 ( .a(newNet_3526), .o(newNet_3527) );
in01f80 g777953 ( .a(n_3717), .o(n_3715) );
no02f80 g777726 ( .a(n_3367), .b(n_3351), .o(n_3352) );
na02f80 g767806 ( .a(n_13119), .b(n_13017), .o(n_13236) );
na02f80 g763528 ( .a(FE_OCP_RBN3081_n_16977), .b(n_15816), .o(n_17164) );
na02f80 g779015 ( .a(n_2150), .b(n_2175), .o(n_2698) );
no02f80 g776234 ( .a(n_4550), .b(n_4549), .o(n_4602) );
in01f80 FE_OCPC1234_n_2414 ( .a(FE_OCPN1233_n_2414), .o(FE_OCPN1234_n_2414) );
no02f80 g770453 ( .a(n_10401), .b(n_44464), .o(n_10586) );
na02f80 g765570 ( .a(n_15142), .b(n_14364), .o(n_15330) );
no02f80 g752176 ( .a(n_44826), .b(n_28106), .o(n_28591) );
in01f80 g749243 ( .a(n_32114), .o(n_32115) );
in01f80 FE_OCPC3175_n_31125 ( .a(n_31125), .o(FE_OCPN3175_n_31125) );
in01f80 FE_RC_752_0 ( .a(n_27968), .o(FE_RN_235_0) );
oa12f80 g737739 ( .a(FE_OCPN885_n_42216), .b(n_42358), .c(n_42562), .o(n_42386) );
in01f80 newInst_2106 ( .a(newNet_2105), .o(newNet_2106) );
no02f80 g779601 ( .a(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_6_), .o(n_1450) );
in01f80 g761950 ( .a(n_18289), .o(n_18290) );
na02f80 g743916 ( .a(n_35578), .b(n_35577), .o(n_35579) );
in01f80 FE_OCP_RBC3076_FE_OFN807_n_46195 ( .a(FE_OFN807_n_46195), .o(FE_OCP_RBN3076_FE_OFN807_n_46195) );
no02f80 g777155 ( .a(n_4864), .b(n_4863), .o(n_4973) );
in01f80 newInst_3279 ( .a(newNet_3278), .o(newNet_3279) );
in01f80 g768368 ( .a(n_12577), .o(n_12578) );
ao12f80 g751774 ( .a(n_44045), .b(n_28941), .c(n_28793), .o(n_29050) );
in01f80 FE_OFC842_n_5067 ( .a(n_5067), .o(FE_OFN842_n_5067) );
ao22s80 g767835 ( .a(n_12787), .b(FE_OCP_RBN1925_cordic_combinational_sub_ln23_0_unr12_z_0__), .c(n_12786), .d(FE_OCP_RBN1923_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_13764) );
ao12f80 g759152 ( .a(n_21259), .b(n_21415), .c(n_21342), .o(n_21526) );
na02f80 g768924 ( .a(n_12213), .b(n_11968), .o(n_12220) );
no02f80 g753458 ( .a(n_26957), .b(n_26956), .o(n_26980) );
in01f80 g777565 ( .a(n_4182), .o(n_4219) );
no02f80 g768535 ( .a(n_12331), .b(n_12341), .o(n_12332) );
no02f80 g778033 ( .a(n_3035), .b(n_3626), .o(n_3065) );
in01f80 g758743 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_8_), .o(n_23267) );
in01f80 g777233 ( .a(n_3661), .o(n_3662) );
no02f80 g772597 ( .a(n_8284), .b(n_8147), .o(n_8325) );
oa22f80 FE_RC_1443_0 ( .a(n_28336), .b(n_44216), .c(n_32287), .d(n_32290), .o(n_32337) );
na02f80 g770325 ( .a(FE_OCP_RBN2886_n_10570), .b(FE_OCP_RBN2621_n_44561), .o(n_10617) );
in01f80 newInst_1462 ( .a(newNet_1461), .o(newNet_1462) );
ao12f80 g766403 ( .a(n_14567), .b(n_14566), .c(n_14565), .o(n_15666) );
ao22s80 FE_RC_3768_0 ( .a(n_17129), .b(n_16985), .c(n_16984), .d(n_16937), .o(n_17243) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_0_ ( .ck(newNet_2795), .d(n_14732), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_) );
no02f80 g745587 ( .a(n_34291), .b(n_33222), .o(n_34353) );
in01f80 g780338 ( .a(n_967), .o(n_1004) );
na02f80 g760710 ( .a(n_19693), .b(n_19661), .o(n_19738) );
in01f80 g753454 ( .a(n_27004), .o(n_27005) );
na02f80 g746769 ( .a(n_32892), .b(n_32946), .o(n_32978) );
ao12f80 g784612 ( .a(n_42874), .b(n_42848), .c(n_42612), .o(n_46940) );
no03m80 FE_RC_2557_0 ( .a(FE_OCPN1020_n_23078), .b(n_22998), .c(n_23044), .o(n_23175) );
no02f80 g769977 ( .a(n_11047), .b(n_10993), .o(n_11043) );
no02f80 g759617 ( .a(n_20684), .b(n_20371), .o(n_20685) );
in01f80 FE_OCP_RBC2205_n_18242 ( .a(FE_OCP_RBN2203_n_18242), .o(FE_OCP_RBN2205_n_18242) );
na02f80 g773801 ( .a(n_7145), .b(n_7062), .o(n_7222) );
in01f80 g756174 ( .a(n_24224), .o(n_24225) );
in01f80 FE_OCP_RBC2575_n_34822 ( .a(n_34822), .o(FE_OCP_RBN2575_n_34822) );
in01f80 newInst_3005 ( .a(newNet_145), .o(newNet_3005) );
ao12f80 g755669 ( .a(n_24449), .b(n_24503), .c(n_24502), .o(n_24568) );
in01f80 g737938 ( .a(n_42296), .o(n_42297) );
oa12f80 g773885 ( .a(n_6987), .b(n_7055), .c(n_6930), .o(n_7088) );
ao22s80 FE_RC_3241_0 ( .a(FE_OFN756_n_44461), .b(n_10225), .c(n_44463), .d(n_10202), .o(n_10401) );
no02f80 g770422 ( .a(n_10575), .b(n_10565), .o(n_10566) );
in01f80 g767064 ( .a(n_13897), .o(n_13967) );
na02f80 g768750 ( .a(n_11998), .b(n_11997), .o(n_11999) );
in01f80 g771740 ( .a(n_9006), .o(n_9007) );
na02f80 g778427 ( .a(n_2616), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .o(n_2663) );
in01f80 g766883 ( .a(n_14341), .o(n_14342) );
in01f80 g764472 ( .a(n_16361), .o(n_16386) );
na02f80 g750067 ( .a(n_29869), .b(n_46960), .o(n_30113) );
na02f80 g762285 ( .a(n_18579), .b(n_18578), .o(n_18968) );
oa22f80 FE_RC_2534_0 ( .a(n_36706), .b(n_36772), .c(n_36771), .d(n_36707), .o(n_36800) );
na02f80 g745366 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35720), .o(n_35849) );
ao12f80 g741001 ( .a(n_38974), .b(FE_OCP_RBN3580_n_44944), .c(n_38989), .o(n_39105) );
in01f80 newInst_1947 ( .a(newNet_1946), .o(newNet_1947) );
no02f80 g772869 ( .a(n_7948), .b(n_7833), .o(n_7985) );
na02f80 g778404 ( .a(n_2502), .b(n_2436), .o(n_2537) );
no02f80 g761135 ( .a(n_19106), .b(n_18707), .o(n_19175) );
na02f80 g756719 ( .a(n_23540), .b(n_22354), .o(n_23626) );
in01f80 g761530 ( .a(n_18868), .o(n_18869) );
no02f80 g752809 ( .a(n_28198), .b(n_28078), .o(n_28728) );
no02f80 g761939 ( .a(n_18300), .b(n_18286), .o(n_18343) );
no02f80 g748634 ( .a(n_31304), .b(FE_OCP_DRV_N3160_n_31303), .o(n_31332) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_18_ ( .ck(newNet_2397), .d(n_36442), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_) );
oa22f80 FE_RC_3043_0 ( .a(FE_OFN803_n_46285), .b(n_12158), .c(FE_OFN771_n_46337), .d(n_12133), .o(n_46348) );
in01f80 newInst_1042 ( .a(newNet_1041), .o(newNet_1042) );
in01f80 FE_RC_152_0 ( .a(n_17889), .o(FE_RN_46_0) );
oa12f80 g749670 ( .a(n_30153), .b(n_30152), .c(n_30151), .o(n_30224) );
na02f80 g742737 ( .a(n_37290), .b(n_37068), .o(n_37300) );
no02f80 g774497 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .o(n_6816) );
na02f80 g740078 ( .a(n_39904), .b(n_39802), .o(n_39919) );
na02f80 g784766 ( .a(n_44881), .b(n_37623), .o(n_47252) );
no02f80 g770872 ( .a(n_9937), .b(n_9967), .o(n_10146) );
no02f80 g769367 ( .a(FE_OCPN858_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_23_), .o(n_12083) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_2_ ( .ck(newNet_2921), .d(n_4623), .o(delay_add_ln22_unr5_stage3_stallmux_q_2_) );
na02f80 g779319 ( .a(n_1654), .b(n_1694), .o(n_1762) );
in01f80 FE_OCP_RBC2269_n_33803 ( .a(FE_OCP_RBN3439_n_33803), .o(FE_OCP_RBN2269_n_33803) );
na02f80 g742562 ( .a(n_37532), .b(n_37351), .o(n_37593) );
ao12f80 g779289 ( .a(n_1713), .b(n_1712), .c(n_1711), .o(n_1766) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_18_ ( .ck(newNet_2864), .d(n_11411), .o(delay_add_ln22_unr8_stage4_stallmux_q_18_) );
in01f80 g743289 ( .a(n_36769), .o(n_36770) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_10_ ( .ck(newNet_3456), .d(n_27090), .o(delay_add_ln22_unr17_stage7_stallmux_q_10_) );
ao22s80 g784417 ( .a(n_36355), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n_46229) );
oa12f80 g747308 ( .a(n_32689), .b(n_32688), .c(n_44962), .o(n_32716) );
in01f80 g757790 ( .a(n_22543), .o(n_22513) );
na02f80 g751873 ( .a(n_28148), .b(n_28187), .o(n_28311) );
no02f80 g751544 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_14_), .o(n_28505) );
ao12f80 g744562 ( .a(n_35363), .b(n_35330), .c(n_35328), .o(n_35414) );
oa12f80 g741873 ( .a(n_38408), .b(n_38407), .c(n_38406), .o(n_38483) );
oa12f80 g751287 ( .a(n_28465), .b(n_28747), .c(FE_OCPN1009_n_28439), .o(n_28790) );
in01f80 g754175 ( .a(n_26020), .o(n_26019) );
ao12f80 g750169 ( .a(n_30899), .b(n_30898), .c(n_30897), .o(n_31275) );
in01f80 g749408 ( .a(n_30624), .o(n_30644) );
no02f80 g743110 ( .a(n_36933), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .o(n_37089) );
no03m80 FE_RC_3809_0 ( .a(n_22212), .b(n_22213), .c(n_22304), .o(n_22445) );
in01f80 g778552 ( .a(n_2340), .o(n_2320) );
na02f80 g738821 ( .a(n_41312), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41353) );
na02f80 g768075 ( .a(FE_OCP_RBN3414_n_12739), .b(n_12221), .o(n_12832) );
na02f80 g764108 ( .a(n_16555), .b(n_16558), .o(n_16606) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_21_ ( .ck(newNet_2386), .d(n_36433), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_) );
no02f80 g766009 ( .a(n_14616), .b(n_14551), .o(n_14617) );
no02f80 g778026 ( .a(n_2991), .b(n_2634), .o(n_3022) );
ao12f80 g777706 ( .a(FE_OCP_RBN2463_n_3076), .b(n_3345), .c(n_3059), .o(n_3346) );
no02f80 g768968 ( .a(FE_OCP_RBN2119_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .o(n_12043) );
in01f80 newInst_2699 ( .a(newNet_2698), .o(newNet_2699) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_29_ ( .ck(newNet_2366), .d(n_36592), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_) );
no02f80 g780698 ( .a(n_646), .b(n_641), .o(n_642) );
in01f80 g736538 ( .a(n_43654), .o(n_43665) );
oa22f80 g770257 ( .a(n_10740), .b(n_10554), .c(n_10681), .d(n_10555), .o(n_10848) );
no02f80 g754032 ( .a(n_26369), .b(FE_OCPN1500_n_26125), .o(n_26126) );
in01f80 newInst_3625 ( .a(newNet_3624), .o(newNet_3625) );
oa22f80 g774841 ( .a(n_6259), .b(n_5333), .c(n_6260), .d(n_5334), .o(n_6323) );
ao12f80 g771800 ( .a(n_8714), .b(n_8766), .c(n_8771), .o(n_8872) );
na02f80 g763482 ( .a(FE_OCP_RBN3079_n_16977), .b(FE_OCP_RBN2867_n_16088), .o(n_17119) );
na02f80 g755125 ( .a(n_25374), .b(n_24395), .o(n_25444) );
in01f80 g746902 ( .a(n_33061), .o(n_33036) );
in01f80 g759660 ( .a(n_20510), .o(n_20509) );
na02f80 g777075 ( .a(n_3806), .b(n_3788), .o(n_3957) );
na02f80 g771762 ( .a(n_8980), .b(FE_OCP_RBN3552_n_44575), .o(n_9053) );
no02f80 g746119 ( .a(n_33825), .b(n_34037), .o(n_33854) );
na02f80 g770134 ( .a(n_45304), .b(FE_OCP_RBN3643_n_44490), .o(n_10807) );
no02f80 g754528 ( .a(n_25430), .b(n_25466), .o(n_27009) );
no02f80 g773246 ( .a(n_7582), .b(n_8840), .o(n_7605) );
in01f80 FE_RC_3580_0 ( .a(n_14466), .o(FE_RN_1559_0) );
oa12f80 g765956 ( .a(n_14734), .b(n_14915), .c(n_14735), .o(n_15092) );
na02f80 g746947 ( .a(n_32857), .b(n_32348), .o(n_32942) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_5_ ( .ck(newNet_3482), .d(n_21486), .o(delay_add_ln22_unr14_stage6_stallmux_q_5_) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_2_ ( .ck(newNet_704), .d(n_46141), .o(delay_xor_ln21_unr6_stage3_stallmux_q_2_) );
no02f80 g768381 ( .a(n_12525), .b(n_12505), .o(n_12584) );
oa12f80 g757972 ( .a(n_21925), .b(n_21974), .c(n_21906), .o(n_22049) );
in01f80 g757863 ( .a(n_22279), .o(n_22318) );
na02f80 g761503 ( .a(n_18997), .b(n_19023), .o(n_19128) );
in01f80 newInst_1659 ( .a(newNet_1658), .o(newNet_1659) );
in01f80 g757273 ( .a(n_23107), .o(n_23108) );
in01f80 g755000 ( .a(n_25481), .o(n_25542) );
no02f80 g736568 ( .a(n_43450), .b(n_43449), .o(n_43532) );
in01f80 newInst_116 ( .a(newNet_115), .o(newNet_116) );
no02f80 FE_RC_1827_0 ( .a(FE_OCP_RBN3283_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(FE_RN_547_0) );
na02f80 g773584 ( .a(n_7456), .b(n_7092), .o(n_7454) );
in01f80 FE_RC_3242_0 ( .a(FE_RN_1433_0), .o(FE_RN_1434_0) );
oa22f80 FE_RC_3466_0 ( .a(n_22907), .b(n_22829), .c(n_22580), .d(n_22800), .o(n_22908) );
in01f80 g755384 ( .a(n_25683), .o(n_25575) );
in01f80 g775541 ( .a(n_5375), .o(n_5486) );
no02f80 g751359 ( .a(n_28788), .b(n_28743), .o(n_28789) );
na02f80 g760620 ( .a(n_19878), .b(n_19877), .o(n_19879) );
in01f80 newInst_1748 ( .a(newNet_1747), .o(newNet_1748) );
in01f80 g766335 ( .a(n_14329), .o(n_14366) );
in01f80 g736849 ( .a(n_43547), .o(n_43548) );
in01f80 g745606 ( .a(n_34816), .o(n_34817) );
no02f80 g754224 ( .a(n_26009), .b(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .o(n_26075) );
in01f80 g754927 ( .a(n_25648), .o(n_25649) );
no02f80 g741809 ( .a(n_38321), .b(n_38121), .o(n_38400) );
in01f80 FE_RC_4172_0 ( .a(n_33326), .o(FE_RN_1819_0) );
in01f80 g737762 ( .a(n_42677), .o(n_42678) );
na02f80 g776862 ( .a(n_3969), .b(n_3498), .o(n_4263) );
na02f80 g740003 ( .a(n_40137), .b(n_40188), .o(n_40191) );
in01f80 g774425 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_2_), .o(n_6551) );
in01f80 g771344 ( .a(n_9410), .o(n_9448) );
na02f80 g778942 ( .a(n_2158), .b(n_2156), .o(n_2157) );
in01f80 newInst_3703 ( .a(newNet_1821), .o(newNet_3703) );
na02f80 g759636 ( .a(n_20639), .b(n_45010), .o(n_20726) );
no02f80 g778658 ( .a(n_2380), .b(n_2379), .o(n_3319) );
na02f80 g773523 ( .a(n_7422), .b(n_7290), .o(n_7426) );
in01f80 FE_OCPC1854_n_13366 ( .a(FE_OCPN1853_n_13366), .o(FE_OCPN1854_n_13366) );
in01f80 newInst_2456 ( .a(newNet_2455), .o(newNet_2456) );
in01f80 g779579 ( .a(n_1434), .o(n_1402) );
ao12f80 g773544 ( .a(n_7443), .b(n_7442), .c(n_7441), .o(n_7496) );
in01f80 g754429 ( .a(n_25729), .o(n_25755) );
na02f80 g750510 ( .a(n_29505), .b(FE_OCPN1432_n_29504), .o(n_29570) );
na02f80 g775546 ( .a(n_5632), .b(FE_OCP_RBN2746_n_47011), .o(n_5823) );
oa12f80 g765986 ( .a(n_14636), .b(n_14584), .c(n_14451), .o(n_14696) );
in01f80 FE_OCP_RBC3413_n_12739 ( .a(n_12739), .o(FE_OCP_RBN3413_n_12739) );
ao12f80 g756758 ( .a(n_24172), .b(n_24171), .c(n_24170), .o(n_25092) );
no02f80 g749465 ( .a(n_30531), .b(n_30172), .o(n_30599) );
oa22f80 g776397 ( .a(n_4294), .b(n_4182), .c(FE_OCP_RBN2789_n_4294), .d(n_4046), .o(n_4552) );
in01f80 g773432 ( .a(n_7540), .o(n_7541) );
in01f80 FE_OCPC879_n_31944 ( .a(FE_OCP_RBN3735_n_31819), .o(FE_OCPN879_n_31944) );
na02f80 g742380 ( .a(n_37772), .b(n_37781), .o(n_37837) );
na02f80 g777780 ( .a(n_3232), .b(n_3130), .o(n_3233) );
in01f80 g763164 ( .a(n_17816), .o(n_17817) );
no02f80 g749075 ( .a(n_30956), .b(FE_OCP_RBN1196_n_30926), .o(n_30990) );
no02f80 g736990 ( .a(n_43242), .b(n_43388), .o(n_43470) );
na02f80 g746908 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_14_), .o(n_33099) );
no03m80 FE_RC_3795_0 ( .a(n_37125), .b(n_37272), .c(n_37447), .o(n_37512) );
in01f80 newInst_870 ( .a(newNet_869), .o(newNet_870) );
oa12f80 g772874 ( .a(n_8005), .b(n_8004), .c(n_8003), .o(n_9525) );
in01f80 newInst_2883 ( .a(newNet_2882), .o(newNet_2883) );
in01f80 g739250 ( .a(n_40883), .o(n_40884) );
in01f80 g772015 ( .a(n_9874), .o(n_9824) );
na02f80 g745650 ( .a(n_34101), .b(n_34121), .o(n_34102) );
na02f80 g758040 ( .a(n_22876), .b(n_22878), .o(n_22953) );
na02f80 g765339 ( .a(FE_OCP_RBN2708_n_15135), .b(n_14225), .o(n_15517) );
na02f80 g759224 ( .a(n_21072), .b(n_45032), .o(n_21188) );
na02f80 g741128 ( .a(n_38990), .b(n_38959), .o(n_39046) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_23_ ( .ck(newNet_2646), .d(n_22778), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_) );
ao12f80 g739394 ( .a(n_40774), .b(FE_OCPN897_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_19_), .o(n_41266) );
in01f80 g780099 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .o(n_1131) );
no02f80 g739321 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_24_), .o(n_40862) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_4_ ( .ck(newNet_2711), .d(n_15488), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_) );
na02f80 g746471 ( .a(n_34940), .b(n_44262), .o(n_34941) );
no02f80 g769769 ( .a(n_11193), .b(n_11194), .o(n_11263) );
in01f80 FE_OCP_RBC3839_n_19513 ( .a(FE_OCP_RBN3838_n_19513), .o(FE_OCP_RBN3839_n_19513) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_27_ ( .ck(newNet_2734), .d(n_17697), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_) );
no02f80 g743672 ( .a(n_37436), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_), .o(n_37437) );
no02f80 g773826 ( .a(n_7118), .b(n_7113), .o(n_7114) );
in01f80 g753084 ( .a(n_27305), .o(n_27306) );
na02f80 g745554 ( .a(n_34381), .b(n_34458), .o(n_34533) );
no02f80 g762613 ( .a(n_18022), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_), .o(n_18045) );
in01f80 FE_OCPC994_n_15552 ( .a(FE_OCPN993_n_15552), .o(FE_OCPN994_n_15552) );
no02f80 g751058 ( .a(n_29886), .b(n_29878), .o(n_30358) );
na02f80 g765894 ( .a(n_14999), .b(n_14998), .o(n_15000) );
no02f80 g746417 ( .a(n_33484), .b(n_33482), .o(n_33483) );
no02f80 FE_RC_1333_0 ( .a(FE_RN_395_0), .b(n_39812), .o(n_39907) );
ao22s80 FE_RC_3793_0 ( .a(n_37065), .b(n_37492), .c(n_37066), .d(n_46952), .o(n_37577) );
na02f80 g778047 ( .a(n_2944), .b(n_2263), .o(n_3031) );
in01f80 g766091 ( .a(FE_OCPN971_n_14716), .o(n_14707) );
no02f80 g763596 ( .a(n_17375), .b(n_17156), .o(n_17577) );
no02f80 g780728 ( .a(n_609), .b(n_477), .o(n_616) );
ao12f80 g760044 ( .a(n_20068), .b(n_20897), .c(n_21019), .o(n_21053) );
oa12f80 g765814 ( .a(n_14970), .b(n_14969), .c(n_15032), .o(n_15091) );
na02f80 g746009 ( .a(n_33908), .b(n_33907), .o(n_33963) );
in01f80 g780481 ( .a(n_1148), .o(n_770) );
no02f80 g736793 ( .a(n_43383), .b(n_43388), .o(n_43392) );
ao12f80 g779354 ( .a(n_1629), .b(n_1628), .c(n_1613), .o(n_1787) );
no02f80 g754704 ( .a(n_26231), .b(n_26230), .o(n_26271) );
in01f80 FE_OFC803_n_46285 ( .a(FE_OFN798_n_46285), .o(FE_OFN803_n_46285) );
in01f80 newInst_2293 ( .a(newNet_2292), .o(newNet_2293) );
oa22f80 g752697 ( .a(n_27240), .b(n_27071), .c(n_27239), .d(n_27072), .o(n_27365) );
in01f80 newInst_2192 ( .a(newNet_1299), .o(newNet_2192) );
no02f80 FE_RC_2843_0 ( .a(FE_RN_1221_0), .b(FE_RN_1222_0), .o(FE_RN_1223_0) );
na02f80 g771626 ( .a(n_9332), .b(n_9331), .o(n_9781) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_25_ ( .ck(newNet_2640), .d(n_22806), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_) );
na02f80 g767641 ( .a(n_13019), .b(n_12815), .o(n_13100) );
no02f80 g765010 ( .a(n_15465), .b(n_15420), .o(n_15535) );
in01f80 g758694 ( .a(n_22397), .o(n_22430) );
no02f80 g744797 ( .a(n_35145), .b(n_30545), .o(n_35204) );
in01f80 g756160 ( .a(n_25258), .o(n_24901) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_3_ ( .ck(newNet_2815), .d(n_10000), .o(delay_add_ln22_unr8_stage4_stallmux_q_3_) );
in01f80 g760092 ( .a(n_20534), .o(n_20535) );
in01f80 g742310 ( .a(n_37833), .o(n_37834) );
in01f80 newInst_170 ( .a(newNet_73), .o(newNet_170) );
no02f80 g757489 ( .a(n_22748), .b(n_22927), .o(n_22958) );
in01f80 FE_OCPC3749_n_34296 ( .a(FE_OCPN3748_n_34296), .o(FE_OCPN3749_n_34296) );
na02f80 g779204 ( .a(n_1837), .b(delay_add_ln22_unr2_stage2_stallmux_q_9_), .o(n_1890) );
in01f80 g767415 ( .a(n_13383), .o(n_13384) );
na02f80 g744024 ( .a(n_44223), .b(n_35598), .o(n_36306) );
in01f80 FE_OCPC1452_n_27518 ( .a(FE_OCPN1451_n_27518), .o(FE_OCPN1452_n_27518) );
no02f80 g770035 ( .a(n_10833), .b(n_44498), .o(n_10859) );
no02f80 g771976 ( .a(n_44498), .b(n_9994), .o(n_10037) );
in01f80 g766039 ( .a(n_14673), .o(n_14714) );
in01f80 g736881 ( .a(n_43599), .o(n_43600) );
in01f80 g751441 ( .a(n_28526), .o(n_28527) );
oa12f80 g756445 ( .a(n_23783), .b(n_23922), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n_23927) );
no03m80 g762178 ( .a(n_18737), .b(n_18625), .c(n_18765), .o(n_18738) );
in01f80 newInst_2167 ( .a(newNet_2166), .o(newNet_2167) );
na02f80 g769734 ( .a(n_11169), .b(n_11141), .o(n_11202) );
in01f80 g738567 ( .a(n_41618), .o(n_41619) );
no02f80 g760212 ( .a(FE_OCP_RBN1332_n_20249), .b(FE_OCPN1044_n_20307), .o(n_20332) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_19_ ( .ck(newNet_2479), .d(n_32281), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_) );
oa12f80 g763124 ( .a(n_17398), .b(n_17481), .c(n_17279), .o(n_17588) );
no02f80 g740205 ( .a(n_39812), .b(n_39536), .o(n_40016) );
in01f80 g780703 ( .a(n_893), .o(n_640) );
na02f80 g763589 ( .a(n_16807), .b(n_44365), .o(n_16899) );
na02f80 g764294 ( .a(n_16330), .b(n_14588), .o(n_16441) );
oa12f80 g775466 ( .a(n_5666), .b(n_5716), .c(n_5665), .o(n_5753) );
na02f80 g738497 ( .a(n_41540), .b(n_41298), .o(n_41669) );
in01f80 newInst_3197 ( .a(newNet_3196), .o(newNet_3197) );
na02f80 g746998 ( .a(n_32822), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_), .o(n_32878) );
in01f80 g777399 ( .a(n_3570), .o(n_3571) );
na02f80 g738240 ( .a(n_41896), .b(n_41753), .o(n_41946) );
no02f80 g745762 ( .a(n_34183), .b(n_34182), .o(n_34247) );
in01f80 FE_OCP_RBC2483_n_14326 ( .a(n_14326), .o(FE_OCP_RBN2483_n_14326) );
in01f80 newInst_2390 ( .a(newNet_1486), .o(newNet_2390) );
na02f80 g753640 ( .a(n_26594), .b(n_26599), .o(n_26595) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_13_ ( .ck(newNet_1540), .d(n_32065), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_) );
na02f80 g739000 ( .a(n_41158), .b(n_40936), .o(n_41186) );
na02f80 g748526 ( .a(n_31677), .b(n_31676), .o(n_31756) );
na02f80 g737619 ( .a(n_42223), .b(n_42208), .o(n_42224) );
no02f80 g736952 ( .a(n_43038), .b(n_42924), .o(n_43270) );
in01f80 g738290 ( .a(n_41776), .o(n_41777) );
in01f80 g780204 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_5_), .o(n_1039) );
ao12f80 g773841 ( .a(n_7087), .b(n_7084), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .o(n_7180) );
in01f80 g755486 ( .a(n_24754), .o(n_24752) );
no02f80 g771843 ( .a(FE_OCPN1388_n_11041), .b(n_10081), .o(n_10156) );
in01f80 newInst_394 ( .a(newNet_393), .o(newNet_394) );
na02f80 g772628 ( .a(n_8252), .b(n_8170), .o(n_8352) );
in01f80 FE_OCP_DRV_C1588_n_31012 ( .a(FE_OCP_DRV_N1587_n_31012), .o(FE_OCP_DRV_N1588_n_31012) );
in01f80 g773954 ( .a(n_7289), .o(n_7290) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_8_ ( .ck(newNet_2990), .d(n_1019), .o(delay_add_ln22_unr2_stage2_stallmux_q_8_) );
oa12f80 g747138 ( .a(n_32887), .b(n_32886), .c(n_32885), .o(n_33756) );
in01f80 FE_RC_3301_0 ( .a(n_17971), .o(FE_RN_1453_0) );
in01f80 g774442 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .o(n_6542) );
in01f80 g765976 ( .a(n_14845), .o(n_14788) );
in01f80 g751369 ( .a(n_29036), .o(n_28771) );
in01f80 newInst_164 ( .a(newNet_163), .o(newNet_164) );
na02f80 g749756 ( .a(n_29905), .b(n_29814), .o(n_29903) );
ao12f80 g738879 ( .a(n_41015), .b(n_41196), .c(n_40886), .o(n_41288) );
in01f80 g745755 ( .a(n_34362), .o(n_34363) );
in01f80 g737178 ( .a(n_46935), .o(n_43010) );
no02f80 g750045 ( .a(n_29869), .b(n_28892), .o(n_29897) );
in01f80 g756787 ( .a(n_23938), .o(n_23991) );
no02f80 g759001 ( .a(n_21571), .b(n_45080), .o(n_21605) );
in01f80 g774234 ( .a(n_6609), .o(n_6610) );
na02f80 g764823 ( .a(n_15623), .b(n_15591), .o(n_15702) );
ms00f80 mux_while_ln12_psv_q_reg_8_ ( .ck(newNet_98), .d(n_265), .o(mux_while_ln12_psv_q_8_) );
ao12f80 g754419 ( .a(n_26386), .b(n_26231), .c(n_26420), .o(n_26941) );
no02f80 g764866 ( .a(n_15557), .b(n_14452), .o(n_15627) );
in01f80 g747850 ( .a(n_32236), .o(n_32237) );
no02f80 g736733 ( .a(n_43362), .b(n_43361), .o(n_43363) );
na02f80 g766190 ( .a(n_14379), .b(n_14378), .o(n_14475) );
no02f80 g758041 ( .a(n_22647), .b(n_22697), .o(n_22698) );
in01f80 FE_OCP_RBC1707_n_20616 ( .a(n_20616), .o(FE_OCP_RBN1707_n_20616) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_7_ ( .ck(newNet_611), .d(n_46378), .o(delay_xor_ln21_unr9_stage4_stallmux_q_7_) );
na02f80 g784137 ( .a(n_7136), .b(n_7135), .o(n_45884) );
na02f80 g779768 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .o(n_1507) );
in01f80 g767318 ( .a(n_13697), .o(n_13716) );
in01f80 g762026 ( .a(n_18458), .o(n_18459) );
na02f80 g738068 ( .a(n_42074), .b(n_42060), .o(n_42137) );
no02f80 g738857 ( .a(n_41285), .b(n_41337), .o(n_41311) );
na02f80 g770279 ( .a(n_10573), .b(n_10592), .o(n_10618) );
in01f80 g751236 ( .a(n_30097), .o(n_30156) );
no02f80 g756730 ( .a(n_23501), .b(n_23465), .o(n_23576) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_28_ ( .ck(newNet_1296), .d(n_1275), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_) );
no02f80 FE_RC_2295_0 ( .a(FE_RN_863_0), .b(n_28200), .o(FE_RN_864_0) );
na02f80 g754098 ( .a(n_26146), .b(n_23467), .o(n_26147) );
na02f80 g767420 ( .a(n_13268), .b(n_13332), .o(n_13361) );
na02f80 g767942 ( .a(n_12694), .b(n_12693), .o(n_12773) );
in01f80 newInst_2463 ( .a(newNet_2462), .o(newNet_2463) );
na02f80 g738433 ( .a(n_41573), .b(n_41672), .o(n_41733) );
na02f80 g781251 ( .a(n_79), .b(n_146), .o(n_165) );
na02f80 g754083 ( .a(n_26068), .b(FE_OCP_RBN2836_FE_RN_745_0), .o(n_26129) );
in01f80 g778097 ( .a(n_3016), .o(n_3041) );
no02f80 g753133 ( .a(n_27392), .b(n_27346), .o(n_27498) );
no02f80 g784755 ( .a(n_47235), .b(n_7730), .o(n_47241) );
no02f80 g777727 ( .a(n_3435), .b(n_3434), .o(n_3436) );
in01f80 g758922 ( .a(n_21330), .o(n_21331) );
no02f80 g776910 ( .a(n_3761), .b(n_3082), .o(n_3851) );
in01f80 newInst_3632 ( .a(newNet_2310), .o(newNet_3632) );
no02f80 g738410 ( .a(n_41743), .b(n_41769), .o(n_41820) );
oa12f80 g749968 ( .a(n_29959), .b(n_29896), .c(FE_OCP_RBN1325_n_29056), .o(n_30488) );
in01f80 g744378 ( .a(n_46212), .o(n_36808) );
no02f80 g762339 ( .a(n_45002), .b(n_18441), .o(n_18834) );
oa22f80 FE_RC_2533_0 ( .a(FE_RN_1032_0), .b(n_17315), .c(FE_OCP_RBN3098_n_17315), .d(n_17510), .o(n_17687) );
na02f80 g748751 ( .a(n_31232), .b(n_31099), .o(n_31266) );
na02f80 g749300 ( .a(n_30625), .b(FE_OCPN1410_n_27014), .o(n_30743) );
in01f80 g741507 ( .a(n_38743), .o(n_38748) );
in01f80 g770042 ( .a(n_11063), .o(n_11064) );
in01f80 g754352 ( .a(n_25890), .o(n_25891) );
in01f80 g762747 ( .a(n_18036), .o(n_18037) );
oa12f80 g756879 ( .a(n_23906), .b(n_24188), .c(n_23863), .o(n_24769) );
in01f80 FE_RC_3019_0 ( .a(n_46426), .o(FE_RN_1324_0) );
ao12f80 g749615 ( .a(n_30459), .b(n_30458), .c(n_30457), .o(n_31504) );
no02f80 g767971 ( .a(FE_OCPN860_n_12880), .b(n_13163), .o(n_13198) );
no02f80 g751539 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_22_), .o(n_28605) );
na02f80 g765354 ( .a(n_15330), .b(n_15373), .o(n_15404) );
in01f80 FE_OCP_RBC2640_n_34921 ( .a(n_34921), .o(FE_OCP_RBN2640_n_34921) );
ao22s80 g772042 ( .a(FE_OCP_RBN2477_n_8599), .b(n_8831), .c(n_8832), .d(n_8599), .o(n_9004) );
no03m80 g752166 ( .a(n_28615), .b(n_28591), .c(n_28105), .o(n_28714) );
na02f80 g750410 ( .a(n_29642), .b(n_29656), .o(n_29739) );
in01f80 g775438 ( .a(n_5796), .o(n_5797) );
no02f80 g776356 ( .a(n_4634), .b(n_4222), .o(n_4680) );
no02f80 g773379 ( .a(n_7528), .b(n_7070), .o(n_7612) );
in01f80 g764763 ( .a(n_15704), .o(n_15772) );
in01f80 FE_OCP_RBC2845_n_10326 ( .a(FE_OCP_RBN2844_n_10326), .o(FE_OCP_RBN2845_n_10326) );
no02f80 g750890 ( .a(n_29080), .b(n_29109), .o(n_29157) );
in01f80 g775473 ( .a(n_5756), .o(n_5757) );
in01f80 FE_OCP_RBC1840_n_19528 ( .a(n_19528), .o(FE_OCP_RBN1840_n_19528) );
no02f80 g768580 ( .a(n_12296), .b(n_12295), .o(n_12297) );
oa22f80 FE_RC_778_0 ( .a(n_8667), .b(n_8388), .c(n_8750), .d(n_8666), .o(n_8782) );
in01f80 g744389 ( .a(n_36793), .o(n_36794) );
no02f80 g741813 ( .a(n_38444), .b(n_38443), .o(n_38445) );
in01f80 FE_OCP_RBC2435_n_14072 ( .a(FE_OCP_RBN2434_n_14072), .o(FE_OCP_RBN2435_n_14072) );
in01f80 g758334 ( .a(n_22466), .o(n_22432) );
in01f80 newInst_2781 ( .a(newNet_122), .o(newNet_2781) );
in01f80 g746383 ( .a(n_33558), .o(n_33610) );
oa22f80 g747773 ( .a(n_33372), .b(n_33576), .c(n_33571), .d(n_33415), .o(n_33862) );
no02f80 g745823 ( .a(n_44102), .b(n_33708), .o(n_34618) );
in01f80 g759898 ( .a(n_21598), .o(n_21561) );
no02f80 g759963 ( .a(n_21051), .b(n_20199), .o(n_21295) );
in01f80 FE_OCP_RBC2742_n_15206 ( .a(n_15206), .o(FE_OCP_RBN2742_n_15206) );
na02f80 g767374 ( .a(n_13406), .b(n_13334), .o(n_13389) );
in01f80 g749054 ( .a(n_32272), .o(n_32273) );
in01f80 g742387 ( .a(n_37778), .o(n_37809) );
ao22s80 FE_RC_543_0 ( .a(n_44441), .b(n_25785), .c(n_25507), .d(n_25818), .o(n_25915) );
in01f80 g743328 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .o(n_36708) );
na02f80 g759705 ( .a(n_21255), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21256) );
no02f80 g752139 ( .a(n_28116), .b(n_28115), .o(n_28139) );
in01f80 g750266 ( .a(n_31213), .o(n_30968) );
in01f80 newInst_2800 ( .a(newNet_2799), .o(newNet_2800) );
in01f80 g784391 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46197) );
in01f80 g767231 ( .a(n_13765), .o(n_13760) );
no02f80 g744053 ( .a(n_44222), .b(n_34752), .o(n_35826) );
no02f80 g748405 ( .a(FE_OCPN1052_n_31674), .b(n_30757), .o(n_31762) );
in01f80 newInst_1013 ( .a(newNet_1012), .o(newNet_1013) );
in01f80 g778141 ( .a(n_2964), .o(n_2965) );
in01f80 g746230 ( .a(n_35629), .o(n_35125) );
in01f80 g744461 ( .a(n_35484), .o(n_35485) );
na02f80 g780131 ( .a(n_1160), .b(n_1159), .o(n_1161) );
na02f80 g773385 ( .a(n_7581), .b(n_7567), .o(n_7609) );
na02f80 g762250 ( .a(n_18608), .b(n_18657), .o(n_18696) );
no02f80 g750072 ( .a(n_29869), .b(n_30111), .o(n_30173) );
in01f80 g780041 ( .a(n_1248), .o(n_1250) );
in01f80 newInst_3090 ( .a(newNet_3089), .o(newNet_3090) );
na02f80 g759925 ( .a(n_21051), .b(n_21246), .o(n_21826) );
in01f80 FE_RC_3701_0 ( .a(n_3492), .o(FE_RN_1629_0) );
no02f80 g739061 ( .a(n_41110), .b(n_40959), .o(n_41138) );
na02f80 g778602 ( .a(FE_OCP_RBN2296_n_2438), .b(n_2744), .o(n_2720) );
in01f80 newInst_2500 ( .a(newNet_2499), .o(newNet_2500) );
na02f80 g754265 ( .a(n_25874), .b(FE_OCPN1514_FE_OFN738_n_22641), .o(n_25919) );
in01f80 g738674 ( .a(n_41607), .o(n_41721) );
in01f80 g764712 ( .a(n_15861), .o(n_15862) );
ao22s80 FE_RC_865_0 ( .a(n_24745), .b(FE_OCPN1474_n_24624), .c(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .d(n_24718), .o(n_24875) );
in01f80 newInst_2976 ( .a(newNet_692), .o(newNet_2976) );
in01f80 g771432 ( .a(n_9089), .o(n_9149) );
in01f80 g763912 ( .a(n_17354), .o(n_17299) );
na02f80 g745564 ( .a(n_34648), .b(n_34674), .o(n_34745) );
no02f80 g758053 ( .a(n_22653), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n_22731) );
na02f80 g744399 ( .a(n_35493), .b(n_35503), .o(n_35494) );
no02f80 g771674 ( .a(n_9066), .b(n_44516), .o(n_10340) );
no02f80 g759200 ( .a(n_21271), .b(n_46967), .o(n_21459) );
in01f80 g737708 ( .a(n_42419), .o(n_42464) );
in01f80 g754447 ( .a(n_25676), .o(n_25677) );
na02f80 g739957 ( .a(n_40085), .b(n_40021), .o(n_40161) );
in01f80 g774026 ( .a(n_6918), .o(n_6919) );
na02f80 g759464 ( .a(n_20907), .b(FE_RN_1585_0), .o(n_20967) );
ao12f80 g742666 ( .a(n_37487), .b(n_37486), .c(n_37485), .o(n_37547) );
in01f80 FE_OCP_RBC3824_n_44061 ( .a(n_44061), .o(FE_OCP_RBN3824_n_44061) );
in01f80 g767562 ( .a(n_12904), .o(n_12945) );
no02f80 g761763 ( .a(n_18564), .b(n_18437), .o(n_18565) );
na02f80 g769833 ( .a(n_11025), .b(n_11062), .o(n_11137) );
na02f80 FE_RC_80_0 ( .a(FE_RN_21_0), .b(FE_RN_22_0), .o(FE_RN_23_0) );
in01f80 newInst_2486 ( .a(newNet_2485), .o(newNet_2486) );
na02f80 g770890 ( .a(n_9992), .b(FE_OFN755_n_44461), .o(n_10107) );
no02f80 g776882 ( .a(n_3739), .b(n_3785), .o(n_3933) );
no02f80 g767699 ( .a(n_13208), .b(n_13197), .o(n_13171) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_27_ ( .ck(newNet_314), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_27_) );
in01f80 newInst_1165 ( .a(newNet_1164), .o(newNet_1165) );
in01f80 g771825 ( .a(n_9955), .o(n_9830) );
oa12f80 g746391 ( .a(n_35021), .b(n_35020), .c(n_35019), .o(n_35633) );
in01f80 g770974 ( .a(n_9856), .o(n_9857) );
in01f80 newInst_724 ( .a(newNet_723), .o(newNet_724) );
na02f80 g746804 ( .a(n_33325), .b(n_33339), .o(n_33404) );
in01f80 newInst_152 ( .a(newNet_151), .o(newNet_152) );
na02f80 g770075 ( .a(n_10950), .b(FE_OCP_RBN2661_n_9292), .o(n_11106) );
no02f80 g756305 ( .a(n_24588), .b(n_24062), .o(n_24606) );
no02f80 FE_RC_3302_0 ( .a(FE_RN_1451_0), .b(FE_RN_1453_0), .o(FE_RN_1454_0) );
in01f80 newInst_1081 ( .a(newNet_1080), .o(newNet_1081) );
ao12f80 g759740 ( .a(n_21374), .b(n_21825), .c(n_21719), .o(n_21781) );
in01f80 g757195 ( .a(n_23195), .o(n_23212) );
in01f80 newInst_539 ( .a(newNet_538), .o(newNet_539) );
oa12f80 g768323 ( .a(n_12510), .b(n_12509), .c(n_12508), .o(n_13590) );
in01f80 g740561 ( .a(n_39722), .o(n_39723) );
oa22f80 FE_RC_1388_0 ( .a(FE_OFN802_n_46285), .b(n_12150), .c(n_12058), .d(FE_OFN771_n_46337), .o(n_46356) );
ao22s80 FE_RC_806_0 ( .a(n_9011), .b(n_7589), .c(n_7588), .d(n_9010), .o(n_9188) );
no02f80 g770313 ( .a(n_10480), .b(FE_OCP_RBN3637_n_44490), .o(n_10488) );
in01f80 g774474 ( .a(n_6857), .o(n_6773) );
na02f80 g763065 ( .a(n_17862), .b(n_17499), .o(n_17937) );
in01f80 FE_OCP_RBC2933_n_31010 ( .a(n_31010), .o(FE_OCP_RBN2933_n_31010) );
na02f80 g768254 ( .a(n_12604), .b(n_12157), .o(n_12662) );
in01f80 g765984 ( .a(n_14722), .o(n_14723) );
in01f80 g742168 ( .a(n_38211), .o(n_38212) );
na02f80 g738507 ( .a(FE_OCP_RBN2313_n_41420), .b(n_41317), .o(n_41635) );
in01f80 g770633 ( .a(n_10377), .o(n_10474) );
no02f80 g755394 ( .a(n_24872), .b(n_22393), .o(n_24873) );
ao12f80 g747305 ( .a(n_32554), .b(FE_OCP_RBN2102_n_44962), .c(delay_xor_ln21_unr21_stage8_stallmux_q_9_), .o(n_32579) );
in01f80 FE_OCP_RBC3683_FE_RN_770_0 ( .a(FE_RN_770_0), .o(FE_OCP_RBN3683_FE_RN_770_0) );
oa22f80 g779884 ( .a(n_44652), .b(n_1144), .c(n_44623), .d(n_1125), .o(n_1351) );
in01f80 newInst_2341 ( .a(newNet_2340), .o(newNet_2341) );
no02f80 g759976 ( .a(n_20336), .b(n_45066), .o(n_20381) );
no02f80 g737321 ( .a(n_42864), .b(n_42488), .o(n_42909) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_21_ ( .ck(newNet_1403), .d(n_36699), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_) );
no02f80 g777138 ( .a(n_3725), .b(n_151), .o(n_3767) );
no02f80 g772319 ( .a(n_8725), .b(n_8724), .o(n_8726) );
oa12f80 g739554 ( .a(n_40634), .b(n_40633), .c(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n_41309) );
no02f80 g736807 ( .a(n_43464), .b(n_43001), .o(n_43346) );
no02f80 g777172 ( .a(n_4371), .b(n_4262), .o(n_5079) );
ao12f80 g748092 ( .a(n_31468), .b(n_31506), .c(n_31519), .o(n_31614) );
in01f80 newInst_373 ( .a(newNet_372), .o(newNet_373) );
in01f80 g740605 ( .a(n_39662), .o(n_39669) );
oa22f80 FE_RC_3247_0 ( .a(n_10446), .b(n_10366), .c(n_10445), .d(n_10365), .o(n_10568) );
in01f80 g748323 ( .a(n_31556), .o(n_31557) );
no02f80 g761961 ( .a(n_18285), .b(n_18263), .o(n_18286) );
in01f80 g737222 ( .a(n_42970), .o(n_42971) );
na02f80 g760193 ( .a(n_20954), .b(n_20051), .o(n_21099) );
ao12f80 g760714 ( .a(n_19692), .b(n_19623), .c(n_19555), .o(n_19877) );
no02f80 g777150 ( .a(n_4773), .b(n_4731), .o(n_4788) );
in01f80 g767880 ( .a(n_46933), .o(n_12823) );
in01f80 FE_OCP_RBC3573_n_44563 ( .a(FE_OCP_RBN3572_n_44563), .o(FE_OCP_RBN3573_n_44563) );
no02f80 g748624 ( .a(n_31422), .b(n_31195), .o(n_31444) );
in01f80 g757485 ( .a(n_22945), .o(n_22900) );
ao12f80 g779064 ( .a(n_1484), .b(n_2023), .c(n_1682), .o(n_2054) );
in01f80 g755180 ( .a(n_25203), .o(n_25204) );
in01f80 g769891 ( .a(n_11132), .o(n_11192) );
no02f80 g760701 ( .a(n_19742), .b(FE_OCP_RBN3842_n_19555), .o(n_19743) );
in01f80 newInst_3656 ( .a(newNet_407), .o(newNet_3656) );
in01f80 newInst_845 ( .a(newNet_844), .o(newNet_845) );
in01f80 g758861 ( .a(n_21579), .o(n_21580) );
no02f80 g750322 ( .a(n_29731), .b(n_29531), .o(n_29808) );
na02f80 g757836 ( .a(n_23085), .b(n_23052), .o(n_23086) );
na02f80 g767433 ( .a(n_13228), .b(n_12910), .o(n_13268) );
na02f80 g759542 ( .a(n_20689), .b(n_20690), .o(n_20732) );
in01f80 g773408 ( .a(n_7567), .o(n_7568) );
na02f80 g779316 ( .a(n_1667), .b(n_1666), .o(n_1768) );
in01f80 g750377 ( .a(n_29648), .o(n_29664) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_7_ ( .ck(newNet_3581), .d(n_15757), .o(delay_add_ln22_unr11_stage5_stallmux_q_7_) );
oa12f80 g760441 ( .a(n_20074), .b(n_20078), .c(n_20073), .o(n_21790) );
in01f80 FE_OFC750_n_45003 ( .a(FE_OFN749_n_45003), .o(FE_OFN750_n_45003) );
in01f80 g765397 ( .a(n_15449), .o(n_15450) );
in01f80 g758884 ( .a(n_21438), .o(n_21439) );
na02f80 FE_RC_1205_0 ( .a(FE_RN_363_0), .b(FE_RN_364_0), .o(FE_RN_365_0) );
na02f80 g754036 ( .a(n_26071), .b(n_25625), .o(n_26153) );
na02f80 g744556 ( .a(n_35365), .b(n_35257), .o(n_35364) );
in01f80 g740455 ( .a(n_39788), .o(n_39789) );
in01f80 FE_OCP_RBC3497_n_13818 ( .a(FE_OCP_RBN3496_n_13818), .o(FE_OCP_RBN3497_n_13818) );
no02f80 g769657 ( .a(n_11257), .b(n_11244), .o(n_11302) );
no02f80 g737673 ( .a(FE_OCPN887_n_42367), .b(n_42710), .o(n_42724) );
no02f80 g747047 ( .a(n_34019), .b(n_33950), .o(n_34075) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_7_ ( .ck(newNet_1898), .d(n_36890), .o(delay_sub_ln22_unr24_stage9_stallmux_q_7_) );
in01f80 g749378 ( .a(n_30609), .o(n_30610) );
in01f80 FE_OCP_RBC3834_n_19241 ( .a(FE_OCP_RBN3833_n_19241), .o(FE_OCP_RBN3834_n_19241) );
in01f80 newInst_317 ( .a(newNet_39), .o(newNet_317) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_11_ ( .ck(newNet_673), .d(n_46365), .o(delay_xor_ln21_unr9_stage4_stallmux_q_11_) );
in01f80 FE_OCPC3782_n_16463 ( .a(n_16463), .o(FE_OCPN3782_n_16463) );
na02f80 g765837 ( .a(n_14972), .b(n_14971), .o(n_14973) );
na02f80 FE_RC_2897_0 ( .a(n_9603), .b(n_9655), .o(FE_RN_1255_0) );
na02f80 g771450 ( .a(FE_OCP_RBN2529_n_9044), .b(n_8992), .o(n_9146) );
in01f80 g767813 ( .a(n_13160), .o(n_13243) );
oa12f80 g751382 ( .a(n_29337), .b(n_29363), .c(n_29336), .o(n_29817) );
na02f80 g737063 ( .a(n_43230), .b(n_42990), .o(n_43424) );
in01f80 g746042 ( .a(n_35258), .o(n_35240) );
in01f80 g776262 ( .a(n_4806), .o(n_4891) );
in01f80 g756205 ( .a(n_24125), .o(n_25228) );
na02f80 FE_RC_81_0 ( .a(FE_RN_23_0), .b(n_17743), .o(n_17841) );
in01f80 g762019 ( .a(n_18506), .o(n_18507) );
oa12f80 g758659 ( .a(n_21803), .b(n_21818), .c(n_21761), .o(n_21898) );
oa12f80 g751617 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .c(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_28742) );
no02f80 g749678 ( .a(n_30079), .b(n_29862), .o(n_30149) );
no02f80 g773782 ( .a(n_7137), .b(n_7119), .o(n_7120) );
in01f80 FE_RC_1503_0 ( .a(n_47258), .o(FE_RN_420_0) );
in01f80 newInst_97 ( .a(newNet_96), .o(newNet_97) );
in01f80 newInst_1883 ( .a(newNet_1882), .o(newNet_1883) );
ao22s80 g750970 ( .a(n_28871), .b(n_28886), .c(n_28967), .d(n_28885), .o(n_30364) );
in01f80 g776468 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_), .o(n_6698) );
na02f80 g743298 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n_36875) );
na02f80 FE_RC_2836_0 ( .a(FE_OCP_RBN2867_n_16088), .b(n_16943), .o(FE_RN_1219_0) );
in01f80 g775384 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .o(n_5884) );
oa22f80 g754450 ( .a(n_25653), .b(n_25427), .c(n_25675), .d(n_25428), .o(n_27416) );
in01f80 FE_OCPC1455_n_18860 ( .a(n_18860), .o(FE_OCPN1455_n_18860) );
no02f80 FE_RC_3897_0 ( .a(FE_RN_1692_0), .b(n_24646), .o(n_24686) );
in01f80 newInst_1230 ( .a(newNet_281), .o(newNet_1230) );
in01f80 g762753 ( .a(n_18183), .o(n_18184) );
in01f80 g759880 ( .a(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_21975) );
in01f80 g770472 ( .a(n_10478), .o(n_10479) );
na02f80 g771616 ( .a(n_9379), .b(n_9378), .o(n_9439) );
in01f80 g743235 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_4_), .o(n_36873) );
no02f80 g767337 ( .a(n_13481), .b(n_13507), .o(n_13547) );
ao12f80 g779196 ( .a(n_1925), .b(n_1924), .c(n_1923), .o(n_1965) );
oa12f80 g771157 ( .a(n_9738), .b(n_9794), .c(n_9737), .o(n_9842) );
in01f80 g763670 ( .a(n_17374), .o(n_17375) );
na02f80 g767536 ( .a(n_13094), .b(n_13063), .o(n_13265) );
na03f80 FE_RC_1053_0 ( .a(n_40878), .b(n_40934), .c(n_40936), .o(n_46947) );
in01f80 g749175 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n_32422) );
in01f80 g747203 ( .a(n_34582), .o(n_33865) );
no02f80 g741572 ( .a(n_38659), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38716) );
in01f80 g759198 ( .a(n_21346), .o(n_21345) );
in01f80 newInst_3489 ( .a(newNet_3488), .o(newNet_3489) );
no02f80 g776131 ( .a(n_4570), .b(n_4523), .o(n_4726) );
no02f80 FE_RC_2714_0 ( .a(n_23122), .b(n_23014), .o(FE_RN_1144_0) );
in01f80 newInst_3746 ( .a(newNet_3141), .o(newNet_3746) );
in01f80 g757450 ( .a(n_23391), .o(n_23031) );
in01f80 g750341 ( .a(n_30719), .o(n_30756) );
na02f80 g740080 ( .a(n_40291), .b(n_40215), .o(n_40328) );
in01f80 g750176 ( .a(n_29888), .o(n_29889) );
in01f80 g758689 ( .a(n_21944), .o(n_21945) );
no02f80 g764963 ( .a(n_15468), .b(n_15385), .o(n_15501) );
na02f80 g773087 ( .a(n_7993), .b(n_8045), .o(n_8086) );
no02f80 g764311 ( .a(n_16398), .b(n_14588), .o(n_16431) );
no02f80 g771936 ( .a(n_8694), .b(n_7601), .o(n_8749) );
ao12f80 g773958 ( .a(n_7257), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .o(n_7404) );
oa12f80 g751699 ( .a(n_28364), .b(n_28363), .c(n_28362), .o(n_29576) );
in01f80 FE_OCP_RBC2317_n_41420 ( .a(FE_OCP_RBN2315_n_41420), .o(FE_OCP_RBN2317_n_41420) );
no02f80 g766373 ( .a(n_14653), .b(n_14137), .o(n_14703) );
in01f80 newInst_1666 ( .a(newNet_1230), .o(newNet_1666) );
na02f80 g740519 ( .a(n_39732), .b(n_39730), .o(n_39778) );
in01f80 newInst_1088 ( .a(newNet_1087), .o(newNet_1088) );
in01f80 newInst_1991 ( .a(newNet_934), .o(newNet_1991) );
no02f80 g746134 ( .a(n_33896), .b(FE_OCP_RBN3439_n_33803), .o(n_33939) );
in01f80 g737180 ( .a(n_43006), .o(n_43418) );
in01f80 g778252 ( .a(n_2829), .o(n_2776) );
no02f80 g743922 ( .a(n_35704), .b(n_44223), .o(n_35872) );
in01f80 newInst_3221 ( .a(newNet_1017), .o(newNet_3221) );
oa12f80 g772677 ( .a(n_7815), .b(n_8131), .c(n_7770), .o(n_8215) );
in01f80 g747796 ( .a(n_33317), .o(n_33296) );
oa12f80 g772345 ( .a(n_8555), .b(n_44058), .c(n_8482), .o(n_8585) );
na02f80 g766138 ( .a(n_14682), .b(n_14655), .o(n_14736) );
in01f80 g759185 ( .a(n_21186), .o(n_21187) );
in01f80 g738223 ( .a(n_41971), .o(n_41972) );
in01f80 g758469 ( .a(n_25824), .o(n_25831) );
no02f80 g748974 ( .a(n_31079), .b(n_30963), .o(n_31132) );
oa22f80 g749115 ( .a(n_32203), .b(n_31625), .c(n_32204), .d(n_31626), .o(n_32256) );
in01f80 g775330 ( .a(n_5816), .o(n_5854) );
in01f80 newInst_2352 ( .a(newNet_439), .o(newNet_2352) );
no02f80 g742641 ( .a(n_37416), .b(n_37152), .o(n_37448) );
in01f80 g738212 ( .a(n_41974), .o(n_41973) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_13_ ( .ck(newNet_3647), .d(n_46979), .o(delay_add_ln22_unr11_stage5_stallmux_q_13_) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_17_ ( .ck(newNet_1416), .d(n_36641), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_) );
na02f80 g757084 ( .a(n_23289), .b(n_23281), .o(n_23303) );
in01f80 g748201 ( .a(n_32122), .o(n_32123) );
oa22f80 g748959 ( .a(n_32273), .b(n_31577), .c(n_32272), .d(n_31576), .o(n_32342) );
na02f80 g780717 ( .a(n_626), .b(n_624), .o(n_625) );
in01f80 newInst_2222 ( .a(newNet_1691), .o(newNet_2222) );
oa12f80 g749692 ( .a(n_29829), .b(n_29970), .c(n_29859), .o(n_30057) );
no02f80 g738114 ( .a(n_42070), .b(n_42054), .o(n_42055) );
no02f80 g769386 ( .a(n_9993), .b(FE_OCP_RBN2105_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11686) );
no02f80 g778119 ( .a(n_2789), .b(n_2226), .o(n_2855) );
ao12f80 g738097 ( .a(n_41772), .b(n_42070), .c(n_41751), .o(n_42085) );
in01f80 g760868 ( .a(n_19511), .o(n_19512) );
na02f80 g768248 ( .a(n_12675), .b(n_12384), .o(n_12698) );
in01f80 g766411 ( .a(n_14271), .o(n_14272) );
na02f80 g751988 ( .a(n_28793), .b(n_28860), .o(n_28904) );
in01f80 g763325 ( .a(n_46973), .o(n_17187) );
no02f80 g742810 ( .a(n_37233), .b(n_37067), .o(n_37232) );
na02f80 g771062 ( .a(n_10001), .b(n_9961), .o(n_9962) );
na02f80 g747097 ( .a(n_32735), .b(n_32799), .o(n_32834) );
na02f80 g736509 ( .a(n_43687), .b(n_43277), .o(n_43714) );
in01f80 newInst_3574 ( .a(newNet_3573), .o(newNet_3574) );
na02f80 g774164 ( .a(n_6769), .b(n_6830), .o(n_7515) );
no02f80 g768964 ( .a(FE_OCP_RBN1138_n_11779), .b(n_11730), .o(n_11819) );
na02f80 FE_RC_2554_0 ( .a(FE_RN_1045_0), .b(FE_RN_1046_0), .o(FE_RN_1047_0) );
in01f80 FE_OCPC3188_n_11012 ( .a(FE_OCPN3187_n_11012), .o(FE_OCPN3188_n_11012) );
no02f80 g771512 ( .a(n_8843), .b(n_8845), .o(n_8951) );
na02f80 g771124 ( .a(n_9594), .b(n_9570), .o(n_9676) );
in01f80 FE_OCPC895_n_6521 ( .a(FE_OCPN894_n_6521), .o(FE_OCPN895_n_6521) );
in01f80 g755842 ( .a(FE_OCPN1500_n_26125), .o(n_26214) );
na02f80 FE_RC_3064_0 ( .a(n_20429), .b(FE_RN_1345_0), .o(FE_RN_1346_0) );
ao12f80 g762798 ( .a(n_17845), .b(FE_OCP_RBN2140_FE_OCPN861_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_12_), .o(n_17868) );
ao12f80 g741346 ( .a(n_38761), .b(n_38801), .c(n_38783), .o(n_38856) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_13_ ( .ck(newNet_366), .d(n_1355), .o(delay_xor_ln22_unr3_stage2_stallmux_q_13_) );
in01f80 g767402 ( .a(n_13335), .o(n_13365) );
oa12f80 g758782 ( .a(n_21379), .b(n_22209), .c(n_21795), .o(n_22242) );
in01f80 g743334 ( .a(n_36736), .o(n_36753) );
no02f80 g762191 ( .a(n_18215), .b(n_18214), .o(n_18240) );
no02f80 g737609 ( .a(n_42389), .b(n_42421), .o(n_42422) );
no02f80 g779582 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .o(n_1595) );
oa22f80 g739277 ( .a(n_45153), .b(n_40594), .c(n_45155), .d(delay_add_ln22_unr27_stage10_stallmux_q_31_), .o(n_40986) );
no02f80 g749071 ( .a(n_31021), .b(n_27315), .o(n_31074) );
oa22f80 FE_RC_2982_0 ( .a(n_6328), .b(n_6347), .c(n_6322), .d(n_6358), .o(n_6487) );
na02f80 g764886 ( .a(n_16137), .b(n_15632), .o(n_16177) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_25_ ( .ck(newNet_2272), .d(n_40554), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_) );
ao12f80 g765775 ( .a(n_15363), .b(n_15362), .c(n_15361), .o(n_15958) );
no02f80 g761522 ( .a(n_18828), .b(n_18798), .o(n_18954) );
oa22f80 FE_RC_401_0 ( .a(n_15154), .b(n_15321), .c(n_15153), .d(n_15284), .o(n_15433) );
in01f80 newInst_1715 ( .a(newNet_1714), .o(newNet_1715) );
na02f80 g762213 ( .a(n_18734), .b(FE_OFN750_n_45003), .o(n_18817) );
in01f80 newInst_1595 ( .a(newNet_1594), .o(newNet_1595) );
in01f80 g752271 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n_27807) );
ao12f80 g750603 ( .a(n_28761), .b(n_29353), .c(n_28742), .o(n_29385) );
in01f80 g758329 ( .a(n_22292), .o(n_22328) );
in01f80 g755205 ( .a(n_25373), .o(n_25551) );
in01f80 g779376 ( .a(n_1593), .o(n_1594) );
in01f80 newInst_1350 ( .a(newNet_1349), .o(newNet_1350) );
no02f80 g774334 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .o(n_7100) );
in01f80 g775876 ( .a(n_5346), .o(n_5347) );
na02f80 g765492 ( .a(FE_OFN765_n_15670), .b(n_15665), .o(n_15969) );
ao12f80 g781258 ( .a(n_7), .b(beta_20), .c(beta_19), .o(n_94) );
in01f80 FE_OCP_RBC2500_n_13896 ( .a(FE_OCP_RBN3528_n_13765), .o(FE_OCP_RBN2500_n_13896) );
in01f80 newInst_1710 ( .a(newNet_798), .o(newNet_1710) );
oa12f80 g772367 ( .a(n_8105), .b(n_8573), .c(n_7996), .o(n_8722) );
no02f80 g739458 ( .a(n_40663), .b(delay_add_ln22_unr27_stage10_stallmux_q_1_), .o(n_40699) );
in01f80 FE_OCP_RBC2104_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(FE_OCP_RBN2004_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN2104_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
na02f80 g742009 ( .a(n_37918), .b(n_37917), .o(n_37919) );
no02f80 g762292 ( .a(n_18498), .b(n_18450), .o(n_18779) );
in01f80 g779239 ( .a(n_1905), .o(n_1906) );
in01f80 g765016 ( .a(n_15933), .o(n_16350) );
in01f80 g749233 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n_30905) );
no02f80 g752196 ( .a(n_28035), .b(n_28034), .o(n_28114) );
in01f80 g739785 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_40494) );
na02f80 FE_RC_4064_0 ( .a(FE_RN_1768_0), .b(n_36280), .o(n_36352) );
no02f80 g742178 ( .a(n_44867), .b(n_38269), .o(n_37937) );
in01f80 g755627 ( .a(n_24636), .o(n_24637) );
in01f80 newInst_2854 ( .a(newNet_2853), .o(newNet_2854) );
na02f80 g780769 ( .a(n_490), .b(n_378), .o(n_505) );
na02f80 g773009 ( .a(n_7789), .b(n_7788), .o(n_7790) );
in01f80 g752269 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .o(n_27938) );
na02f80 g737746 ( .a(n_42233), .b(n_42202), .o(n_42259) );
in01f80 newInst_2711 ( .a(newNet_2710), .o(newNet_2711) );
in01f80 g750752 ( .a(n_29339), .o(n_29368) );
in01f80 g742983 ( .a(n_37072), .o(n_36970) );
ao12f80 g773043 ( .a(FE_OCP_RBN3461_n_7886), .b(n_8045), .c(n_7982), .o(n_8113) );
na02f80 g762361 ( .a(n_45118), .b(n_17859), .o(n_18579) );
in01f80 g747134 ( .a(n_32931), .o(n_32888) );
oa22f80 g742958 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_9_), .c(n_37082), .d(n_36151), .o(n_37319) );
na02f80 g737764 ( .a(n_42351), .b(n_42350), .o(n_42352) );
in01f80 g776031 ( .a(n_4957), .o(n_4958) );
na02f80 g737929 ( .a(n_42201), .b(n_42036), .o(n_42414) );
no02f80 g759122 ( .a(n_21312), .b(n_45070), .o(n_21350) );
na02f80 g768977 ( .a(n_12085), .b(n_12013), .o(n_12281) );
na02f80 g765960 ( .a(n_14699), .b(n_14727), .o(n_14826) );
in01f80 FE_OCPC971_n_14716 ( .a(FE_OCPN970_n_14716), .o(FE_OCPN971_n_14716) );
na02f80 g771407 ( .a(n_9641), .b(n_9640), .o(n_9786) );
na02f80 g769946 ( .a(n_11042), .b(n_10154), .o(n_11180) );
na02f80 g768356 ( .a(n_12445), .b(n_12364), .o(n_12446) );
no02f80 g742138 ( .a(n_38324), .b(n_38373), .o(n_38450) );
na02f80 g744236 ( .a(n_46209), .b(n_36838), .o(n_36880) );
oa12f80 g759026 ( .a(n_21381), .b(n_21526), .c(n_21456), .o(n_21642) );
in01f80 g743463 ( .a(n_37747), .o(n_37748) );
no02f80 g779580 ( .a(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .o(n_1434) );
ao22s80 g758201 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .c(n_22658), .d(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22813) );
in01f80 FE_OCP_RBC3597_FE_OCPN1243_n_44460 ( .a(FE_OCPN1243_n_44460), .o(FE_OCP_RBN3597_FE_OCPN1243_n_44460) );
oa12f80 g778994 ( .a(n_2196), .b(n_2195), .c(n_2194), .o(n_2228) );
in01f80 g777377 ( .a(n_3692), .o(n_3693) );
na02f80 g748843 ( .a(n_31061), .b(n_30891), .o(n_31058) );
in01f80 FE_RC_4178_0 ( .a(n_33368), .o(FE_RN_1825_0) );
in01f80 FE_OCP_RBC2636_n_38806 ( .a(n_38806), .o(FE_OCP_RBN2636_n_38806) );
oa22f80 g743324 ( .a(n_36719), .b(n_36604), .c(n_36718), .d(n_36579), .o(n_36766) );
in01f80 newInst_1551 ( .a(newNet_133), .o(newNet_1551) );
in01f80 FE_OCPC1228_n_46101 ( .a(n_46101), .o(FE_OCPN1228_n_46101) );
in01f80 g772046 ( .a(n_8898), .o(n_8899) );
no02f80 g736704 ( .a(n_43148), .b(n_43120), .o(n_43233) );
in01f80 g781261 ( .a(n_75), .o(n_76) );
na02f80 g736761 ( .a(n_43062), .b(n_43070), .o(n_43071) );
na02f80 g745603 ( .a(n_34285), .b(n_33542), .o(n_34380) );
ao12f80 g763951 ( .a(n_16583), .b(n_16560), .c(n_16562), .o(n_16640) );
oa22f80 FE_RC_27_0 ( .a(FE_OFN84_n_46137), .b(n_6479), .c(FE_OFN806_n_46196), .d(n_46993), .o(n_46181) );
na02f80 g759983 ( .a(n_20606), .b(n_20529), .o(n_20607) );
in01f80 g740211 ( .a(n_39861), .o(n_39898) );
in01f80 FE_OCP_DRV_C1554_n_19314 ( .a(FE_OCP_DRV_N1553_n_19314), .o(FE_OCP_DRV_N1554_n_19314) );
oa22f80 g764135 ( .a(n_16886), .b(n_16132), .c(n_16885), .d(n_16131), .o(n_17014) );
na02f80 g748521 ( .a(n_31446), .b(FE_OCP_DRV_N1606_n_31445), .o(n_31519) );
no02f80 g751994 ( .a(n_28793), .b(n_28942), .o(n_28955) );
in01f80 FE_OCP_RBC3841_n_19419 ( .a(n_19419), .o(FE_OCP_RBN3841_n_19419) );
na02f80 g770090 ( .a(n_10893), .b(n_10746), .o(n_10952) );
in01f80 g748904 ( .a(n_32498), .o(n_32482) );
no02f80 g777763 ( .a(n_3270), .b(n_2486), .o(n_3316) );
no02f80 g743071 ( .a(n_37085), .b(n_36929), .o(n_37139) );
ao22s80 FE_RC_3890_0 ( .a(n_28628), .b(n_29035), .c(n_28629), .d(n_29034), .o(n_29143) );
in01f80 g736410 ( .a(n_43820), .o(n_43821) );
in01f80 g739109 ( .a(n_40997), .o(n_41051) );
in01f80 g754513 ( .a(n_25566), .o(n_25629) );
in01f80 g750838 ( .a(n_29167), .o(n_29160) );
no02f80 g765783 ( .a(n_14905), .b(n_14758), .o(n_14941) );
in01f80 g780208 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_7_), .o(n_1038) );
in01f80 g763457 ( .a(n_17311), .o(n_17312) );
na02f80 FE_RC_3998_0 ( .a(n_29929), .b(FE_RN_1733_0), .o(n_30298) );
no02f80 g757552 ( .a(FE_OCP_RBN3817_n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .o(n_22799) );
in01f80 g757882 ( .a(n_22238), .o(n_22239) );
in01f80 g774429 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .o(n_6506) );
in01f80 g769304 ( .a(n_11669), .o(n_11759) );
no02f80 g748943 ( .a(n_31198), .b(n_31197), .o(n_31230) );
in01f80 g740340 ( .a(n_40353), .o(n_40354) );
in01f80 g738234 ( .a(n_41956), .o(n_42374) );
na02f80 g766691 ( .a(n_13850), .b(n_12799), .o(n_13980) );
no02f80 g770068 ( .a(n_10898), .b(n_10875), .o(n_10932) );
in01f80 g770584 ( .a(n_10280), .o(n_10360) );
in01f80 newInst_1354 ( .a(newNet_1353), .o(newNet_1354) );
no02f80 g755890 ( .a(n_25570), .b(n_25604), .o(n_25689) );
oa12f80 g741920 ( .a(n_38073), .b(n_38074), .c(n_37941), .o(n_38126) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_20_ ( .ck(newNet_3224), .d(n_36439), .o(delay_add_ln22_unr23_stage9_stallmux_q_20_) );
na02f80 g754458 ( .a(n_26831), .b(n_26832), .o(n_26833) );
no02f80 g754968 ( .a(n_25182), .b(n_25147), .o(n_25183) );
na03f80 g774155 ( .a(n_6619), .b(n_6656), .c(n_6543), .o(n_6734) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_26_ ( .ck(newNet_3609), .d(n_17782), .o(delay_add_ln22_unr11_stage5_stallmux_q_26_) );
in01f80 g744572 ( .a(n_35333), .o(n_35334) );
no02f80 g742010 ( .a(n_37951), .b(n_37950), .o(n_37952) );
in01f80 FE_OCP_RBC3619_n_15135 ( .a(n_15135), .o(FE_OCP_RBN3619_n_15135) );
in01f80 g765589 ( .a(n_15748), .o(n_15512) );
no02f80 g764445 ( .a(n_16158), .b(n_16194), .o(n_16288) );
in01f80 newInst_728 ( .a(newNet_727), .o(newNet_728) );
in01f80 g768327 ( .a(n_12502), .o(n_12503) );
na02f80 g771473 ( .a(n_9121), .b(n_9041), .o(n_9204) );
na02f80 g778238 ( .a(n_47025), .b(n_2766), .o(n_2799) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_18_ ( .ck(newNet_2570), .d(n_27622), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_) );
no02f80 g775437 ( .a(n_5742), .b(n_4819), .o(n_5874) );
in01f80 g747407 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .o(n_32622) );
na02f80 g765055 ( .a(n_16133), .b(n_16175), .o(n_16176) );
no02f80 g773038 ( .a(n_8049), .b(n_8060), .o(n_8120) );
na02f80 g775828 ( .a(n_5339), .b(n_5294), .o(n_5295) );
oa12f80 g757468 ( .a(n_23344), .b(n_23343), .c(n_23342), .o(n_23954) );
no02f80 g754326 ( .a(n_25783), .b(n_25445), .o(n_25828) );
na02f80 g750613 ( .a(n_29491), .b(n_28349), .o(n_29583) );
no02f80 g752933 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_), .o(n_28076) );
in01f80 g745354 ( .a(n_34262), .o(n_34263) );
na02f80 g748287 ( .a(FE_OCP_RBN3735_n_31819), .b(FE_OCP_RBN2933_n_31010), .o(n_32044) );
na02f80 g773929 ( .a(n_7001), .b(n_6903), .o(n_7060) );
no02f80 g776115 ( .a(n_44862), .b(n_5009), .o(n_5010) );
in01f80 g755667 ( .a(n_26419), .o(n_25524) );
na02f80 g751904 ( .a(n_28940), .b(n_28939), .o(n_28941) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_4_ ( .ck(newNet_1801), .d(n_16411), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_) );
in01f80 FE_OCP_RBC2637_n_38806 ( .a(FE_OCP_RBN2636_n_38806), .o(FE_OCP_RBN2637_n_38806) );
na02f80 g773948 ( .a(n_7000), .b(n_47210), .o(n_7001) );
na02f80 g771052 ( .a(n_9360), .b(n_8362), .o(n_9504) );
na02f80 g778214 ( .a(n_2829), .b(n_2665), .o(n_2860) );
ao22s80 FE_RC_607_0 ( .a(n_38183), .b(n_38499), .c(n_38184), .d(n_38500), .o(n_38569) );
in01f80 g746152 ( .a(n_35109), .o(n_35190) );
in01f80 newInst_1161 ( .a(newNet_1160), .o(newNet_1161) );
no02f80 g755531 ( .a(n_24650), .b(n_22393), .o(n_24651) );
no02f80 g775965 ( .a(n_5101), .b(n_3625), .o(n_5149) );
na02f80 g765068 ( .a(n_15240), .b(n_15283), .o(n_15429) );
in01f80 g736997 ( .a(n_43297), .o(n_43391) );
in01f80 g774894 ( .a(n_6419), .o(n_6392) );
in01f80 g768463 ( .a(n_12434), .o(n_12435) );
in01f80 g762814 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_23_), .o(n_17692) );
in01f80 fopt783670 ( .a(n_45322), .o(n_45321) );
no02f80 g768916 ( .a(FE_OCPN867_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_12_), .o(n_12055) );
no02f80 g741473 ( .a(n_38767), .b(n_38766), .o(n_38768) );
no02f80 g758261 ( .a(FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_10_), .o(n_22695) );
na02f80 g772491 ( .a(n_8469), .b(n_8468), .o(n_8470) );
na02f80 g755892 ( .a(n_25741), .b(n_25680), .o(n_25950) );
na02f80 g742460 ( .a(n_37562), .b(n_37057), .o(n_37607) );
in01f80 g762769 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_18_), .o(n_17892) );
oa12f80 g761181 ( .a(n_18310), .b(FE_OCP_RBN3826_n_18951), .c(n_18339), .o(n_19062) );
in01f80 FE_OCP_RBC3100_n_22502 ( .a(n_22502), .o(FE_OCP_RBN3100_n_22502) );
in01f80 newInst_3722 ( .a(newNet_3721), .o(newNet_3722) );
ao12f80 g768509 ( .a(n_12370), .b(n_45659), .c(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .o(n_12488) );
na02f80 g763668 ( .a(n_17212), .b(n_17093), .o(n_17609) );
ao12f80 g741929 ( .a(n_38070), .b(n_38092), .c(n_38069), .o(n_38820) );
no02f80 g774469 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n_6742) );
in01f80 newInst_535 ( .a(newNet_358), .o(newNet_535) );
no02f80 FE_RC_3633_0 ( .a(n_23278), .b(n_24291), .o(FE_RN_1592_0) );
na02f80 FE_RC_3982_0 ( .a(n_13945), .b(n_13944), .o(FE_RN_1726_0) );
oa12f80 g779328 ( .a(n_1616), .b(n_1690), .c(n_1644), .o(n_1699) );
na02f80 g742413 ( .a(n_37742), .b(n_37741), .o(n_37777) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_8_ ( .ck(newNet_2895), .d(n_5379), .o(delay_add_ln22_unr5_stage3_stallmux_q_8_) );
in01f80 newInst_462 ( .a(newNet_461), .o(newNet_462) );
na02f80 g758808 ( .a(n_21789), .b(n_21788), .o(n_21871) );
in01f80 g763390 ( .a(n_17036), .o(n_17135) );
in01f80 newInst_1672 ( .a(newNet_554), .o(newNet_1672) );
no02f80 g759436 ( .a(n_21699), .b(n_21254), .o(n_21673) );
na02f80 g737016 ( .a(n_43230), .b(n_42596), .o(n_43493) );
no02f80 g750059 ( .a(n_29869), .b(FE_OCP_RBN2265_n_29033), .o(n_30010) );
na02f80 g748836 ( .a(n_31296), .b(n_31231), .o(n_31354) );
na02f80 g748378 ( .a(n_31476), .b(n_31504), .o(n_31522) );
in01f80 g752925 ( .a(n_28156), .o(n_28077) );
na02f80 g768419 ( .a(n_12404), .b(FE_OCPN1002_n_45660), .o(n_12461) );
na02f80 g741633 ( .a(n_38569), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38584) );
in01f80 g755617 ( .a(n_24598), .o(n_24646) );
in01f80 g748664 ( .a(n_31484), .o(n_31485) );
na02f80 g763748 ( .a(n_16708), .b(n_16668), .o(n_16731) );
na02f80 g775097 ( .a(n_6025), .b(n_5791), .o(n_6049) );
na02f80 g738483 ( .a(n_41582), .b(n_41292), .o(n_41830) );
in01f80 g767620 ( .a(n_12940), .o(n_12941) );
in01f80 g753749 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_1_), .o(n_28034) );
in01f80 newInst_3502 ( .a(newNet_3501), .o(newNet_3502) );
in01f80 newInst_32 ( .a(newNet_0), .o(newNet_32) );
in01f80 g747839 ( .a(n_33701), .o(n_33532) );
no02f80 g739702 ( .a(n_40471), .b(n_40522), .o(n_40523) );
in01f80 g754121 ( .a(n_26061), .o(n_26062) );
in01f80 g767742 ( .a(n_13045), .o(n_13046) );
oa22f80 FE_RC_1391_0 ( .a(n_46956), .b(n_27315), .c(n_31017), .d(n_27366), .o(n_31101) );
no02f80 g772831 ( .a(n_8022), .b(n_8070), .o(n_8175) );
no02f80 g760969 ( .a(n_19300), .b(n_19350), .o(n_19420) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_18_ ( .ck(newNet_1626), .d(n_27200), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_18_) );
na02f80 g769202 ( .a(n_11897), .b(n_11960), .o(n_12470) );
oa12f80 g745273 ( .a(n_36083), .b(FE_OCP_RBN2994_n_35539), .c(n_36118), .o(n_36176) );
oa12f80 g765913 ( .a(n_14744), .b(n_14743), .c(n_14898), .o(n_14916) );
in01f80 FE_OCP_RBC2861_n_10399 ( .a(FE_OCP_RBN2859_n_10399), .o(FE_OCP_RBN2861_n_10399) );
no02f80 g770178 ( .a(n_10669), .b(n_10601), .o(n_10791) );
in01f80 FE_OCP_RBC2546_n_44944 ( .a(n_44944), .o(FE_OCP_RBN2546_n_44944) );
oa22f80 g780169 ( .a(n_997), .b(n_1098), .c(n_45819), .d(n_1099), .o(n_1124) );
in01f80 g752391 ( .a(n_27884), .o(n_27937) );
no02f80 g768600 ( .a(n_12296), .b(n_11885), .o(n_12312) );
na02f80 g773515 ( .a(n_7436), .b(n_7426), .o(n_7500) );
na02f80 g772795 ( .a(n_8136), .b(n_8135), .o(n_8182) );
na02f80 g749870 ( .a(FE_OCP_RBN3010_n_31117), .b(n_31213), .o(n_31570) );
oa22f80 g753700 ( .a(n_27096), .b(n_26891), .c(n_27095), .d(n_26890), .o(n_27165) );
no02f80 g757046 ( .a(n_23700), .b(n_23699), .o(n_23748) );
in01f80 FE_OCP_RBC2165_n_28249 ( .a(n_28249), .o(FE_OCP_RBN2165_n_28249) );
na02f80 g770312 ( .a(FE_OCP_RBN2936_n_10626), .b(n_10682), .o(n_10719) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_7_ ( .ck(newNet_2900), .d(n_5323), .o(delay_add_ln22_unr5_stage3_stallmux_q_7_) );
no02f80 g750319 ( .a(n_29705), .b(n_29688), .o(n_29751) );
in01f80 g744662 ( .a(n_36598), .o(n_36619) );
na02f80 g746956 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_33289) );
in01f80 g759127 ( .a(n_21487), .o(n_21488) );
na02f80 g756213 ( .a(n_24083), .b(n_24071), .o(n_24181) );
in01f80 FE_RC_1069_0 ( .a(n_12311), .o(FE_RN_315_0) );
oa12f80 g738353 ( .a(n_41408), .b(n_41517), .c(n_41452), .o(n_41596) );
in01f80 g741549 ( .a(n_38724), .o(n_38725) );
na02f80 g778276 ( .a(n_2623), .b(n_2622), .o(n_2724) );
in01f80 g744768 ( .a(n_35198), .o(n_35199) );
no02f80 g738980 ( .a(n_41207), .b(n_40989), .o(n_41241) );
na02f80 g747158 ( .a(n_32867), .b(n_32905), .o(n_32970) );
na02f80 g748690 ( .a(n_31183), .b(n_31271), .o(n_31301) );
no02f80 g742239 ( .a(FE_OCP_RBN3425_n_44881), .b(n_38047), .o(n_38078) );
in01f80 g764591 ( .a(n_16541), .o(n_16542) );
no02f80 g748638 ( .a(n_31488), .b(n_31490), .o(n_31491) );
in01f80 g749836 ( .a(n_31224), .o(n_31187) );
na02f80 g759605 ( .a(n_20684), .b(n_20473), .o(n_20767) );
in01f80 newInst_3073 ( .a(newNet_3072), .o(newNet_3073) );
in01f80 g776014 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_5_), .o(n_5139) );
no02f80 g744296 ( .a(n_44180), .b(n_35897), .o(n_36001) );
ao12f80 g767711 ( .a(n_13204), .b(n_13084), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n_13320) );
in01f80 g756733 ( .a(n_23431), .o(n_23432) );
no02f80 g769394 ( .a(n_44336), .b(n_10293), .o(n_11473) );
in01f80 g766189 ( .a(n_14475), .o(n_14476) );
na02f80 g777629 ( .a(n_3414), .b(n_3191), .o(n_3415) );
na02f80 g769231 ( .a(n_11627), .b(FE_OCP_RBN2949_n_10852), .o(n_11715) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_19_ ( .ck(newNet_568), .d(n_17752), .o(delay_xor_ln22_unr12_stage5_stallmux_q_19_) );
in01f80 newInst_1829 ( .a(newNet_1828), .o(newNet_1829) );
in01f80 g777418 ( .a(n_3690), .o(n_3794) );
no02f80 g750686 ( .a(n_29279), .b(n_28800), .o(n_29280) );
in01f80 g738521 ( .a(n_41583), .o(n_41624) );
in01f80 g757535 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_24_), .o(n_23653) );
in01f80 FE_OCP_RBC3442_n_37945 ( .a(n_37945), .o(FE_OCP_RBN3442_n_37945) );
in01f80 newInst_669 ( .a(newNet_371), .o(newNet_669) );
na02f80 g745741 ( .a(n_34479), .b(n_34328), .o(n_34569) );
na02f80 g738464 ( .a(n_41387), .b(n_41473), .o(n_41513) );
in01f80 g777506 ( .a(n_4556), .o(n_4875) );
no02f80 g783678 ( .a(n_15856), .b(n_15942), .o(n_45332) );
na02f80 g755586 ( .a(n_24451), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24476) );
oa22f80 g784354 ( .a(FE_OFN86_n_46137), .b(n_6043), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_6063), .o(n_46160) );
in01f80 newInst_2257 ( .a(newNet_2256), .o(newNet_2257) );
na02f80 g759744 ( .a(n_47175), .b(n_45065), .o(n_20348) );
in01f80 newInst_1593 ( .a(newNet_994), .o(newNet_1593) );
na02f80 g756996 ( .a(n_47337), .b(n_23267), .o(n_23287) );
oa12f80 g751266 ( .a(n_29759), .b(n_29758), .c(n_29757), .o(n_30095) );
in01f80 FE_OCP_RBC2489_n_3338 ( .a(FE_OCP_RBN2487_n_3338), .o(FE_OCP_RBN2489_n_3338) );
no02f80 g779130 ( .a(n_2015), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .o(n_2061) );
na02f80 g748436 ( .a(n_31730), .b(n_31107), .o(n_31721) );
in01f80 newInst_1872 ( .a(newNet_1871), .o(newNet_1872) );
na02f80 FE_RC_3096_0 ( .a(n_30526), .b(n_30527), .o(FE_RN_1368_0) );
na02f80 g746722 ( .a(n_33234), .b(n_33097), .o(n_33235) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_1_ ( .ck(newNet_3321), .d(n_31008), .o(delay_add_ln22_unr20_stage8_stallmux_q_1_) );
na02f80 g776671 ( .a(n_4214), .b(n_4247), .o(n_4434) );
in01f80 g770736 ( .a(n_10190), .o(n_10191) );
no02f80 g736645 ( .a(n_43475), .b(n_43352), .o(n_43526) );
na02f80 g767922 ( .a(n_12669), .b(n_12654), .o(n_12799) );
oa12f80 FE_RC_2187_0 ( .a(FE_RN_782_0), .b(n_22750), .c(n_22801), .o(n_22794) );
na02f80 g781316 ( .a(beta_31), .b(beta_25), .o(n_103) );
ao12f80 g761170 ( .a(n_19084), .b(n_19083), .c(n_19082), .o(n_21028) );
no02f80 g756923 ( .a(n_23703), .b(n_23702), .o(n_23751) );
na02f80 g744861 ( .a(n_35033), .b(n_35010), .o(n_35099) );
na02f80 FE_RC_3103_0 ( .a(FE_RN_1371_0), .b(n_21233), .o(FE_RN_1372_0) );
in01f80 g743475 ( .a(n_37725), .o(n_37726) );
in01f80 g742671 ( .a(n_37416), .o(n_37417) );
ao12f80 g750575 ( .a(n_29443), .b(n_29396), .c(n_29322), .o(n_29542) );
oa12f80 g765157 ( .a(n_15879), .b(n_15827), .c(FE_OFN765_n_15670), .o(n_15974) );
in01f80 newInst_2220 ( .a(newNet_2219), .o(newNet_2220) );
ao12f80 g743868 ( .a(n_46250), .b(n_36434), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37138) );
in01f80 g741020 ( .a(n_39209), .o(n_39210) );
in01f80 newInst_213 ( .a(newNet_60), .o(newNet_213) );
oa12f80 g739867 ( .a(n_39908), .b(n_40200), .c(n_39902), .o(n_40261) );
in01f80 g741111 ( .a(n_39048), .o(n_39049) );
na02f80 g740144 ( .a(FE_OCP_RBN3721_n_39913), .b(n_39459), .o(n_40187) );
in01f80 g779405 ( .a(n_1513), .o(n_1547) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_13_ ( .ck(newNet_2119), .d(n_5913), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_) );
in01f80 FE_OCPC873_n_44672 ( .a(n_44672), .o(FE_OCPN873_n_44672) );
no02f80 g746350 ( .a(n_34868), .b(n_34867), .o(n_34916) );
in01f80 FE_OCP_RBC1342_n_19077 ( .a(FE_OCP_RBN1341_n_19077), .o(FE_OCP_RBN1342_n_19077) );
ao12f80 g779507 ( .a(n_1554), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .o(n_1609) );
in01f80 g750996 ( .a(n_29892), .o(n_28995) );
ao12f80 g756847 ( .a(n_23331), .b(n_23266), .c(delay_add_ln22_unr14_stage6_stallmux_q_9_), .o(n_23506) );
na02f80 g754919 ( .a(n_25270), .b(FE_OCP_RBN2307_n_24288), .o(n_25389) );
in01f80 newInst_2113 ( .a(newNet_2112), .o(newNet_2113) );
in01f80 g760937 ( .a(n_19386), .o(n_19387) );
in01f80 g736337 ( .a(n_43854), .o(n_43855) );
na02f80 g775672 ( .a(n_5658), .b(n_5727), .o(n_5688) );
no02f80 g763292 ( .a(n_17391), .b(n_17390), .o(n_17392) );
in01f80 FE_OCP_RBC3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN3361_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
no02f80 g760792 ( .a(n_19592), .b(n_19602), .o(n_19593) );
in01f80 newInst_3022 ( .a(newNet_3021), .o(newNet_3022) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_3_ ( .ck(newNet_559), .d(n_16804), .o(delay_xor_ln22_unr12_stage5_stallmux_q_3_) );
no02f80 g748127 ( .a(n_31904), .b(n_31835), .o(n_31951) );
no03m80 FE_RC_1656_0 ( .a(n_23378), .b(n_23022), .c(n_23379), .o(n_23411) );
in01f80 g775944 ( .a(n_4858), .o(n_4903) );
ao12f80 g780322 ( .a(n_831), .b(n_851), .c(n_45809), .o(n_908) );
in01f80 g766751 ( .a(n_16246), .o(n_14433) );
ao12f80 g752249 ( .a(n_28001), .b(FE_OCP_RBN2126_n_44734), .c(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n_28030) );
in01f80 g746408 ( .a(n_33427), .o(n_33428) );
in01f80 FE_RC_205_0 ( .a(FE_RN_68_0), .o(n_11765) );
in01f80 g775137 ( .a(n_6080), .o(n_6006) );
in01f80 newInst_3438 ( .a(newNet_2577), .o(newNet_3438) );
no02f80 FE_RC_985_0 ( .a(FE_RN_283_0), .b(FE_RN_282_0), .o(FE_RN_284_0) );
in01f80 g749683 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_), .o(n_32356) );
in01f80 g738046 ( .a(n_42148), .o(n_42391) );
no02f80 g766550 ( .a(n_14457), .b(n_14110), .o(n_14531) );
na02f80 g738525 ( .a(FE_OCP_RBN2312_n_41420), .b(n_41175), .o(n_41546) );
oa22f80 g752512 ( .a(n_27665), .b(n_24350), .c(n_27644), .d(n_27796), .o(n_27708) );
in01f80 g777651 ( .a(n_3505), .o(n_3506) );
in01f80 g775396 ( .a(n_5888), .o(n_5911) );
oa22f80 FE_RC_3148_0 ( .a(n_21326), .b(n_21443), .c(n_21442), .d(n_21327), .o(n_21581) );
in01f80 g779428 ( .a(n_1460), .o(n_1461) );
no02f80 g779421 ( .a(n_1501), .b(n_1515), .o(n_1502) );
na02f80 g767411 ( .a(n_13232), .b(FE_OCP_RBN3419_n_12739), .o(n_13244) );
in01f80 g755753 ( .a(n_24463), .o(n_24489) );
no02f80 g769903 ( .a(n_10966), .b(n_10917), .o(n_11011) );
in01f80 FE_OCP_RBC2855_n_10112 ( .a(n_10112), .o(FE_OCP_RBN2855_n_10112) );
na02f80 g765587 ( .a(n_15599), .b(n_14434), .o(n_16136) );
in01f80 g751514 ( .a(n_29175), .o(n_29176) );
ao22s80 FE_RC_862_0 ( .a(FE_OCP_RBN2559_n_44576), .b(n_9584), .c(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .d(FE_OCP_RBN2747_n_9584), .o(n_9747) );
no02f80 g754852 ( .a(n_25359), .b(n_25358), .o(n_25360) );
in01f80 g739437 ( .a(n_40766), .o(n_40721) );
ao12f80 g781090 ( .a(n_248), .b(n_247), .c(n_246), .o(n_424) );
in01f80 newInst_1152 ( .a(newNet_1151), .o(newNet_1152) );
na02f80 g760783 ( .a(n_20137), .b(n_19762), .o(n_20155) );
na02f80 g778248 ( .a(n_45506), .b(n_2480), .o(n_2692) );
na02f80 g756586 ( .a(n_23601), .b(n_23636), .o(n_24001) );
na02f80 g770374 ( .a(n_10689), .b(n_9829), .o(n_10720) );
no02f80 FE_RC_2136_0 ( .a(FE_RN_746_0), .b(n_26553), .o(FE_RN_747_0) );
no02f80 g768364 ( .a(n_12464), .b(delay_add_ln22_unr8_stage4_stallmux_q_13_), .o(n_12483) );
na02f80 g779144 ( .a(n_1870), .b(n_1442), .o(n_1958) );
na02f80 g748828 ( .a(n_31178), .b(n_31200), .o(n_31234) );
no02f80 g743251 ( .a(n_36865), .b(n_36883), .o(n_36904) );
in01f80 FE_OCPC1011_n_7802 ( .a(FE_OCPN1010_n_7802), .o(FE_OCPN1011_n_7802) );
in01f80 g774790 ( .a(n_6354), .o(n_6355) );
na02f80 g746369 ( .a(n_33412), .b(n_33434), .o(n_33491) );
in01f80 FE_RC_4082_0 ( .a(n_16923), .o(FE_RN_1782_0) );
in01f80 FE_OCPC1041_n_3673 ( .a(n_3673), .o(FE_OCPN1041_n_3673) );
oa12f80 g755064 ( .a(n_25196), .b(n_25715), .c(n_25217), .o(n_25803) );
no02f80 g769608 ( .a(n_11351), .b(n_11269), .o(n_11352) );
in01f80 newInst_2065 ( .a(newNet_2064), .o(newNet_2065) );
no02f80 g775168 ( .a(n_5818), .b(n_4759), .o(n_5926) );
na02f80 g780828 ( .a(n_567), .b(n_427), .o(n_614) );
no02f80 g773872 ( .a(n_7083), .b(FE_OCPN895_n_6521), .o(n_7087) );
in01f80 g757147 ( .a(n_23803), .o(n_24059) );
ao12f80 g741828 ( .a(n_38387), .b(n_38386), .c(n_38385), .o(n_39324) );
ao22s80 g736355 ( .a(n_43836), .b(n_43598), .c(n_43837), .d(n_43597), .o(n_43867) );
na02f80 g755590 ( .a(n_24637), .b(n_24713), .o(n_24780) );
in01f80 g758736 ( .a(n_21818), .o(n_21833) );
in01f80 g752627 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_15_), .o(n_28473) );
in01f80 g738008 ( .a(n_42189), .o(n_42192) );
in01f80 newInst_972 ( .a(newNet_971), .o(newNet_972) );
no02f80 g738919 ( .a(n_41280), .b(n_41279), .o(n_41281) );
in01f80 newInst_1614 ( .a(newNet_1613), .o(newNet_1614) );
no02f80 g749949 ( .a(n_30050), .b(n_30116), .o(n_30143) );
ao22s80 FE_RC_3331_0 ( .a(FE_OFN779_n_17093), .b(n_19008), .c(n_17783), .d(n_19033), .o(n_19110) );
in01f80 FE_RC_2255_0 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(FE_RN_832_0) );
na02f80 g774012 ( .a(n_6889), .b(n_6597), .o(n_6890) );
na02f80 g772881 ( .a(n_7930), .b(n_8676), .o(n_7981) );
na02f80 g768751 ( .a(n_12125), .b(n_12124), .o(n_12126) );
in01f80 g748643 ( .a(n_33362), .o(n_33396) );
ao12f80 g766391 ( .a(n_14028), .b(n_14026), .c(n_14101), .o(n_14133) );
in01f80 g746982 ( .a(n_32911), .o(n_32999) );
na02f80 g780893 ( .a(n_374), .b(n_385), .o(n_409) );
in01f80 g773499 ( .a(n_7519), .o(n_7520) );
na02f80 g756624 ( .a(n_24192), .b(n_24152), .o(n_24193) );
na02f80 g744262 ( .a(n_44180), .b(n_34765), .o(n_35590) );
in01f80 g780048 ( .a(n_1245), .o(n_1246) );
no02f80 g777380 ( .a(n_3652), .b(n_3749), .o(n_3792) );
no02f80 g753667 ( .a(n_26596), .b(n_26562), .o(n_26563) );
in01f80 FE_OCP_RBC1153_n_29053 ( .a(n_29053), .o(FE_OCP_RBN1153_n_29053) );
no02f80 g753778 ( .a(n_26519), .b(n_26336), .o(n_26580) );
na02f80 g775497 ( .a(n_5457), .b(n_4556), .o(n_5568) );
in01f80 g748734 ( .a(n_31379), .o(n_31380) );
oa12f80 g759792 ( .a(n_21622), .b(n_21374), .c(n_21562), .o(n_21563) );
oa12f80 g752848 ( .a(n_26982), .b(n_27047), .c(n_26913), .o(n_27058) );
no02f80 g779565 ( .a(n_1471), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n_1493) );
in01f80 g749789 ( .a(n_31313), .o(n_31314) );
in01f80 g758011 ( .a(n_22338), .o(n_22339) );
in01f80 FE_OCPC1856_n_33341 ( .a(FE_OCPN1855_n_33341), .o(FE_OCPN1856_n_33341) );
in01f80 newInst_3312 ( .a(newNet_3311), .o(newNet_3312) );
na02f80 g743863 ( .a(n_46250), .b(n_46236), .o(n_37027) );
no02f80 g783840 ( .a(n_18237), .b(n_45527), .o(n_45528) );
oa12f80 g778400 ( .a(n_2049), .b(n_45488), .c(n_2017), .o(n_2528) );
in01f80 g778688 ( .a(n_2745), .o(n_2705) );
no02f80 g778678 ( .a(FE_OCP_RBN2294_n_2438), .b(n_2472), .o(n_2661) );
no02f80 g773034 ( .a(n_7679), .b(n_7666), .o(n_7803) );
in01f80 newInst_2925 ( .a(newNet_2924), .o(newNet_2925) );
no02f80 g739036 ( .a(n_41093), .b(n_41042), .o(n_41144) );
ao12f80 g761526 ( .a(n_19549), .b(n_19548), .c(n_19547), .o(n_19983) );
in01f80 g769127 ( .a(n_11743), .o(n_11744) );
na02f80 g776870 ( .a(n_4010), .b(n_4064), .o(n_4281) );
no02f80 g755853 ( .a(n_24252), .b(n_23849), .o(n_24294) );
in01f80 g746950 ( .a(n_32939), .o(n_32940) );
na02f80 g779303 ( .a(n_1699), .b(n_1698), .o(n_1700) );
in01f80 g740742 ( .a(n_39889), .o(n_39520) );
no02f80 g763818 ( .a(n_17154), .b(n_17260), .o(n_18141) );
in01f80 g759858 ( .a(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_22089) );
na02f80 FE_RC_2704_0 ( .a(n_7536), .b(FE_RN_1136_0), .o(n_8409) );
no02f80 g739161 ( .a(n_40942), .b(n_40941), .o(n_40957) );
in01f80 g775059 ( .a(n_6041), .o(n_6064) );
no02f80 g746608 ( .a(FE_OCP_RBN2600_n_34388), .b(n_34497), .o(n_34815) );
in01f80 newInst_1292 ( .a(newNet_1291), .o(newNet_1292) );
in01f80 newInst_2689 ( .a(newNet_2688), .o(newNet_2689) );
in01f80 g746259 ( .a(n_33728), .o(n_33750) );
in01f80 g739743 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_18_), .o(n_40514) );
ao22s80 FE_RC_3882_0 ( .a(n_20690), .b(n_20730), .c(n_20647), .d(n_20731), .o(n_20886) );
in01f80 g748950 ( .a(n_31194), .o(n_31195) );
in01f80 g759130 ( .a(n_21977), .o(n_21978) );
na02f80 g745640 ( .a(n_34369), .b(n_33662), .o(n_34627) );
in01f80 FE_OFC797_n_46285 ( .a(n_46285), .o(FE_OFN797_n_46285) );
in01f80 newInst_1853 ( .a(newNet_1852), .o(newNet_1853) );
na02f80 g768074 ( .a(FE_OCP_RBN3414_n_12739), .b(n_12224), .o(n_12811) );
no02f80 g766380 ( .a(n_14191), .b(n_14190), .o(n_14192) );
in01f80 g743837 ( .a(n_35878), .o(n_35876) );
na02f80 g740834 ( .a(n_39291), .b(n_39012), .o(n_39354) );
in01f80 FE_OCPC1387_n_11041 ( .a(n_11041), .o(FE_OCPN1387_n_11041) );
in01f80 g768527 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_19_), .o(n_12338) );
no02f80 g743785 ( .a(n_36046), .b(n_35693), .o(n_36108) );
no02f80 g750131 ( .a(FE_OCPN1786_n_30134), .b(n_30399), .o(n_30443) );
no02f80 g736752 ( .a(n_43276), .b(n_43174), .o(n_43277) );
na02f80 g741653 ( .a(n_38579), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38623) );
in01f80 FE_RC_2675_0 ( .a(n_3790), .o(FE_RN_1118_0) );
na02f80 g749863 ( .a(n_31311), .b(n_30718), .o(n_31526) );
in01f80 g738124 ( .a(n_42052), .o(n_42053) );
na02f80 g765243 ( .a(n_15407), .b(n_15335), .o(n_15453) );
oa22f80 FE_RC_1168_0 ( .a(n_32687), .b(n_32647), .c(n_32612), .d(FE_OCP_RBN2130_n_32647), .o(n_32770) );
na02f80 g777964 ( .a(n_3045), .b(n_3044), .o(n_3046) );
na02f80 g748600 ( .a(n_31492), .b(n_27536), .o(n_31494) );
in01f80 newInst_2397 ( .a(newNet_2396), .o(newNet_2397) );
oa12f80 g781209 ( .a(n_166), .b(n_165), .c(beta_3), .o(n_501) );
in01f80 FE_RC_1165_0 ( .a(n_28012), .o(FE_RN_352_0) );
na02f80 g762144 ( .a(n_18817), .b(n_18772), .o(n_19610) );
in01f80 FE_OCP_RBC2981_n_26591 ( .a(n_26591), .o(FE_OCP_RBN2981_n_26591) );
na02f80 g764665 ( .a(n_15809), .b(n_15855), .o(n_15992) );
na02f80 g767684 ( .a(n_12956), .b(n_13000), .o(n_13022) );
no02f80 g748307 ( .a(n_31605), .b(n_31610), .o(n_31736) );
in01f80 drc784752 ( .a(n_47235), .o(n_47236) );
in01f80 FE_RC_4043_0 ( .a(FE_OCP_DRV_N1603_n_19961), .o(FE_RN_1757_0) );
in01f80 newInst_475 ( .a(newNet_474), .o(newNet_475) );
na02f80 g754088 ( .a(n_26100), .b(n_26027), .o(n_26101) );
no02f80 g737557 ( .a(n_42266), .b(n_42221), .o(n_42508) );
no02f80 g772815 ( .a(n_7985), .b(n_8091), .o(n_8092) );
in01f80 newInst_239 ( .a(newNet_9), .o(newNet_239) );
in01f80 g775912 ( .a(n_5087), .o(n_5125) );
na02f80 g770621 ( .a(n_10418), .b(n_10489), .o(n_10565) );
no02f80 g767791 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_30_), .o(n_13120) );
no02f80 g756086 ( .a(n_24246), .b(FE_OCP_RBN2279_n_24199), .o(n_24247) );
in01f80 g755057 ( .a(n_25661), .o(n_25662) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_0_ ( .ck(newNet_1773), .d(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(cordic_combinational_sub_ln23_0_unr20_z_0_) );
in01f80 newInst_275 ( .a(newNet_274), .o(newNet_275) );
no02f80 g777702 ( .a(n_3279), .b(n_3173), .o(n_3327) );
no03m80 g767589 ( .a(n_12857), .b(n_13136), .c(n_12854), .o(n_13306) );
oa12f80 g773540 ( .a(n_6783), .b(n_7434), .c(n_6936), .o(n_7480) );
no02f80 g777936 ( .a(n_3111), .b(n_3087), .o(n_3088) );
na02f80 g736627 ( .a(n_43156), .b(n_43158), .o(n_43159) );
in01f80 g748351 ( .a(n_31914), .o(n_31915) );
in01f80 g746892 ( .a(n_33057), .o(n_33102) );
na02f80 g778059 ( .a(n_2960), .b(n_2959), .o(n_2961) );
ao12f80 g774936 ( .a(n_5241), .b(n_6160), .c(n_5368), .o(n_6209) );
in01f80 g771020 ( .a(n_9890), .o(n_9901) );
na02f80 g756636 ( .a(n_23555), .b(n_23554), .o(n_23631) );
no02f80 g740594 ( .a(n_39576), .b(n_45840), .o(n_39607) );
no02f80 g738214 ( .a(n_41939), .b(n_41750), .o(n_41962) );
in01f80 newInst_571 ( .a(newNet_570), .o(newNet_571) );
oa22f80 g739753 ( .a(n_40423), .b(n_40324), .c(n_40424), .d(n_40325), .o(n_40465) );
oa12f80 g781221 ( .a(n_146), .b(n_78), .c(n_12), .o(n_162) );
no02f80 g755240 ( .a(n_24977), .b(n_24976), .o(n_24978) );
ao22s80 g750386 ( .a(n_29610), .b(n_29633), .c(n_29584), .d(n_29565), .o(n_29677) );
in01f80 g773936 ( .a(n_7050), .o(n_7051) );
in01f80 g776206 ( .a(n_4530), .o(n_4531) );
no02f80 g741944 ( .a(n_38121), .b(n_38059), .o(n_38141) );
in01f80 g779684 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_1_), .o(n_1365) );
na02f80 g752182 ( .a(n_27941), .b(n_27896), .o(n_27975) );
in01f80 g757676 ( .a(n_22819), .o(n_22792) );
ao12f80 g777838 ( .a(n_2964), .b(n_3176), .c(n_2999), .o(n_3232) );
na02f80 g770564 ( .a(n_10278), .b(n_9188), .o(n_10396) );
in01f80 newInst_299 ( .a(newNet_298), .o(newNet_299) );
na02f80 g745377 ( .a(FE_OCP_RBN2987_n_35539), .b(n_35884), .o(n_35962) );
na02f80 g769593 ( .a(n_11381), .b(n_11380), .o(n_11425) );
na02f80 g753103 ( .a(n_27303), .b(n_27302), .o(n_27304) );
in01f80 g744825 ( .a(n_35102), .o(n_35101) );
na02f80 g772800 ( .a(n_8089), .b(n_47236), .o(n_8109) );
in01f80 g765262 ( .a(n_15671), .o(n_15672) );
in01f80 newInst_1726 ( .a(newNet_1725), .o(newNet_1726) );
na02f80 g749205 ( .a(n_30825), .b(n_30845), .o(n_30930) );
in01f80 g765567 ( .a(n_15293), .o(n_15373) );
oa12f80 g774254 ( .a(n_6676), .b(n_6862), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n_6818) );
in01f80 g766542 ( .a(n_14121), .o(n_14091) );
no02f80 g755810 ( .a(n_24359), .b(FE_OCP_RBN2306_n_24288), .o(n_24397) );
in01f80 newInst_2027 ( .a(newNet_1619), .o(newNet_2027) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_18_ ( .ck(newNet_1755), .d(n_22361), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_) );
no02f80 g762395 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18488), .o(n_18524) );
in01f80 newInst_3735 ( .a(newNet_3734), .o(newNet_3735) );
oa22f80 FE_RC_111_0 ( .a(n_19738), .b(n_19920), .c(n_19737), .d(n_19890), .o(n_20020) );
in01f80 g767827 ( .a(n_12967), .o(n_13138) );
in01f80 g756555 ( .a(n_23736), .o(n_23768) );
in01f80 g747365 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .o(n_32624) );
na02f80 g746886 ( .a(FE_OCP_RBN3387_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_28_), .o(n_33326) );
in01f80 newInst_2000 ( .a(newNet_1999), .o(newNet_2000) );
in01f80 g740274 ( .a(n_40210), .o(n_40211) );
na02f80 g769953 ( .a(n_11071), .b(n_11126), .o(n_11212) );
na02f80 g761320 ( .a(n_19850), .b(n_19849), .o(n_19851) );
in01f80 FE_OCP_RBC3039_n_46337 ( .a(n_46337), .o(FE_OCP_RBN3039_n_46337) );
in01f80 newInst_2333 ( .a(newNet_2332), .o(newNet_2333) );
no02f80 g742840 ( .a(n_37188), .b(n_37081), .o(n_37215) );
in01f80 newInst_1340 ( .a(newNet_960), .o(newNet_1340) );
in01f80 g752846 ( .a(n_27076), .o(n_27077) );
in01f80 g756139 ( .a(FE_OCP_RBN2525_n_24902), .o(n_24981) );
ao12f80 g741796 ( .a(n_38398), .b(n_38397), .c(n_38396), .o(n_38872) );
in01f80 g741465 ( .a(n_38770), .o(n_38763) );
in01f80 fopt782908 ( .a(n_44356), .o(n_44355) );
in01f80 g756341 ( .a(n_24018), .o(n_24019) );
in01f80 g758372 ( .a(n_22185), .o(n_22186) );
in01f80 g757604 ( .a(n_22889), .o(n_22890) );
na02f80 g754318 ( .a(n_25907), .b(FE_OCPN1522_n_26054), .o(n_25924) );
no02f80 g775766 ( .a(n_5420), .b(n_5050), .o(n_5539) );
na02f80 g780518 ( .a(n_986), .b(n_1053), .o(n_1070) );
in01f80 g765302 ( .a(n_15871), .o(n_15872) );
in01f80 g768629 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_), .o(n_12229) );
no03m80 FE_RC_2183_0 ( .a(n_22292), .b(n_22383), .c(n_22291), .o(FE_RN_780_0) );
na02f80 g773199 ( .a(n_7730), .b(n_7715), .o(n_7805) );
na02f80 g771140 ( .a(n_9789), .b(n_8240), .o(n_9999) );
in01f80 g744724 ( .a(n_35253), .o(n_35229) );
na02f80 g778267 ( .a(n_2921), .b(n_2975), .o(n_3014) );
in01f80 g775243 ( .a(n_5957), .o(n_5958) );
in01f80 newInst_938 ( .a(newNet_937), .o(newNet_938) );
in01f80 g749584 ( .a(n_31692), .o(n_31693) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_9_ ( .ck(newNet_3465), .d(n_21851), .o(delay_add_ln22_unr14_stage6_stallmux_q_9_) );
ao12f80 g772990 ( .a(n_7312), .b(n_7745), .c(n_7325), .o(n_7810) );
in01f80 newInst_2 ( .a(newNet_1), .o(newNet_2) );
in01f80 g744974 ( .a(n_36403), .o(n_36404) );
in01f80 newInst_3615 ( .a(newNet_513), .o(newNet_3615) );
in01f80 g748311 ( .a(n_31802), .o(n_31803) );
in01f80 g759297 ( .a(n_21261), .o(n_21262) );
in01f80 FE_RC_1840_0 ( .a(n_23074), .o(FE_RN_557_0) );
in01f80 FE_OCP_RBC1336_n_20941 ( .a(n_20941), .o(FE_OCP_RBN1336_n_20941) );
oa12f80 g762294 ( .a(n_18060), .b(n_18008), .c(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_18176) );
na02f80 g746987 ( .a(n_32857), .b(n_32347), .o(n_32934) );
in01f80 g754767 ( .a(n_26856), .o(n_26896) );
in01f80 FE_OCP_RBC2956_n_26231 ( .a(FE_OCP_RBN2955_n_26231), .o(FE_OCP_RBN2956_n_26231) );
ao12f80 g767424 ( .a(n_13475), .b(n_13474), .c(n_13473), .o(n_13934) );
na02f80 FE_RC_1108_0 ( .a(FE_RN_330_0), .b(FE_RN_331_0), .o(FE_RN_332_0) );
na02f80 g766029 ( .a(n_14716), .b(n_13563), .o(n_14718) );
in01f80 g756041 ( .a(n_25053), .o(n_25054) );
na02f80 g740570 ( .a(n_45740), .b(n_39678), .o(n_39697) );
na02f80 g781138 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_5_), .o(n_221) );
no02f80 g774490 ( .a(n_6556), .b(n_6061), .o(n_6862) );
na02f80 g755581 ( .a(n_24612), .b(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24644) );
in01f80 g749857 ( .a(n_31289), .o(n_31219) );
na02f80 g762740 ( .a(n_17892), .b(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_17946) );
ao12f80 g753922 ( .a(n_26215), .b(n_26267), .c(n_26214), .o(n_26370) );
na02f80 g770079 ( .a(n_10940), .b(n_10953), .o(n_10986) );
in01f80 FE_RC_2711_0 ( .a(n_12945), .o(FE_RN_1142_0) );
ao12f80 g746457 ( .a(n_33345), .b(n_33344), .c(n_33343), .o(n_34118) );
na02f80 g738088 ( .a(n_42072), .b(n_42013), .o(n_42073) );
in01f80 newInst_1173 ( .a(newNet_1172), .o(newNet_1173) );
in01f80 newInst_1091 ( .a(newNet_1090), .o(newNet_1091) );
no02f80 g757811 ( .a(n_23121), .b(n_23120), .o(n_23185) );
in01f80 g742730 ( .a(n_37912), .o(n_37495) );
in01f80 g748514 ( .a(n_31678), .o(n_31700) );
na02f80 g736620 ( .a(n_43442), .b(n_43320), .o(n_43444) );
na02f80 g738191 ( .a(n_41985), .b(n_41792), .o(n_41999) );
in01f80 g753488 ( .a(n_26875), .o(n_26876) );
ao12f80 g738041 ( .a(n_41687), .b(n_42145), .c(n_41602), .o(n_42163) );
no02f80 g747118 ( .a(n_32870), .b(n_32717), .o(n_32890) );
no02f80 g772845 ( .a(n_7821), .b(n_7378), .o(n_7869) );
no02f80 g779213 ( .a(n_1862), .b(n_1632), .o(n_1864) );
no02f80 g749929 ( .a(n_30195), .b(n_30050), .o(n_30197) );
in01f80 FE_OCP_RBC2215_FE_OCPN950_n_28595 ( .a(FE_OCP_RBN2214_FE_OCPN950_n_28595), .o(FE_OCP_RBN2215_FE_OCPN950_n_28595) );
na02f80 g775301 ( .a(n_5806), .b(n_5607), .o(n_5866) );
oa22f80 g752495 ( .a(n_27653), .b(n_24350), .c(n_27635), .d(n_27796), .o(n_27687) );
in01f80 g777346 ( .a(n_4702), .o(n_4773) );
na02f80 g748188 ( .a(FE_OCP_RBN3712_n_31466), .b(n_31558), .o(n_31666) );
in01f80 newInst_231 ( .a(newNet_230), .o(newNet_231) );
in01f80 newInst_361 ( .a(newNet_217), .o(newNet_361) );
in01f80 newInst_2439 ( .a(newNet_1459), .o(newNet_2439) );
na02f80 g736721 ( .a(n_43140), .b(n_43230), .o(n_43231) );
no02f80 g766416 ( .a(n_14002), .b(n_13958), .o(n_14071) );
na02f80 g768044 ( .a(n_12721), .b(n_12289), .o(n_12775) );
na02f80 g781331 ( .a(n_1), .b(beta_7), .o(n_58) );
in01f80 g767706 ( .a(n_13028), .o(n_13029) );
no02f80 g751857 ( .a(n_28209), .b(n_28218), .o(n_28299) );
oa12f80 g780263 ( .a(n_766), .b(n_786), .c(n_765), .o(n_791) );
in01f80 g751324 ( .a(n_29598), .o(n_29599) );
in01f80 g760100 ( .a(n_20533), .o(n_20575) );
na02f80 g769932 ( .a(n_11022), .b(n_11014), .o(n_11075) );
na02f80 g751057 ( .a(n_29909), .b(n_30165), .o(n_30061) );
no02f80 g744965 ( .a(n_34976), .b(n_34992), .o(n_35075) );
in01f80 g775815 ( .a(n_5304), .o(n_5305) );
no02f80 g760922 ( .a(n_19360), .b(n_19218), .o(n_19438) );
oa12f80 g738881 ( .a(n_41047), .b(n_41194), .c(n_41229), .o(n_41258) );
in01f80 g771854 ( .a(n_10159), .o(n_10119) );
ao22s80 g736423 ( .a(n_43744), .b(n_43354), .c(n_43745), .d(n_43353), .o(n_43785) );
in01f80 g752447 ( .a(n_27720), .o(n_27698) );
in01f80 g760652 ( .a(n_19833), .o(n_19834) );
na02f80 g737081 ( .a(n_43103), .b(n_42781), .o(n_43199) );
na02f80 g765135 ( .a(n_15204), .b(n_14215), .o(n_15237) );
no02f80 g761879 ( .a(n_18595), .b(n_18549), .o(n_18639) );
no02f80 g751801 ( .a(n_29131), .b(n_29101), .o(n_29203) );
in01f80 g743316 ( .a(n_36787), .o(n_36788) );
oa22f80 FE_RC_784_0 ( .a(n_40598), .b(FE_OCP_RBN3138_n_40568), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_40568), .o(n_40580) );
na02f80 g767986 ( .a(n_12884), .b(n_13078), .o(n_13504) );
in01f80 newInst_129 ( .a(newNet_128), .o(newNet_129) );
in01f80 g768605 ( .a(n_12334), .o(n_12291) );
in01f80 g756724 ( .a(n_24107), .o(n_24047) );
in01f80 g746039 ( .a(n_33977), .o(n_34033) );
oa22f80 g761956 ( .a(n_18203), .b(n_18149), .c(n_18248), .d(n_18150), .o(n_18287) );
na02f80 g753681 ( .a(n_26560), .b(n_26764), .o(n_26647) );
no02f80 g778468 ( .a(n_2628), .b(delay_add_ln22_unr2_stage2_stallmux_q_25_), .o(n_2734) );
in01f80 g741408 ( .a(n_38804), .o(n_38805) );
oa12f80 g778085 ( .a(n_2775), .b(n_2938), .c(n_2739), .o(n_2980) );
na02f80 g771202 ( .a(n_9057), .b(n_8232), .o(n_9144) );
no02f80 g756939 ( .a(n_24007), .b(n_24074), .o(n_24664) );
no02f80 g776585 ( .a(n_4051), .b(n_4032), .o(n_4125) );
na02f80 g770253 ( .a(n_10666), .b(n_10647), .o(n_10754) );
na02f80 FE_RC_4042_0 ( .a(FE_OCP_RBN2629_n_14590), .b(n_16319), .o(FE_RN_1756_0) );
na02f80 g751864 ( .a(n_28188), .b(delay_add_ln22_unr17_stage7_stallmux_q_6_), .o(n_28250) );
no03m80 g751820 ( .a(n_29129), .b(n_29046), .c(n_29071), .o(n_29130) );
na02f80 g750649 ( .a(n_29440), .b(FE_OCPN3747_n_29439), .o(n_29516) );
in01f80 g772809 ( .a(n_8224), .o(n_8121) );
no02f80 g759644 ( .a(FE_OCP_RBN1707_n_20616), .b(n_20337), .o(n_20643) );
in01f80 newInst_674 ( .a(newNet_455), .o(newNet_674) );
no02f80 g773159 ( .a(n_7743), .b(n_7812), .o(n_7996) );
no02f80 g753648 ( .a(n_26538), .b(n_23564), .o(n_26985) );
in01f80 FE_OCP_RBC2263_n_29033 ( .a(n_29033), .o(FE_OCP_RBN2263_n_29033) );
oa22f80 g778509 ( .a(n_2296), .b(n_2360), .c(n_2295), .d(n_2359), .o(n_3721) );
ao12f80 g749978 ( .a(n_30161), .b(n_30925), .c(n_30062), .o(n_30976) );
na02f80 g738715 ( .a(n_41378), .b(n_41402), .o(n_41419) );
no02f80 g771950 ( .a(n_44463), .b(n_9681), .o(n_9771) );
in01f80 newInst_551 ( .a(newNet_550), .o(newNet_551) );
na02f80 g770547 ( .a(n_10337), .b(n_10279), .o(n_10467) );
in01f80 g776960 ( .a(n_3633), .o(n_3681) );
in01f80 g770694 ( .a(n_10417), .o(n_10418) );
oa22f80 g770722 ( .a(FE_OCP_RBN3653_n_10100), .b(n_9197), .c(FE_OCP_RBN2775_n_10100), .d(n_9114), .o(n_10456) );
na02f80 g765358 ( .a(n_15224), .b(n_15223), .o(n_15256) );
no02f80 g773837 ( .a(n_7118), .b(n_6951), .o(n_7153) );
no02f80 g770164 ( .a(n_10862), .b(n_10608), .o(n_10863) );
na02f80 g752039 ( .a(n_28143), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .o(n_28222) );
no02f80 g767669 ( .a(n_13371), .b(n_13356), .o(n_13391) );
in01f80 newInst_3439 ( .a(newNet_3438), .o(newNet_3439) );
na02f80 g775294 ( .a(n_5894), .b(n_5005), .o(n_5944) );
in01f80 FE_OCPC1251_n_8210 ( .a(FE_OCP_RBN3500_n_8187), .o(FE_OCPN1251_n_8210) );
no02f80 g780594 ( .a(n_745), .b(n_773), .o(n_793) );
in01f80 g757655 ( .a(n_22674), .o(n_23035) );
na02f80 g778243 ( .a(n_2697), .b(n_2393), .o(n_2772) );
in01f80 g774181 ( .a(n_6639), .o(n_6640) );
na02f80 g749202 ( .a(n_30739), .b(n_45489), .o(n_30773) );
in01f80 FE_OCP_RBC3665_n_4604 ( .a(n_4604), .o(FE_OCP_RBN3665_n_4604) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_6_ ( .ck(newNet_434), .d(n_27797), .o(delay_xor_ln22_unr18_stage7_stallmux_q_6_) );
na02f80 g781046 ( .a(cos_out_6), .b(FE_OFN2_n_43918), .o(n_319) );
no02f80 g749762 ( .a(n_31118), .b(n_31067), .o(n_31174) );
ao12f80 g761169 ( .a(n_19768), .b(n_19769), .c(n_19767), .o(n_21105) );
no02f80 FE_RC_2596_0 ( .a(FE_RN_1074_0), .b(n_2937), .o(FE_RN_1075_0) );
ao12f80 g739226 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_15_), .b(n_45146), .c(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n_40679) );
in01f80 newInst_506 ( .a(newNet_505), .o(newNet_506) );
no02f80 FE_RC_4162_0 ( .a(n_33181), .b(n_33186), .o(FE_RN_1813_0) );
no03m80 FE_RC_685_0 ( .a(n_40825), .b(n_40826), .c(n_40725), .o(n_40866) );
na02f80 g744789 ( .a(n_35099), .b(n_30633), .o(n_35148) );
na02f80 g766283 ( .a(n_14202), .b(n_14203), .o(n_14334) );
no02f80 g756514 ( .a(n_23679), .b(n_23607), .o(n_23714) );
in01f80 g766838 ( .a(n_13645), .o(n_13664) );
na02f80 g762043 ( .a(n_18930), .b(n_18807), .o(n_18934) );
na02f80 FE_RC_1846_0 ( .a(FE_RN_561_0), .b(n_36108), .o(FE_RN_562_0) );
in01f80 newInst_2592 ( .a(newNet_2591), .o(newNet_2592) );
no02f80 g742432 ( .a(n_37774), .b(n_37752), .o(n_38698) );
na02f80 FE_RC_3506_0 ( .a(n_29110), .b(FE_RN_1514_0), .o(n_29154) );
na02f80 g750618 ( .a(n_29380), .b(n_29239), .o(n_29381) );
no02f80 g768887 ( .a(n_11847), .b(n_11723), .o(n_11848) );
in01f80 g774264 ( .a(n_6670), .o(n_6646) );
in01f80 g761384 ( .a(n_18980), .o(n_19082) );
no02f80 g759669 ( .a(n_20638), .b(n_20682), .o(n_20761) );
oa12f80 g747264 ( .a(n_33887), .b(n_45753), .c(n_33885), .o(n_34497) );
in01f80 FE_OCP_RBC3491_n_29553 ( .a(n_29553), .o(FE_OCP_RBN3491_n_29553) );
no02f80 FE_RC_3354_0 ( .a(FE_RN_1463_0), .b(FE_RN_1325_0), .o(n_21218) );
ao12f80 g755192 ( .a(n_24978), .b(n_24977), .c(n_24976), .o(n_26626) );
in01f80 FE_OCP_RBC2455_n_14157 ( .a(n_14157), .o(FE_OCP_RBN2455_n_14157) );
no02f80 g736661 ( .a(n_43329), .b(n_43370), .o(n_43371) );
no02f80 FE_RC_1517_0 ( .a(n_31716), .b(n_32223), .o(FE_RN_427_0) );
in01f80 newInst_962 ( .a(newNet_961), .o(newNet_962) );
ao22s80 FE_RC_1293_0 ( .a(n_8934), .b(n_8899), .c(n_8891), .d(n_8898), .o(n_9075) );
in01f80 newInst_3753 ( .a(newNet_3752), .o(newNet_3753) );
in01f80 newInst_401 ( .a(newNet_400), .o(newNet_401) );
in01f80 g750710 ( .a(n_29477), .o(n_30111) );
na02f80 g744003 ( .a(n_36198), .b(n_36191), .o(n_36301) );
ao22s80 FE_RC_2974_0 ( .a(n_14741), .b(n_14790), .c(n_14791), .d(n_14720), .o(n_14905) );
in01f80 g773713 ( .a(n_7311), .o(n_7896) );
in01f80 g775600 ( .a(n_5663), .o(n_5695) );
in01f80 g775063 ( .a(n_6146), .o(n_6137) );
na02f80 g774454 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n_6849) );
no02f80 g742675 ( .a(n_37486), .b(n_37485), .o(n_37487) );
in01f80 newInst_1782 ( .a(newNet_1781), .o(newNet_1782) );
no02f80 g768286 ( .a(n_12644), .b(n_12642), .o(n_12643) );
in01f80 g763903 ( .a(n_17104), .o(n_17055) );
oa12f80 g741830 ( .a(n_38118), .b(n_38386), .c(n_38082), .o(n_38389) );
in01f80 newInst_635 ( .a(newNet_51), .o(newNet_635) );
in01f80 FE_OCP_RBC3425_n_44881 ( .a(n_44881), .o(FE_OCP_RBN3425_n_44881) );
ao22s80 FE_RC_3415_0 ( .a(FE_OCP_RBN1131_n_24179), .b(n_24312), .c(FE_OCP_RBN1130_n_24179), .d(n_24311), .o(n_24503) );
na02f80 g781036 ( .a(sin_out_13), .b(FE_OFN3_n_43918), .o(n_300) );
in01f80 g768496 ( .a(n_12408), .o(n_12409) );
no02f80 g761276 ( .a(n_20011), .b(n_19980), .o(n_20050) );
no02f80 g738921 ( .a(n_41224), .b(n_40984), .o(n_41265) );
na02f80 g755521 ( .a(n_25468), .b(n_25467), .o(n_25469) );
oa12f80 g755080 ( .a(n_25718), .b(n_25717), .c(n_25716), .o(n_26510) );
in01f80 g758129 ( .a(n_23152), .o(n_23153) );
in01f80 g765904 ( .a(n_14891), .o(n_14824) );
na02f80 g745625 ( .a(n_34369), .b(FE_OCP_RBN1353_n_33584), .o(n_34454) );
na02f80 g774519 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .o(n_6782) );
in01f80 g761805 ( .a(n_18564), .o(n_18517) );
ao12f80 g739477 ( .a(n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n_40826) );
no02f80 g740651 ( .a(n_39586), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39604) );
ao12f80 g780733 ( .a(n_603), .b(n_608), .c(n_602), .o(n_808) );
no02f80 g745582 ( .a(n_34291), .b(n_34293), .o(n_34318) );
in01f80 g763661 ( .a(n_16893), .o(n_16894) );
na02f80 g762926 ( .a(n_17763), .b(n_15892), .o(n_17864) );
no02f80 g763322 ( .a(n_17179), .b(n_17216), .o(n_17384) );
in01f80 FE_OCPC869_n_16086 ( .a(FE_OCPN868_n_16086), .o(FE_OCPN869_n_16086) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_19_ ( .ck(newNet_1524), .d(n_32257), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_) );
no03m80 g777857 ( .a(n_2706), .b(n_3212), .c(n_2661), .o(n_3213) );
na02f80 g751784 ( .a(n_28291), .b(n_28290), .o(n_28292) );
oa22f80 FE_RC_1226_0 ( .a(n_6465), .b(n_6576), .c(n_6466), .d(n_47335), .o(n_6774) );
no02f80 g780792 ( .a(n_412), .b(n_1108), .o(n_413) );
in01f80 g775997 ( .a(n_5085), .o(n_5086) );
oa22f80 FE_RC_1393_0 ( .a(n_16554), .b(n_16489), .c(n_16553), .d(n_16514), .o(n_16638) );
in01f80 g749629 ( .a(n_31740), .o(n_30284) );
na02f80 g769873 ( .a(n_11072), .b(n_11035), .o(n_11110) );
in01f80 g758612 ( .a(n_21922), .o(n_21937) );
no02f80 g771586 ( .a(n_8983), .b(n_9012), .o(n_9013) );
oa12f80 g752530 ( .a(n_27256), .b(n_27602), .c(n_27601), .o(n_27610) );
oa12f80 g746424 ( .a(n_33469), .b(n_33468), .c(n_33467), .o(n_34127) );
in01f80 g770667 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .o(n_10419) );
in01f80 g749184 ( .a(n_30776), .o(n_30777) );
in01f80 FE_OCP_RBC2975_n_5531 ( .a(FE_OCP_RBN2974_n_5531), .o(FE_OCP_RBN2975_n_5531) );
in01f80 newInst_1556 ( .a(newNet_157), .o(newNet_1556) );
in01f80 g771330 ( .a(n_9090), .o(n_9111) );
no02f80 g770705 ( .a(n_10290), .b(n_10768), .o(n_10390) );
oa12f80 g780806 ( .a(n_363), .b(n_379), .c(n_371), .o(n_386) );
no02f80 g779627 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .o(n_1913) );
na02f80 g766166 ( .a(n_14839), .b(n_14838), .o(n_14840) );
oa12f80 g758779 ( .a(n_22178), .b(n_22177), .c(n_22176), .o(n_22245) );
no02f80 g779561 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_17_), .o(n_1881) );
in01f80 newInst_51 ( .a(newNet_50), .o(newNet_51) );
na02f80 g756428 ( .a(n_23615), .b(n_23587), .o(n_23588) );
in01f80 g759159 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_4_), .o(n_21457) );
oa12f80 g741090 ( .a(n_38804), .b(n_38856), .c(n_38816), .o(n_38968) );
na02f80 FE_RC_2374_0 ( .a(FE_RN_922_0), .b(n_42600), .o(n_42652) );
no02f80 g765117 ( .a(n_15142), .b(n_15456), .o(n_15525) );
na02f80 g758102 ( .a(FE_OCPN979_n_21973), .b(FE_OCP_RBN1845_n_20910), .o(n_22047) );
no02f80 FE_RC_2157_0 ( .a(n_14420), .b(n_15314), .o(FE_RN_763_0) );
in01f80 g776614 ( .a(n_4252), .o(n_4253) );
in01f80 g771850 ( .a(n_10120), .o(n_10121) );
na02f80 g755681 ( .a(n_25063), .b(n_25092), .o(n_25093) );
in01f80 FE_OCPC963_n_27287 ( .a(n_27287), .o(FE_OCPN963_n_27287) );
in01f80 g757932 ( .a(n_22470), .o(n_22471) );
in01f80 g747318 ( .a(FE_OCPN1236_n_32791), .o(n_32553) );
ao22s80 FE_RC_3732_0 ( .a(n_44711), .b(n_6439), .c(n_6438), .d(n_44710), .o(n_6567) );
in01f80 newInst_3406 ( .a(newNet_3405), .o(newNet_3406) );
no02f80 g769355 ( .a(n_10419), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11727) );
oa12f80 g758872 ( .a(n_22062), .b(n_22061), .c(n_22060), .o(n_22118) );
in01f80 g745000 ( .a(n_34836), .o(n_35824) );
na02f80 g740923 ( .a(n_39087), .b(n_39276), .o(n_39308) );
in01f80 g737615 ( .a(n_42251), .o(n_42252) );
in01f80 fopt783261 ( .a(n_7659), .o(n_44829) );
in01f80 newInst_3053 ( .a(newNet_3052), .o(newNet_3053) );
in01f80 FE_OFC824_n_3500 ( .a(FE_OFN840_n_3500), .o(FE_OFN824_n_3500) );
ao12f80 g747700 ( .a(n_33392), .b(n_33532), .c(n_33227), .o(n_33603) );
no02f80 g740938 ( .a(n_39213), .b(n_39063), .o(n_39286) );
no02f80 g762680 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_24_), .b(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n_17813) );
no02f80 g751277 ( .a(n_29744), .b(n_29204), .o(n_29745) );
in01f80 newInst_2189 ( .a(newNet_2031), .o(newNet_2189) );
na02f80 g746261 ( .a(n_33674), .b(n_33232), .o(n_33707) );
na02f80 g778665 ( .a(n_2256), .b(n_2250), .o(n_2325) );
in01f80 g746776 ( .a(n_34739), .o(n_34155) );
in01f80 g742728 ( .a(n_37518), .o(n_37545) );
in01f80 FE_OCPC1523_n_45072 ( .a(n_45072), .o(FE_OCPN1523_n_45072) );
oa12f80 g752120 ( .a(n_28639), .b(n_28638), .c(n_28637), .o(n_28899) );
no02f80 g770223 ( .a(n_10696), .b(n_10667), .o(n_10759) );
oa22f80 FE_RC_392_0 ( .a(n_13152), .b(n_12715), .c(n_12714), .d(n_13151), .o(n_13334) );
in01f80 g755727 ( .a(n_25063), .o(n_25438) );
na04m80 g751374 ( .a(n_28722), .b(n_28650), .c(n_28770), .d(n_28720), .o(n_28788) );
na02f80 g778229 ( .a(n_2689), .b(n_2688), .o(n_2690) );
oa12f80 g764946 ( .a(n_16351), .b(n_16350), .c(n_16349), .o(n_16411) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_14_ ( .ck(newNet_3165), .d(n_40458), .o(delay_add_ln22_unr27_stage10_stallmux_q_14_) );
oa22f80 g776271 ( .a(n_4376), .b(FE_OCP_RBN2691_FE_OCPN843_n_3912), .c(FE_OCP_RBN2766_n_4376), .d(FE_OCPN960_n_3951), .o(n_4554) );
in01f80 newInst_3558 ( .a(newNet_3452), .o(newNet_3558) );
no02f80 g780064 ( .a(n_1223), .b(n_885), .o(n_1230) );
in01f80 fopt783928 ( .a(n_24506), .o(n_45635) );
na02f80 g743649 ( .a(n_36352), .b(n_35954), .o(n_36382) );
na02f80 g742861 ( .a(n_37128), .b(n_37008), .o(n_37214) );
in01f80 g751598 ( .a(n_28698), .o(n_28735) );
in01f80 g750219 ( .a(n_29809), .o(n_29846) );
na02f80 FE_RC_2098_0 ( .a(FE_RN_721_0), .b(n_14873), .o(FE_RN_722_0) );
no02f80 g772590 ( .a(n_8337), .b(n_7892), .o(n_8369) );
no02f80 g773105 ( .a(n_7980), .b(n_7964), .o(n_8706) );
na02f80 g766659 ( .a(n_13887), .b(n_13886), .o(n_13931) );
na02f80 g777873 ( .a(n_3185), .b(n_3243), .o(n_3244) );
na02f80 g737373 ( .a(n_42806), .b(n_42625), .o(n_42837) );
in01f80 g778474 ( .a(n_2681), .o(n_2682) );
oa22f80 FE_RC_3328_0 ( .a(n_33404), .b(n_33875), .c(n_33900), .d(n_33405), .o(n_33976) );
ao22s80 FE_RC_4005_0 ( .a(n_34703), .b(n_35026), .c(n_34702), .d(n_35048), .o(n_35132) );
ao12f80 g779430 ( .a(n_1595), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_9_), .o(n_1842) );
in01f80 g780773 ( .a(FE_OCPN1408_n_672), .o(n_556) );
in01f80 g740079 ( .a(n_40328), .o(n_40329) );
in01f80 g773641 ( .a(n_7378), .o(n_7379) );
in01f80 FE_OCPC3183_n_22294 ( .a(n_22294), .o(FE_OCPN3183_n_22294) );
no02f80 g782645 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_19_), .b(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n_44039) );
oa12f80 g784644 ( .a(n_16840), .b(n_16811), .c(n_16785), .o(n_46974) );
in01f80 FE_OCP_RBC2790_n_4462 ( .a(n_4462), .o(FE_OCP_RBN2790_n_4462) );
in01f80 newInst_3642 ( .a(newNet_3641), .o(newNet_3642) );
na02f80 g779275 ( .a(n_1727), .b(n_912), .o(n_1814) );
no02f80 g745062 ( .a(n_34788), .b(n_34563), .o(n_34826) );
in01f80 g746129 ( .a(n_33778), .o(n_33779) );
na02f80 g759901 ( .a(n_21374), .b(n_21373), .o(n_21478) );
na02f80 g737520 ( .a(n_42532), .b(n_42403), .o(n_42455) );
na02f80 g777897 ( .a(n_3164), .b(n_3148), .o(n_4022) );
ao12f80 g768819 ( .a(n_11872), .b(n_12005), .c(n_11875), .o(n_12176) );
in01f80 g767486 ( .a(n_13228), .o(n_13245) );
ao12f80 g759072 ( .a(n_20661), .b(n_21143), .c(n_20786), .o(n_21197) );
na02f80 g770246 ( .a(n_10569), .b(n_10592), .o(n_10620) );
no02f80 g738987 ( .a(n_41147), .b(n_41146), .o(n_41148) );
in01f80 g767545 ( .a(n_13324), .o(n_13325) );
na02f80 g777252 ( .a(n_3565), .b(n_3581), .o(n_3666) );
no02f80 g748078 ( .a(n_31746), .b(n_31735), .o(n_31747) );
no02f80 g774864 ( .a(n_6176), .b(FE_OCP_RBN3696_n_5284), .o(n_6240) );
no02f80 g766801 ( .a(n_13703), .b(n_13702), .o(n_13713) );
na02f80 g760160 ( .a(n_20299), .b(FE_OCP_RBN1692_n_19052), .o(n_20413) );
na02f80 FE_RC_1278_0 ( .a(FE_RN_375_0), .b(FE_RN_376_0), .o(FE_RN_377_0) );
in01f80 newInst_2289 ( .a(newNet_751), .o(newNet_2289) );
in01f80 g755132 ( .a(n_25535), .o(n_25499) );
na02f80 g740216 ( .a(n_39892), .b(n_39942), .o(n_40003) );
in01f80 newInst_2063 ( .a(newNet_2062), .o(newNet_2063) );
no02f80 g766438 ( .a(n_14100), .b(n_13240), .o(n_14123) );
in01f80 g777738 ( .a(n_3343), .o(n_3344) );
na02f80 g767930 ( .a(n_12817), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .o(n_12954) );
oa22f80 FE_RC_1489_0 ( .a(n_24059), .b(n_27727), .c(n_27796), .d(n_27705), .o(n_27749) );
oa22f80 g780348 ( .a(n_921), .b(n_840), .c(n_920), .d(n_919), .o(n_990) );
in01f80 g777900 ( .a(n_3259), .o(n_3260) );
in01f80 g777078 ( .a(n_4070), .o(n_4049) );
in01f80 g756707 ( .a(n_23579), .o(n_23544) );
in01f80 FE_RC_2727_0 ( .a(n_18339), .o(FE_RN_1154_0) );
oa22f80 g780536 ( .a(n_923), .b(n_893), .c(n_890), .d(n_640), .o(n_1059) );
no02f80 g753436 ( .a(n_27589), .b(n_26817), .o(n_27613) );
ms00f80 cos_out_reg_26_ ( .ck(newNet_3708), .d(n_43891), .o(cos_out_26) );
na02f80 g754896 ( .a(FE_OCP_RBN2594_n_25181), .b(FE_OCP_RBN2278_n_24173), .o(n_25276) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_28_ ( .ck(newNet_3207), .d(n_36608), .o(delay_add_ln22_unr23_stage9_stallmux_q_28_) );
no02f80 g744931 ( .a(n_34972), .b(n_34654), .o(n_35049) );
na02f80 g777637 ( .a(n_3433), .b(n_3473), .o(n_3548) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_29_ ( .ck(newNet_2454), .d(n_32518), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_) );
no02f80 g776059 ( .a(n_5059), .b(n_5058), .o(n_5060) );
na02f80 g741780 ( .a(n_38423), .b(n_38422), .o(n_38424) );
na02f80 g774538 ( .a(n_6416), .b(n_6387), .o(n_6491) );
in01f80 g762344 ( .a(n_18726), .o(n_18727) );
in01f80 g777759 ( .a(n_5062), .o(n_3323) );
no02f80 g765213 ( .a(n_15338), .b(n_15337), .o(n_15457) );
no02f80 g779002 ( .a(n_2161), .b(delay_add_ln22_unr2_stage2_stallmux_q_17_), .o(n_2181) );
ao12f80 g738180 ( .a(n_42010), .b(n_42009), .c(n_42008), .o(n_42066) );
na02f80 g776340 ( .a(n_4541), .b(n_4540), .o(n_4629) );
no02f80 g775503 ( .a(n_5759), .b(FE_OCP_RBN2817_n_4458), .o(n_5812) );
in01f80 newInst_1628 ( .a(newNet_1627), .o(newNet_1628) );
no02f80 g760811 ( .a(n_19479), .b(n_19478), .o(n_19480) );
na02f80 FE_RC_2060_0 ( .a(n_26620), .b(n_26664), .o(FE_RN_698_0) );
no02f80 g776779 ( .a(n_4127), .b(n_3910), .o(n_4257) );
in01f80 newInst_1497 ( .a(newNet_1454), .o(newNet_1497) );
in01f80 FE_OCP_RBC2560_n_3437 ( .a(n_3437), .o(FE_OCP_RBN2560_n_3437) );
in01f80 FE_OCP_RBC2741_n_15206 ( .a(n_15206), .o(FE_OCP_RBN2741_n_15206) );
in01f80 newInst_2771 ( .a(newNet_2770), .o(newNet_2771) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_25_ ( .ck(newNet_2736), .d(n_17686), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_) );
in01f80 g775005 ( .a(n_6148), .o(n_6173) );
no02f80 g736712 ( .a(n_43180), .b(n_43082), .o(n_43370) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_26_ ( .ck(newNet_1304), .d(n_1272), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_) );
in01f80 FE_OCP_RBC2839_n_4692 ( .a(FE_OCP_RBN2838_n_4692), .o(FE_OCP_RBN2839_n_4692) );
in01f80 g754521 ( .a(n_26611), .o(n_26612) );
no02f80 g738143 ( .a(n_42066), .b(n_42065), .o(n_42067) );
ao22s80 FE_RC_3373_0 ( .a(n_19222), .b(FE_OCP_RBN2260_n_18899), .c(FE_OFN779_n_17093), .d(n_18899), .o(n_19005) );
oa12f80 g774023 ( .a(n_6958), .b(n_6957), .c(n_6956), .o(n_7707) );
in01f80 g766069 ( .a(n_14642), .o(n_14643) );
na02f80 g761701 ( .a(n_18795), .b(n_18748), .o(n_18749) );
no02f80 g763600 ( .a(n_16712), .b(n_16716), .o(n_16717) );
oa12f80 g736288 ( .a(n_307), .b(n_43856), .c(FE_OFN3_n_43918), .o(n_43888) );
in01f80 newInst_642 ( .a(newNet_641), .o(newNet_642) );
in01f80 g762955 ( .a(n_17836), .o(n_17837) );
in01f80 g740119 ( .a(n_40322), .o(n_40323) );
oa12f80 g771731 ( .a(n_9326), .b(n_9325), .c(n_9324), .o(n_9437) );
in01f80 g776890 ( .a(n_3867), .o(n_3740) );
na02f80 g776225 ( .a(n_4831), .b(n_4515), .o(n_4889) );
no02f80 g779053 ( .a(n_2104), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .o(n_2153) );
in01f80 g773749 ( .a(n_7321), .o(n_8135) );
oa22f80 g771552 ( .a(n_9009), .b(FE_OCP_RBN3543_n_44575), .c(FE_OCP_RBN2585_n_9009), .d(n_44563), .o(n_9185) );
oa22f80 FE_RC_3430_0 ( .a(n_26331), .b(n_26400), .c(n_26399), .d(n_26364), .o(n_26522) );
no02f80 g758008 ( .a(n_22264), .b(n_22045), .o(n_22341) );
na02f80 FE_RC_2629_0 ( .a(FE_RN_1094_0), .b(n_12423), .o(n_12492) );
na02f80 g772682 ( .a(n_8236), .b(n_7702), .o(n_8493) );
ao12f80 g737659 ( .a(n_42236), .b(n_42235), .c(n_42234), .o(n_43019) );
na02f80 g745385 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35926), .o(n_36171) );
in01f80 g745148 ( .a(n_34677), .o(n_34678) );
oa12f80 g784440 ( .a(n_46204), .b(n_37992), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_46252) );
na02f80 g751727 ( .a(n_28348), .b(delay_add_ln22_unr17_stage7_stallmux_q_10_), .o(n_28403) );
na02f80 FE_RC_2364_0 ( .a(FE_RN_914_0), .b(n_1741), .o(FE_RN_915_0) );
na02f80 g739663 ( .a(n_40536), .b(n_40250), .o(n_40548) );
in01f80 newInst_1003 ( .a(newNet_696), .o(newNet_1003) );
ao12f80 g746015 ( .a(n_34008), .b(n_34007), .c(n_34006), .o(n_34055) );
ao22s80 g743066 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .c(n_36992), .d(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37571) );
na02f80 g752338 ( .a(n_45200), .b(FE_OCP_RBN3306_n_44722), .o(n_27911) );
no02f80 g747789 ( .a(n_33571), .b(n_33683), .o(n_33970) );
na02f80 FE_RC_2929_0 ( .a(n_27291), .b(FE_RN_1276_0), .o(n_27548) );
no02f80 g772407 ( .a(n_8414), .b(n_8323), .o(n_8521) );
no02f80 g750402 ( .a(n_29632), .b(n_29593), .o(n_29667) );
no02f80 g766454 ( .a(n_14116), .b(n_14089), .o(n_14228) );
oa12f80 g744594 ( .a(n_35350), .b(n_35349), .c(n_35348), .o(n_35378) );
ao22s80 g736376 ( .a(n_43834), .b(n_43463), .c(n_43819), .d(n_43462), .o(n_43878) );
na02f80 g776590 ( .a(n_4383), .b(n_4501), .o(n_4614) );
in01f80 g776152 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_4_), .o(n_4948) );
in01f80 g772422 ( .a(n_44058), .o(n_8542) );
in01f80 newInst_1405 ( .a(newNet_1404), .o(newNet_1405) );
oa22f80 FE_RC_759_0 ( .a(n_11588), .b(n_11652), .c(n_11587), .d(n_11702), .o(n_11873) );
na02f80 g773597 ( .a(n_7427), .b(n_45863), .o(n_7450) );
ao12f80 g770914 ( .a(n_9434), .b(n_10131), .c(n_9505), .o(n_10218) );
oa22f80 FE_RC_1627_0 ( .a(FE_OFN737_n_22641), .b(n_25890), .c(n_23259), .d(n_25891), .o(n_25983) );
in01f80 FE_RC_3776_0 ( .a(FE_RN_1657_0), .o(FE_RN_1656_0) );
in01f80 newInst_480 ( .a(newNet_479), .o(newNet_480) );
oa12f80 g763179 ( .a(n_17474), .b(n_17473), .c(n_17472), .o(n_18860) );
na02f80 g755888 ( .a(n_25407), .b(n_25003), .o(n_25467) );
in01f80 FE_RC_3816_0 ( .a(FE_RN_1239_0), .o(FE_RN_1664_0) );
in01f80 g780638 ( .a(n_865), .o(n_866) );
na02f80 g772603 ( .a(n_8445), .b(n_8444), .o(n_8555) );
oa12f80 g767080 ( .a(n_13611), .b(n_13610), .c(n_13609), .o(n_15462) );
no02f80 g767049 ( .a(FE_OCP_RBN2457_n_13765), .b(n_13289), .o(n_13895) );
in01f80 g763844 ( .a(n_16667), .o(n_16668) );
ao12f80 g772562 ( .a(n_8216), .b(n_8256), .c(n_8182), .o(n_8374) );
in01f80 g769131 ( .a(n_11799), .o(n_11800) );
in01f80 g765127 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_), .o(n_17347) );
ao12f80 g739095 ( .a(n_41018), .b(n_41017), .c(n_41016), .o(n_41447) );
in01f80 newInst_1478 ( .a(newNet_922), .o(newNet_1478) );
na02f80 g775424 ( .a(n_5886), .b(n_5702), .o(n_5887) );
ao12f80 g757940 ( .a(n_22788), .b(n_22737), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_22811) );
in01f80 newInst_599 ( .a(newNet_598), .o(newNet_599) );
no02f80 g776587 ( .a(n_4589), .b(n_4493), .o(n_4708) );
in01f80 newInst_24 ( .a(newNet_23), .o(newNet_24) );
ao22s80 FE_RC_263_0 ( .a(n_21149), .b(n_20658), .c(n_20659), .d(n_21150), .o(n_21312) );
ao12f80 g747696 ( .a(n_33392), .b(n_33513), .c(n_33512), .o(n_33515) );
in01f80 g739998 ( .a(n_40295), .o(n_40333) );
no02f80 g778091 ( .a(n_2884), .b(n_2216), .o(n_2897) );
na02f80 g770756 ( .a(FE_OCP_RBN2775_n_10100), .b(n_9148), .o(n_10304) );
in01f80 g778976 ( .a(n_2216), .o(n_2217) );
no02f80 g748046 ( .a(n_32086), .b(n_31744), .o(n_31879) );
oa12f80 g761291 ( .a(n_19846), .b(n_19983), .c(n_20086), .o(n_21022) );
na02f80 g770048 ( .a(n_10855), .b(n_10457), .o(n_10882) );
in01f80 g751894 ( .a(n_29101), .o(n_29334) );
no02f80 g745620 ( .a(FE_OCP_RBN3433_n_33664), .b(n_34369), .o(n_34564) );
na02f80 g780721 ( .a(n_616), .b(n_484), .o(n_618) );
in01f80 FE_OCP_RBC3457_n_33872 ( .a(FE_OCP_RBN3456_n_33872), .o(FE_OCP_RBN3457_n_33872) );
no02f80 g761151 ( .a(n_19101), .b(n_17900), .o(n_19146) );
in01f80 newInst_3118 ( .a(newNet_3117), .o(newNet_3118) );
in01f80 g750811 ( .a(n_29120), .o(n_29121) );
oa12f80 g780704 ( .a(n_632), .b(n_631), .c(n_630), .o(n_893) );
ao12f80 g763855 ( .a(n_17425), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .o(n_17986) );
no02f80 g751261 ( .a(n_29745), .b(n_29248), .o(n_29800) );
in01f80 g748142 ( .a(n_31990), .o(n_31991) );
in01f80 g766855 ( .a(n_13742), .o(n_15643) );
no02f80 g778603 ( .a(n_2652), .b(n_2612), .o(n_2655) );
ao12f80 g760557 ( .a(n_20353), .b(n_20354), .c(n_19934), .o(n_20451) );
no02f80 g755572 ( .a(n_24598), .b(FE_OCPN1480_n_23872), .o(n_24616) );
in01f80 newInst_1302 ( .a(newNet_1301), .o(newNet_1302) );
in01f80 g751316 ( .a(n_28747), .o(n_28707) );
no02f80 g777803 ( .a(n_3287), .b(n_3286), .o(n_3288) );
no02f80 g757742 ( .a(FE_OCP_RBN3823_n_44061), .b(n_22517), .o(n_22559) );
no02f80 g739073 ( .a(n_41097), .b(n_41120), .o(n_41151) );
no02f80 g765795 ( .a(n_14978), .b(n_14977), .o(n_15070) );
na02f80 g746782 ( .a(n_32941), .b(n_32939), .o(n_33023) );
in01f80 g754280 ( .a(n_25931), .o(n_25932) );
in01f80 FE_OCPC1479_n_23872 ( .a(n_23872), .o(FE_OCPN1479_n_23872) );
in01f80 g773418 ( .a(n_7547), .o(n_7548) );
na02f80 g780757 ( .a(n_547), .b(n_396), .o(n_548) );
no03m80 g766808 ( .a(n_14454), .b(n_14352), .c(n_14456), .o(n_14489) );
in01f80 newInst_3080 ( .a(newNet_3079), .o(newNet_3080) );
in01f80 g774231 ( .a(n_6596), .o(n_6597) );
no02f80 g747578 ( .a(n_33481), .b(n_33440), .o(n_33465) );
no02f80 g738575 ( .a(n_41688), .b(n_41654), .o(n_41689) );
na02f80 g766788 ( .a(n_13667), .b(n_13634), .o(n_13691) );
in01f80 FE_OCP_RBC2189_n_7346 ( .a(n_7346), .o(FE_OCP_RBN2189_n_7346) );
in01f80 g778727 ( .a(n_2269), .o(n_2326) );
no02f80 g762031 ( .a(n_18206), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_), .o(n_18300) );
no02f80 g743375 ( .a(n_36689), .b(n_36579), .o(n_36705) );
no02f80 FE_RC_3995_0 ( .a(FE_RN_1732_0), .b(FE_OCP_RBN1332_n_20249), .o(n_20289) );
in01f80 newInst_1759 ( .a(newNet_1758), .o(newNet_1759) );
oa12f80 g780148 ( .a(n_1156), .b(n_1162), .c(n_1155), .o(n_1189) );
in01f80 newInst_2325 ( .a(newNet_2324), .o(newNet_2325) );
in01f80 newInst_880 ( .a(newNet_879), .o(newNet_880) );
na02f80 g737931 ( .a(n_42270), .b(n_42542), .o(n_42624) );
ao22s80 FE_RC_3695_0 ( .a(n_11819), .b(n_11830), .c(n_11829), .d(n_11881), .o(n_11978) );
na02f80 g777785 ( .a(n_3391), .b(FE_OCP_RBN3489_n_3390), .o(n_3488) );
in01f80 FE_RC_1757_0 ( .a(n_45685), .o(FE_RN_499_0) );
na02f80 FE_RC_2327_0 ( .a(FE_RN_886_0), .b(n_33099), .o(FE_RN_887_0) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_16_ ( .ck(newNet_2775), .d(n_46976), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_) );
in01f80 newInst_444 ( .a(newNet_443), .o(newNet_444) );
ms00f80 delay_sub_ln23_0_unr14_stage6_stallmux_q_reg ( .ck(newNet_1779), .d(n_20252), .o(n_44061) );
na02f80 g765900 ( .a(n_14826), .b(FE_OCPN1046_n_13570), .o(n_14906) );
no02f80 g759929 ( .a(n_21406), .b(n_21405), .o(n_21448) );
no02f80 g761338 ( .a(n_20069), .b(n_19993), .o(n_20117) );
in01f80 fopt783364 ( .a(n_38830), .o(n_44944) );
na02f80 g742522 ( .a(n_37535), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37560) );
na02f80 g739455 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .o(n_40809) );
in01f80 g774348 ( .a(n_6998), .o(n_6999) );
no02f80 g736837 ( .a(n_43215), .b(n_43214), .o(n_43258) );
na02f80 g778436 ( .a(n_2433), .b(n_2102), .o(n_2444) );
in01f80 fopt782969 ( .a(n_32338), .o(n_44432) );
na02f80 g744380 ( .a(n_35854), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36838) );
no02f80 g756270 ( .a(n_24673), .b(n_24672), .o(n_24674) );
no02f80 g768952 ( .a(n_11661), .b(n_11555), .o(n_11662) );
ao22s80 FE_RC_99_0 ( .a(FE_OCP_RBN1174_n_18981), .b(n_17815), .c(n_18981), .d(n_17783), .o(n_19075) );
na02f80 g742224 ( .a(FE_OCP_RBN3425_n_44881), .b(n_37598), .o(n_38049) );
no02f80 FE_RC_1916_0 ( .a(FE_RN_602_0), .b(n_19206), .o(FE_RN_603_0) );
ao12f80 g755249 ( .a(n_24881), .b(n_24975), .c(n_24823), .o(n_24989) );
no02f80 g751532 ( .a(n_28453), .b(n_28452), .o(n_28471) );
ao12f80 g768617 ( .a(n_12155), .b(n_12154), .c(n_12153), .o(n_12871) );
no02f80 g784404 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .o(n_46216) );
na02f80 g740423 ( .a(FE_OCP_RBN3029_n_39942), .b(n_39577), .o(n_40169) );
oa22f80 g764717 ( .a(n_15804), .b(n_15259), .c(n_15851), .d(n_15298), .o(n_15900) );
in01f80 g778563 ( .a(n_2342), .o(n_2406) );
in01f80 g740671 ( .a(n_39992), .o(n_39602) );
ao12f80 g766086 ( .a(n_14947), .b(n_14894), .c(n_14386), .o(n_14996) );
na02f80 g763921 ( .a(FE_OCP_RBN3294_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_), .o(n_17202) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_2_ ( .ck(newNet_2826), .d(n_9842), .o(delay_add_ln22_unr8_stage4_stallmux_q_2_) );
in01f80 g778744 ( .a(n_2251), .o(n_2252) );
in01f80 newInst_3164 ( .a(newNet_3163), .o(newNet_3164) );
na02f80 g761449 ( .a(n_19787), .b(n_19873), .o(n_19901) );
in01f80 g778006 ( .a(n_3580), .o(n_3563) );
in01f80 newInst_3626 ( .a(newNet_2595), .o(newNet_3626) );
in01f80 newInst_3117 ( .a(newNet_3116), .o(newNet_3117) );
in01f80 newInst_626 ( .a(newNet_625), .o(newNet_626) );
no02f80 g774308 ( .a(FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .o(n_6560) );
no02f80 g753399 ( .a(n_27041), .b(n_27040), .o(n_27361) );
no02f80 g762076 ( .a(FE_OCP_RBN2204_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_20_), .o(n_19014) );
no02f80 g755358 ( .a(n_24963), .b(n_24962), .o(n_25035) );
na02f80 g740718 ( .a(n_39449), .b(n_39418), .o(n_39523) );
no02f80 g773390 ( .a(n_7585), .b(n_7614), .o(n_7660) );
in01f80 g739448 ( .a(n_40769), .o(n_40718) );
in01f80 g772859 ( .a(n_8052), .o(n_8053) );
ao12f80 g760343 ( .a(n_20105), .b(n_20104), .c(n_20103), .o(n_21896) );
in01f80 FE_OCP_DRV_C3157_n_27062 ( .a(n_27062), .o(FE_OCP_DRV_N3157_n_27062) );
in01f80 g776094 ( .a(n_4867), .o(n_4868) );
in01f80 newInst_290 ( .a(newNet_197), .o(newNet_290) );
in01f80 g744313 ( .a(n_46245), .o(n_36849) );
ms00f80 sin_out_reg_10_ ( .ck(newNet_91), .d(n_43803), .o(sin_out_10) );
oa22f80 FE_RC_1484_0 ( .a(n_32287), .b(n_32546), .c(n_28336), .d(n_32513), .o(n_32594) );
in01f80 newInst_2920 ( .a(newNet_2051), .o(newNet_2920) );
in01f80 g774995 ( .a(n_6059), .o(n_6078) );
na02f80 g740155 ( .a(FE_OCP_RBN3721_n_39913), .b(n_39905), .o(n_40186) );
in01f80 g768018 ( .a(n_12651), .o(n_12652) );
no02f80 g740016 ( .a(n_39812), .b(n_39906), .o(n_39957) );
no02f80 g767353 ( .a(n_13447), .b(n_13404), .o(n_13508) );
in01f80 g747526 ( .a(n_32546), .o(n_32513) );
in01f80 g769939 ( .a(n_11158), .o(n_11249) );
na02f80 g758947 ( .a(n_21642), .b(n_21641), .o(n_21643) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_28_ ( .ck(newNet_2266), .d(FE_OCP_RBN3139_n_40568), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_) );
in01f80 g762231 ( .a(n_18148), .o(n_18190) );
in01f80 FE_OCP_RBC2840_n_4692 ( .a(FE_OCP_RBN2839_n_4692), .o(FE_OCP_RBN2840_n_4692) );
in01f80 newInst_351 ( .a(newNet_350), .o(newNet_351) );
na02f80 FE_RC_3608_0 ( .a(FE_RN_1577_0), .b(n_18954), .o(n_18984) );
in01f80 g763085 ( .a(n_17349), .o(n_17350) );
in01f80 newInst_3247 ( .a(newNet_3246), .o(newNet_3247) );
no02f80 g746940 ( .a(n_32862), .b(n_32861), .o(n_32879) );
in01f80 g777601 ( .a(n_5242), .o(n_3472) );
na02f80 FE_RC_2573_0 ( .a(FE_RN_1057_0), .b(n_43775), .o(n_43788) );
in01f80 g758963 ( .a(n_21636), .o(n_21637) );
no02f80 g778762 ( .a(n_2381), .b(n_2021), .o(n_2455) );
na02f80 g750396 ( .a(n_30590), .b(n_30589), .o(n_30591) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_6_ ( .ck(newNet_1926), .d(n_36885), .o(delay_sub_ln21_unr24_stage9_stallmux_q_6_) );
na02f80 g769381 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_11933) );
in01f80 g764352 ( .a(n_16392), .o(n_16393) );
in01f80 FE_OCP_RBC2995_n_35539 ( .a(FE_OCP_RBN2991_n_35539), .o(FE_OCP_RBN2995_n_35539) );
in01f80 g738995 ( .a(n_41492), .o(n_41187) );
oa12f80 g751348 ( .a(n_29433), .b(n_29432), .c(n_29431), .o(n_29908) );
in01f80 FE_RC_2096_0 ( .a(n_14758), .o(FE_RN_721_0) );
in01f80 g749793 ( .a(n_31625), .o(n_31626) );
ao12f80 g762853 ( .a(n_17840), .b(n_17839), .c(n_17838), .o(n_19354) );
oa12f80 g737360 ( .a(n_42580), .b(n_42807), .c(n_42514), .o(n_42848) );
ao12f80 g774224 ( .a(n_6644), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_8_), .o(n_6731) );
no02f80 g755169 ( .a(n_25045), .b(FE_OCPN1792_n_25044), .o(n_25116) );
na02f80 g755176 ( .a(n_25045), .b(FE_OCPN1792_n_25044), .o(n_25069) );
no02f80 g752284 ( .a(FE_OCP_RBN2126_n_44734), .b(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .o(n_28001) );
na02f80 g741753 ( .a(n_38493), .b(n_39324), .o(n_38494) );
in01f80 newInst_851 ( .a(newNet_850), .o(newNet_851) );
in01f80 g749104 ( .a(n_46956), .o(n_31017) );
in01f80 g757263 ( .a(n_23490), .o(n_23491) );
no02f80 FE_RC_3454_0 ( .a(FE_RN_1485_0), .b(FE_RN_772_0), .o(n_26753) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_22_ ( .ck(newNet_2651), .d(n_22718), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_) );
ao12f80 g760527 ( .a(n_20386), .b(n_20385), .c(n_20384), .o(n_21244) );
in01f80 g766981 ( .a(n_13557), .o(n_13556) );
in01f80 g777118 ( .a(n_3841), .o(n_3842) );
in01f80 g742660 ( .a(n_37618), .o(n_37548) );
in01f80 FE_RC_2042_0 ( .a(n_24794), .o(FE_RN_684_0) );
no02f80 g779081 ( .a(n_2087), .b(n_1832), .o(n_2100) );
in01f80 g775853 ( .a(n_5003), .o(n_6131) );
na02f80 g771981 ( .a(FE_OFN754_n_44461), .b(n_9369), .o(n_9516) );
no02f80 g749951 ( .a(FE_OCP_RBN2634_n_30213), .b(n_30278), .o(n_30292) );
in01f80 g755820 ( .a(n_24423), .o(n_24424) );
na02f80 g738370 ( .a(n_41700), .b(FE_OCP_RBN2314_n_41420), .o(n_41793) );
no02f80 g769737 ( .a(n_11254), .b(n_11253), .o(n_11269) );
in01f80 g780172 ( .a(n_1163), .o(n_1151) );
in01f80 newInst_2087 ( .a(newNet_234), .o(newNet_2087) );
in01f80 newInst_1684 ( .a(newNet_1683), .o(newNet_1684) );
in01f80 g780182 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_28_), .o(n_1095) );
in01f80 g779645 ( .a(n_1790), .o(n_1791) );
na02f80 g755239 ( .a(n_25096), .b(n_23891), .o(n_25176) );
no02f80 g740575 ( .a(n_39680), .b(n_38712), .o(n_39695) );
in01f80 g738297 ( .a(n_41823), .o(n_41824) );
in01f80 g749718 ( .a(n_31576), .o(n_31577) );
na02f80 g778262 ( .a(n_2895), .b(n_2894), .o(n_2918) );
in01f80 g750804 ( .a(n_31116), .o(n_30393) );
in01f80 FE_OCP_RBC2147_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2144_FE_OCPN861_n_45450), .o(FE_OCP_RBN2147_FE_OCPN861_n_45450) );
in01f80 g780672 ( .a(n_694), .o(n_713) );
in01f80 g736957 ( .a(n_43254), .o(n_43352) );
na02f80 g778259 ( .a(n_2836), .b(n_2894), .o(n_2887) );
oa12f80 FE_RC_1930_0 ( .a(FE_RN_611_0), .b(FE_RN_610_0), .c(n_29273), .o(n_29378) );
in01f80 g753653 ( .a(n_26622), .o(n_26652) );
no02f80 g769043 ( .a(FE_OCP_RBN2116_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n_11643) );
ao12f80 g743800 ( .a(n_44180), .b(n_35878), .c(n_35555), .o(n_35923) );
na02f80 g779105 ( .a(n_1987), .b(n_1834), .o(n_1988) );
ao12f80 g777391 ( .a(n_3217), .b(n_3416), .c(n_3199), .o(n_3424) );
no02f80 g769374 ( .a(n_45659), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n_12078) );
na02f80 g755138 ( .a(n_25551), .b(n_45635), .o(n_25645) );
in01f80 g765763 ( .a(FE_OCP_RBN2716_n_14982), .o(n_15103) );
no02f80 g749521 ( .a(n_30497), .b(n_30142), .o(n_30529) );
in01f80 FE_RC_145_0 ( .a(n_12039), .o(FE_RN_43_0) );
no02f80 FE_RC_3164_0 ( .a(FE_RN_1402_0), .b(FE_OCP_RBN3726_FE_RN_1787_0), .o(n_17137) );
no03m80 FE_RC_1642_0 ( .a(n_17289), .b(n_17410), .c(n_17485), .o(n_17517) );
in01f80 FE_RC_358_0 ( .a(n_17349), .o(FE_RN_105_0) );
in01f80 FE_OFC836_n_4575 ( .a(n_4575), .o(FE_OFN836_n_4575) );
in01f80 g747183 ( .a(n_32867), .o(n_32868) );
no02f80 g751729 ( .a(n_28348), .b(delay_add_ln22_unr17_stage7_stallmux_q_10_), .o(n_28357) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_21_ ( .ck(newNet_3143), .d(n_40486), .o(delay_add_ln22_unr27_stage10_stallmux_q_21_) );
na02f80 g775534 ( .a(n_5485), .b(n_5494), .o(n_5572) );
in01f80 FE_RC_4080_0 ( .a(FE_OCP_RBN2851_n_46982), .o(FE_RN_1780_0) );
oa12f80 g765629 ( .a(n_14851), .b(n_14830), .c(n_14794), .o(n_14944) );
in01f80 g752952 ( .a(n_27875), .o(n_27953) );
no02f80 FE_RC_2408_0 ( .a(FE_RN_948_0), .b(n_6959), .o(FE_RN_949_0) );
na02f80 g761031 ( .a(FE_OCP_RBN3829_n_19204), .b(n_19131), .o(n_19317) );
no02f80 g737352 ( .a(n_42830), .b(n_42368), .o(n_42839) );
in01f80 newInst_2214 ( .a(newNet_14), .o(newNet_2214) );
in01f80 newInst_1036 ( .a(newNet_1035), .o(newNet_1036) );
no02f80 g742107 ( .a(n_37892), .b(n_37851), .o(n_38010) );
in01f80 g765416 ( .a(n_15567), .o(n_15568) );
oa22f80 g780398 ( .a(n_881), .b(n_780), .c(n_803), .d(n_1159), .o(n_835) );
in01f80 g751804 ( .a(n_28960), .o(n_29008) );
in01f80 newInst_3396 ( .a(newNet_3395), .o(newNet_3396) );
in01f80 FE_RC_2997_0 ( .a(n_6447), .o(FE_RN_1311_0) );
no02f80 g741298 ( .a(n_44955), .b(n_38147), .o(n_38957) );
ao22s80 FE_RC_1254_0 ( .a(n_41325), .b(n_41344), .c(n_41353), .d(n_41340), .o(n_41364) );
na02f80 g761657 ( .a(n_19521), .b(n_19520), .o(n_19522) );
no02f80 g777871 ( .a(n_3157), .b(n_3156), .o(n_3158) );
in01f80 g746104 ( .a(n_33940), .o(n_34060) );
no02f80 g778314 ( .a(n_2798), .b(n_2797), .o(n_2847) );
na02f80 g752200 ( .a(n_28589), .b(n_28588), .o(n_28590) );
in01f80 newInst_2983 ( .a(newNet_2982), .o(newNet_2983) );
in01f80 g756830 ( .a(n_24153), .o(n_24131) );
no02f80 g780553 ( .a(n_713), .b(n_420), .o(n_754) );
in01f80 g762456 ( .a(n_18001), .o(n_18002) );
no02f80 FE_RC_181_0 ( .a(FE_RN_59_0), .b(n_12297), .o(n_12342) );
no02f80 FE_RC_3979_0 ( .a(n_29643), .b(FE_RN_1724_0), .o(n_29658) );
no02f80 g769912 ( .a(n_10992), .b(n_44463), .o(n_11048) );
na02f80 g739388 ( .a(n_45145), .b(n_40342), .o(n_40787) );
na02f80 g763151 ( .a(n_17479), .b(n_17478), .o(n_17580) );
in01f80 FE_OCPC959_n_3951 ( .a(FE_OCPN958_n_3951), .o(FE_OCPN959_n_3951) );
in01f80 g753266 ( .a(n_27256), .o(n_27295) );
in01f80 g765288 ( .a(n_16306), .o(n_16307) );
in01f80 newInst_191 ( .a(newNet_190), .o(newNet_191) );
in01f80 newInst_253 ( .a(newNet_74), .o(newNet_253) );
in01f80 newInst_1703 ( .a(newNet_1702), .o(newNet_1703) );
na02f80 g769064 ( .a(n_11659), .b(n_45224), .o(n_11769) );
in01f80 g748216 ( .a(n_32778), .o(n_32779) );
na02f80 g759635 ( .a(n_20727), .b(n_45067), .o(n_20793) );
in01f80 newInst_1652 ( .a(newNet_1583), .o(newNet_1652) );
in01f80 g757947 ( .a(n_22233), .o(n_22234) );
na02f80 g765649 ( .a(FE_OCP_RBN1189_n_14911), .b(n_14758), .o(n_14963) );
oa12f80 g777212 ( .a(n_3356), .b(n_3507), .c(n_3309), .o(n_3547) );
no02f80 g745693 ( .a(n_34367), .b(n_34430), .o(n_34481) );
in01f80 g742815 ( .a(n_37256), .o(n_37281) );
in01f80 g764805 ( .a(n_15700), .o(n_15699) );
in01f80 g764748 ( .a(n_15980), .o(n_15981) );
na02f80 g773541 ( .a(n_7474), .b(n_7473), .o(n_7475) );
ao12f80 g754985 ( .a(n_25774), .b(n_25773), .c(n_25772), .o(n_25867) );
in01f80 newInst_2238 ( .a(newNet_2237), .o(newNet_2238) );
na02f80 g753988 ( .a(n_26979), .b(n_26862), .o(n_27033) );
no02f80 g741956 ( .a(n_37976), .b(n_37902), .o(n_38041) );
no02f80 g747672 ( .a(n_32087), .b(n_31809), .o(n_32148) );
na02f80 g743169 ( .a(n_36879), .b(n_36897), .o(n_36912) );
na02f80 g767973 ( .a(n_12883), .b(n_13159), .o(n_13520) );
in01f80 g762169 ( .a(n_18247), .o(n_18201) );
na02f80 g759601 ( .a(n_20911), .b(n_20842), .o(n_20874) );
na02f80 g773817 ( .a(n_7144), .b(n_7063), .o(n_7145) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_4_ ( .ck(newNet_785), .d(n_1345), .o(delay_xor_ln21_unr3_stage2_stallmux_q_4_) );
in01f80 g744636 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n_36637) );
na02f80 g770219 ( .a(n_10741), .b(n_10786), .o(n_10902) );
in01f80 FE_OCP_RBC3536_n_13765 ( .a(FE_OCP_RBN3531_n_13765), .o(FE_OCP_RBN3536_n_13765) );
in01f80 g780550 ( .a(n_936), .o(n_750) );
in01f80 g737518 ( .a(n_42475), .o(n_42454) );
in01f80 g741990 ( .a(n_38108), .o(n_38109) );
in01f80 g738100 ( .a(n_42102), .o(n_42569) );
in01f80 g743803 ( .a(n_36369), .o(n_36370) );
oa12f80 g747395 ( .a(n_33747), .b(n_33746), .c(n_33745), .o(n_34389) );
in01f80 g750300 ( .a(n_29784), .o(n_29785) );
no02f80 g738564 ( .a(n_41604), .b(n_41725), .o(n_41761) );
oa12f80 g740929 ( .a(n_39064), .b(n_39214), .c(n_38994), .o(n_39306) );
oa12f80 g761101 ( .a(n_19037), .b(n_19142), .c(n_19081), .o(n_19152) );
ao12f80 g763714 ( .a(n_16603), .b(n_16646), .c(n_16641), .o(n_16690) );
oa22f80 FE_RC_3370_0 ( .a(n_32566), .b(n_32518), .c(n_28336), .d(n_32470), .o(n_32571) );
in01f80 newInst_1107 ( .a(newNet_874), .o(newNet_1107) );
no02f80 g779142 ( .a(n_1993), .b(n_1992), .o(n_1994) );
in01f80 g775575 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_10_), .o(n_5619) );
no02f80 g754435 ( .a(n_25635), .b(n_25401), .o(n_25656) );
no02f80 g743510 ( .a(n_37713), .b(n_46238), .o(n_37676) );
no02f80 g779011 ( .a(n_2174), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .o(n_2209) );
na02f80 g760920 ( .a(n_19313), .b(n_19286), .o(n_19362) );
in01f80 FE_OCP_RBC2288_n_2268 ( .a(n_2268), .o(FE_OCP_RBN2288_n_2268) );
oa12f80 g772609 ( .a(n_7423), .b(n_8191), .c(n_7384), .o(n_8261) );
in01f80 g757439 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_6_), .o(n_22828) );
no02f80 g746977 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .o(n_33104) );
in01f80 newInst_3338 ( .a(newNet_3337), .o(newNet_3338) );
na02f80 g760682 ( .a(n_19673), .b(n_19441), .o(n_19707) );
ao12f80 g741342 ( .a(n_38845), .b(n_38844), .c(n_38843), .o(n_39763) );
na02f80 g746103 ( .a(n_33874), .b(n_33850), .o(n_33959) );
in01f80 newInst_108 ( .a(newNet_107), .o(newNet_108) );
oa22f80 FE_RC_1643_0 ( .a(n_18956), .b(n_18509), .c(n_18955), .d(n_18510), .o(n_19064) );
na02f80 g773606 ( .a(n_47176), .b(n_6942), .o(n_7427) );
na02f80 g772880 ( .a(n_7992), .b(n_7991), .o(n_8039) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_13_ ( .ck(newNet_663), .d(n_46360), .o(delay_xor_ln21_unr9_stage4_stallmux_q_13_) );
no02f80 g766804 ( .a(n_13745), .b(n_13644), .o(n_13789) );
in01f80 g774816 ( .a(n_6395), .o(n_6370) );
na02f80 g760246 ( .a(FE_OCPN1261_n_20242), .b(n_19497), .o(n_20657) );
no02f80 g755863 ( .a(n_25193), .b(n_25140), .o(n_25199) );
oa22f80 FE_RC_871_0 ( .a(n_27493), .b(n_27723), .c(n_27724), .d(n_27492), .o(n_27835) );
na02f80 g773831 ( .a(FE_RN_953_0), .b(n_7134), .o(n_7416) );
no02f80 g760352 ( .a(n_20127), .b(FE_OCP_RBN2512_n_19884), .o(n_20153) );
no02f80 g752810 ( .a(n_27792), .b(n_27929), .o(n_28338) );
na02f80 g753158 ( .a(n_27327), .b(n_27375), .o(n_27484) );
na02f80 FE_RC_3723_0 ( .a(n_14960), .b(n_14846), .o(FE_RN_1638_0) );
no02f80 g767047 ( .a(n_14758), .b(n_14170), .o(n_14291) );
in01f80 FE_OCP_DRV_C1598_n_35644 ( .a(FE_OCP_DRV_N1597_n_35644), .o(FE_OCP_DRV_N1598_n_35644) );
in01f80 g755224 ( .a(n_25173), .o(n_25201) );
no03m80 g746874 ( .a(n_34074), .b(n_34082), .c(n_33701), .o(n_34169) );
oa12f80 FE_RC_3861_0 ( .a(FE_RN_1686_0), .b(FE_RN_1380_0), .c(n_31246), .o(n_31404) );
in01f80 newInst_1889 ( .a(newNet_442), .o(newNet_1889) );
ao12f80 g761293 ( .a(n_19787), .b(n_19983), .c(n_19571), .o(n_20010) );
no02f80 g776802 ( .a(n_4099), .b(n_2531), .o(n_4277) );
in01f80 g747538 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_), .o(n_32540) );
in01f80 newInst_2774 ( .a(newNet_2773), .o(newNet_2774) );
na02f80 g752202 ( .a(n_44825), .b(n_28130), .o(n_28635) );
na02f80 g740932 ( .a(n_39088), .b(n_39016), .o(n_39113) );
no02f80 g761553 ( .a(n_18948), .b(n_18919), .o(n_18920) );
oa12f80 g765105 ( .a(n_15976), .b(n_15884), .c(n_15874), .o(n_16310) );
in01f80 g758699 ( .a(n_21811), .o(n_21843) );
in01f80 FE_OCP_RBC2557_n_44576 ( .a(FE_OCP_RBN3550_n_44575), .o(FE_OCP_RBN2557_n_44576) );
na02f80 g770346 ( .a(n_10639), .b(n_10656), .o(n_10781) );
in01f80 g741818 ( .a(n_38418), .o(n_38419) );
na02f80 g776494 ( .a(n_4447), .b(n_4351), .o(n_4476) );
no02f80 g744001 ( .a(n_36098), .b(n_36144), .o(n_36268) );
na02f80 g776181 ( .a(n_4462), .b(n_4236), .o(n_4524) );
no02f80 g777131 ( .a(n_3767), .b(n_3756), .o(n_3985) );
ao22s80 g736422 ( .a(n_43727), .b(n_43548), .c(n_43726), .d(n_43547), .o(n_43770) );
in01f80 newInst_20 ( .a(newNet_19), .o(newNet_20) );
in01f80 newInst_3375 ( .a(newNet_3374), .o(newNet_3375) );
in01f80 g773391 ( .a(n_7764), .o(n_7765) );
in01f80 FE_OCP_RBC2539_n_8781 ( .a(n_8781), .o(FE_OCP_RBN2539_n_8781) );
in01f80 FE_OCP_RBC1132_n_12827 ( .a(n_12827), .o(FE_OCP_RBN1132_n_12827) );
na02f80 g749064 ( .a(n_30940), .b(n_30915), .o(n_30998) );
in01f80 newInst_3092 ( .a(newNet_3091), .o(newNet_3092) );
na02f80 g749353 ( .a(n_30542), .b(n_27014), .o(n_30611) );
in01f80 g777827 ( .a(n_3697), .o(n_3663) );
in01f80 g766980 ( .a(n_13557), .o(n_13577) );
no02f80 g745357 ( .a(n_36154), .b(n_36079), .o(n_36209) );
oa12f80 g780103 ( .a(n_1210), .b(n_45818), .c(n_1208), .o(n_1217) );
ao12f80 g752054 ( .a(n_28014), .b(FE_OCPN877_n_44734), .c(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .o(n_28229) );
in01f80 newInst_3398 ( .a(newNet_3397), .o(newNet_3398) );
in01f80 g738758 ( .a(n_41479), .o(n_41480) );
na02f80 g774363 ( .a(n_6844), .b(n_6939), .o(n_7449) );
oa12f80 g745173 ( .a(n_34405), .b(n_34656), .c(n_34340), .o(n_34784) );
no02f80 g776769 ( .a(n_3737), .b(n_2988), .o(n_3858) );
ao22s80 g737408 ( .a(n_42732), .b(n_42698), .c(n_42731), .d(n_42699), .o(n_43106) );
in01f80 g772879 ( .a(n_8039), .o(n_8040) );
in01f80 g739324 ( .a(n_40843), .o(n_40886) );
in01f80 FE_OCP_RBC3401_n_37670 ( .a(n_37670), .o(FE_OCP_RBN3401_n_37670) );
ms00f80 cos_out_reg_30_ ( .ck(newNet_3694), .d(n_43906), .o(cos_out_30) );
no02f80 g748368 ( .a(n_32726), .b(n_32725), .o(n_32727) );
in01f80 FE_RC_3588_0 ( .a(FE_RN_1565_0), .o(FE_RN_1564_0) );
in01f80 newInst_1017 ( .a(newNet_388), .o(newNet_1017) );
na02f80 g758078 ( .a(n_44277), .b(n_21216), .o(n_22232) );
in01f80 FE_OCPC1778_n_37744 ( .a(FE_OCPN1777_n_37744), .o(FE_OCPN1778_n_37744) );
in01f80 FE_OCP_RBC1990_delay_xor_ln23_unr6_stage3_stallmux_q ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .o(FE_OCP_RBN1990_delay_xor_ln23_unr6_stage3_stallmux_q) );
ao22s80 g780301 ( .a(n_950), .b(n_1098), .c(n_864), .d(n_1099), .o(n_998) );
in01f80 g756816 ( .a(n_24032), .o(n_24033) );
no02f80 FE_RC_4050_0 ( .a(n_36015), .b(FE_RN_1760_0), .o(FE_RN_1761_0) );
oa12f80 g770301 ( .a(FE_OCP_RBN3654_n_10100), .b(n_10541), .c(n_8908), .o(n_10569) );
in01f80 g740764 ( .a(n_39514), .o(n_39515) );
na02f80 g750043 ( .a(n_29809), .b(n_28830), .o(n_29901) );
no02f80 g766787 ( .a(n_14081), .b(FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_14082) );
in01f80 FE_OFC833_n_19885 ( .a(n_19885), .o(FE_OFN833_n_19885) );
na02f80 g755576 ( .a(n_24436), .b(n_22111), .o(n_24452) );
na02f80 FE_RC_2676_0 ( .a(FE_RN_1118_0), .b(n_4233), .o(FE_RN_1119_0) );
no02f80 g771885 ( .a(n_8743), .b(n_7577), .o(n_8788) );
in01f80 FE_RC_1077_0 ( .a(n_12543), .o(FE_RN_319_0) );
in01f80 FE_OCP_RBC3840_n_19513 ( .a(FE_OCP_RBN3839_n_19513), .o(FE_OCP_RBN3840_n_19513) );
na02f80 g774475 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .o(n_6857) );
in01f80 FE_RC_2580_0 ( .a(n_2880), .o(FE_RN_1064_0) );
ao12f80 g747089 ( .a(n_33996), .b(n_33995), .c(n_33994), .o(n_34696) );
oa22f80 g758602 ( .a(n_22431), .b(n_21777), .c(n_22453), .d(n_21776), .o(n_22548) );
no02f80 g740381 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39881), .o(n_40274) );
na02f80 g762625 ( .a(n_18294), .b(n_18293), .o(n_18295) );
oa12f80 g780299 ( .a(n_750), .b(n_903), .c(n_795), .o(n_960) );
in01f80 FE_OCP_RBC3626_n_38870 ( .a(FE_OCP_RBN2685_n_38870), .o(FE_OCP_RBN3626_n_38870) );
na02f80 g737581 ( .a(n_42402), .b(n_42364), .o(n_42425) );
in01f80 newInst_1932 ( .a(newNet_1756), .o(newNet_1932) );
no02f80 g768503 ( .a(n_45659), .b(delay_xor_ln21_unr9_stage4_stallmux_q_16_), .o(n_12355) );
no02f80 g760404 ( .a(n_20125), .b(FE_OCP_RBN3844_FE_RN_1242_0), .o(n_20187) );
in01f80 FE_OCPC913_n_43022 ( .a(FE_OCPN911_n_43022), .o(FE_OCPN913_n_43022) );
ao12f80 g747390 ( .a(n_32634), .b(FE_OCP_RBN2103_n_44962), .c(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .o(n_32651) );
oa12f80 g783846 ( .a(n_25824), .b(n_25678), .c(n_25707), .o(n_45532) );
na02f80 g751589 ( .a(FE_OCP_RBN2192_n_28597), .b(n_28646), .o(n_28718) );
in01f80 FE_OCP_DRV_C1606_n_31445 ( .a(FE_OCP_DRV_N1605_n_31445), .o(FE_OCP_DRV_N1606_n_31445) );
in01f80 g779103 ( .a(n_2076), .o(n_2065) );
in01f80 g751764 ( .a(n_28303), .o(n_28304) );
in01f80 newInst_42 ( .a(newNet_24), .o(newNet_42) );
na02f80 g771753 ( .a(n_10159), .b(n_10208), .o(n_10239) );
oa12f80 g775476 ( .a(n_5617), .b(n_5624), .c(n_5616), .o(n_5724) );
ao22s80 g763134 ( .a(n_17481), .b(n_17435), .c(n_17397), .d(n_17434), .o(n_18854) );
na02f80 g780815 ( .a(n_380), .b(n_379), .o(n_381) );
na02f80 g746531 ( .a(n_33450), .b(n_33377), .o(n_33451) );
oa22f80 g758738 ( .a(n_21794), .b(n_21759), .c(n_21733), .d(n_21760), .o(n_21851) );
in01f80 newInst_102 ( .a(newNet_60), .o(newNet_102) );
in01f80 FE_RC_4068_0 ( .a(FE_OCPN1783_n_26801), .o(FE_RN_1771_0) );
in01f80 fopt782745 ( .a(n_21119), .o(n_44158) );
in01f80 g763662 ( .a(n_16900), .o(n_16893) );
in01f80 g751883 ( .a(n_29073), .o(n_29074) );
in01f80 g749797 ( .a(n_31454), .o(n_31428) );
in01f80 FE_OCP_RBC2201_n_12808 ( .a(n_12808), .o(FE_OCP_RBN2201_n_12808) );
in01f80 g770544 ( .a(n_10363), .o(n_10364) );
no02f80 g779764 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .o(n_1619) );
oa22f80 g763871 ( .a(n_16961), .b(n_16308), .c(n_16960), .d(n_16309), .o(n_17102) );
in01f80 g758575 ( .a(n_21997), .o(n_21998) );
ao12f80 g750353 ( .a(n_30636), .b(n_30663), .c(n_30635), .o(n_31210) );
in01f80 FE_RC_2246_0 ( .a(n_37092), .o(FE_RN_825_0) );
in01f80 FE_OCPC898_n_44776 ( .a(FE_OCPN896_n_44776), .o(FE_OCPN898_n_44776) );
no02f80 g758950 ( .a(n_21573), .b(n_21352), .o(n_21610) );
na03f80 g747229 ( .a(n_33498), .b(n_33764), .c(n_33513), .o(n_33931) );
oa12f80 g778546 ( .a(n_2720), .b(n_3297), .c(n_2744), .o(n_3489) );
oa22f80 FE_RC_946_0 ( .a(n_20231), .b(n_22875), .c(n_22833), .d(n_44329), .o(n_22949) );
no02f80 g739286 ( .a(n_40850), .b(n_40849), .o(n_40878) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_0_ ( .ck(newNet_2429), .d(n_35210), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_) );
in01f80 g747553 ( .a(n_32311), .o(n_32286) );
na02f80 g737923 ( .a(n_42201), .b(n_42304), .o(n_42360) );
in01f80 g772914 ( .a(n_46991), .o(n_8071) );
in01f80 g748568 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_), .o(n_31650) );
in01f80 FE_RC_53_0 ( .a(n_4407), .o(FE_RN_13_0) );
ao12f80 g761777 ( .a(n_19198), .b(n_19197), .c(n_19196), .o(n_19291) );
in01f80 FE_OCP_RBC3072_n_43230 ( .a(FE_OCP_RBN3069_n_43230), .o(FE_OCP_RBN3072_n_43230) );
no02f80 g740657 ( .a(n_39524), .b(n_39529), .o(n_39571) );
ao12f80 g752061 ( .a(n_28263), .b(n_28709), .c(n_28214), .o(n_28757) );
in01f80 newInst_1219 ( .a(newNet_1218), .o(newNet_1219) );
in01f80 g750282 ( .a(n_30835), .o(n_30836) );
ao22s80 FE_RC_4271_0 ( .a(FE_OCP_RBN3799_delay_xor_ln22_unr12_stage5_stallmux_q_0_), .b(FE_OCP_RBN3214_n_44365), .c(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .d(FE_OCP_RBN3205_n_44365), .o(n_16799) );
oa12f80 g741769 ( .a(n_38456), .b(n_38455), .c(n_38454), .o(n_38553) );
in01f80 g742920 ( .a(n_37116), .o(n_37117) );
in01f80 g759738 ( .a(n_21409), .o(n_21566) );
in01f80 newInst_3111 ( .a(newNet_2683), .o(newNet_3111) );
ao12f80 g756886 ( .a(n_23803), .b(n_23986), .c(n_23985), .o(n_23987) );
in01f80 g741943 ( .a(n_38141), .o(n_38142) );
na02f80 g748806 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .o(n_32558) );
oa12f80 g779140 ( .a(n_1886), .b(n_1885), .c(n_1884), .o(n_2363) );
in01f80 g766349 ( .a(n_14197), .o(n_14196) );
na02f80 g752587 ( .a(FE_OCP_RBN3102_n_27571), .b(n_27504), .o(n_27597) );
no02f80 g740007 ( .a(n_40189), .b(n_40033), .o(n_40226) );
oa12f80 g768133 ( .a(n_11892), .b(n_12623), .c(n_12083), .o(n_12645) );
na02f80 g744840 ( .a(n_35063), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35119) );
no02f80 g771974 ( .a(n_44498), .b(n_9939), .o(n_9951) );
na02f80 g754868 ( .a(n_25626), .b(n_25591), .o(n_25670) );
na02f80 g741016 ( .a(n_38837), .b(FE_OCP_RBN2639_n_38806), .o(n_38897) );
na02f80 g769931 ( .a(n_11006), .b(n_9742), .o(n_11076) );
no02f80 g777986 ( .a(n_3031), .b(n_2333), .o(n_3032) );
oa22f80 FE_RC_800_0 ( .a(n_8189), .b(n_8835), .c(FE_OCP_RBN3475_n_7886), .d(FE_OCP_RBN2497_n_8835), .o(n_8953) );
in01f80 g748800 ( .a(n_32537), .o(n_32452) );
na02f80 g759922 ( .a(FE_OCP_RBN3677_n_21051), .b(n_20157), .o(n_21299) );
na02f80 g768417 ( .a(n_12381), .b(FE_OCPN1002_n_45660), .o(n_12414) );
in01f80 g762661 ( .a(n_18253), .o(n_18254) );
in01f80 g758997 ( .a(n_21572), .o(n_21606) );
na02f80 g777095 ( .a(n_3899), .b(n_3700), .o(n_4071) );
oa22f80 FE_RC_1520_0 ( .a(n_22458), .b(n_22745), .c(n_22457), .d(n_22707), .o(n_22901) );
in01f80 g737236 ( .a(FE_OCP_RBN2915_n_42947), .o(n_42961) );
na02f80 g769724 ( .a(n_11293), .b(n_11292), .o(n_11374) );
no02f80 g740830 ( .a(n_39218), .b(n_39301), .o(n_39351) );
in01f80 g760558 ( .a(n_20018), .o(n_20019) );
no02f80 g742093 ( .a(FE_OCP_RBN3452_n_37945), .b(n_37567), .o(n_38102) );
na02f80 FE_RC_3523_0 ( .a(FE_RN_1522_0), .b(n_34767), .o(FE_RN_1523_0) );
na02f80 g775228 ( .a(n_6003), .b(n_6011), .o(n_6127) );
in01f80 g762348 ( .a(n_18497), .o(n_18582) );
ao12f80 g738329 ( .a(n_41553), .b(n_41596), .c(n_41552), .o(n_42209) );
no02f80 g776227 ( .a(n_4814), .b(n_4487), .o(n_4860) );
in01f80 g776682 ( .a(n_5603), .o(n_3971) );
in01f80 g751288 ( .a(n_29744), .o(n_29722) );
no03m80 g777047 ( .a(n_5091), .b(n_4974), .c(n_5090), .o(n_5092) );
no02f80 g742998 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n_37000) );
in01f80 g776546 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .o(n_6761) );
oa12f80 g777591 ( .a(n_3165), .b(n_3414), .c(n_3123), .o(n_3507) );
in01f80 newInst_2082 ( .a(newNet_2081), .o(newNet_2082) );
no02f80 g784603 ( .a(n_16241), .b(n_14805), .o(n_46426) );
no02f80 g762073 ( .a(FE_OCP_RBN2205_n_18242), .b(n_18329), .o(n_18426) );
no02f80 g736609 ( .a(n_43624), .b(n_43467), .o(n_43644) );
no02f80 g756577 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n_23878) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_13_ ( .ck(newNet_2021), .d(n_11061), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_) );
ao22s80 FE_RC_3046_0 ( .a(n_27315), .b(FE_OCP_RBN2934_n_31010), .c(n_27366), .d(n_31010), .o(n_31111) );
in01f80 newInst_2163 ( .a(newNet_2162), .o(newNet_2163) );
no02f80 g778434 ( .a(n_3127), .b(FE_OCPN1234_n_2414), .o(n_2563) );
oa12f80 g775485 ( .a(n_5535), .b(n_5622), .c(n_5412), .o(n_5690) );
no02f80 FE_RC_2046_0 ( .a(FE_RN_687_0), .b(n_25588), .o(FE_RN_688_0) );
ao22s80 g777234 ( .a(n_3639), .b(n_3113), .c(n_3638), .d(n_4719), .o(n_3661) );
in01f80 newInst_908 ( .a(newNet_907), .o(newNet_908) );
oa12f80 g741912 ( .a(n_38319), .b(n_38170), .c(n_38317), .o(n_38432) );
in01f80 newInst_1 ( .a(newNet_0), .o(newNet_1) );
no02f80 g762743 ( .a(FE_OCP_RBN2145_FE_OCPN861_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .o(n_17967) );
in01f80 newInst_443 ( .a(newNet_442), .o(newNet_443) );
in01f80 g768932 ( .a(n_11938), .o(n_11939) );
na02f80 g755683 ( .a(n_25371), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25372) );
no02f80 g755489 ( .a(n_24601), .b(n_24602), .o(n_24603) );
in01f80 g777544 ( .a(n_4606), .o(n_4759) );
no02f80 g737251 ( .a(n_42914), .b(n_42610), .o(n_42930) );
in01f80 FE_OCPC1028_n_4182 ( .a(FE_OCPN1027_n_4182), .o(FE_OCPN1028_n_4182) );
in01f80 newInst_543 ( .a(newNet_542), .o(newNet_543) );
no02f80 g775279 ( .a(n_5609), .b(n_4759), .o(n_5653) );
in01f80 FE_OCP_RBC2949_n_10852 ( .a(FE_OCP_RBN3693_n_10852), .o(FE_OCP_RBN2949_n_10852) );
in01f80 drc1 ( .a(n_47236), .o(n_47239) );
in01f80 g756953 ( .a(n_23701), .o(n_23989) );
in01f80 newInst_3304 ( .a(newNet_3303), .o(newNet_3304) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_3_ ( .ck(newNet_2154), .d(n_1167), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_) );
in01f80 newInst_2940 ( .a(newNet_2939), .o(newNet_2940) );
na02f80 g740379 ( .a(n_39803), .b(n_39881), .o(n_39852) );
ao22s80 g780739 ( .a(n_601), .b(n_571), .c(n_599), .d(n_572), .o(n_744) );
in01f80 g779563 ( .a(n_1554), .o(n_1555) );
na02f80 g744552 ( .a(n_35438), .b(n_35437), .o(n_35439) );
in01f80 g757743 ( .a(n_22820), .o(n_22595) );
no02f80 g776773 ( .a(FE_OCP_RBN3602_n_3913), .b(n_3625), .o(n_4056) );
na02f80 g754237 ( .a(n_25954), .b(n_25748), .o(n_25989) );
oa12f80 g762306 ( .a(n_18384), .b(n_18383), .c(n_18382), .o(n_18734) );
na02f80 g753117 ( .a(n_27175), .b(n_27143), .o(n_27348) );
na02f80 FE_RC_2807_0 ( .a(n_13634), .b(n_13616), .o(FE_RN_1201_0) );
oa12f80 g784691 ( .a(n_3100), .b(n_2940), .c(n_3049), .o(n_47021) );
oa22f80 FE_RC_3199_0 ( .a(n_16801), .b(n_16745), .c(n_16802), .d(n_16746), .o(n_16987) );
no02f80 g755105 ( .a(n_24161), .b(n_25201), .o(n_25319) );
no02f80 g769778 ( .a(n_11284), .b(n_11283), .o(n_11303) );
in01f80 FE_OCPC1405_n_25859 ( .a(n_25859), .o(FE_OCPN1405_n_25859) );
no02f80 FE_RC_1094_0 ( .a(FE_RN_321_0), .b(FE_RN_322_0), .o(FE_RN_323_0) );
in01f80 g781352 ( .a(beta_18), .o(n_11) );
no02f80 g756169 ( .a(n_24102), .b(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24128) );
no02f80 FE_RC_412_0 ( .a(FE_RN_120_0), .b(FE_RN_121_0), .o(FE_RN_122_0) );
no02f80 g772401 ( .a(n_8513), .b(FE_OCP_RBN3464_n_7886), .o(n_8544) );
na02f80 g762276 ( .a(n_45002), .b(n_18414), .o(n_18624) );
no02f80 g765088 ( .a(n_16101), .b(n_16098), .o(n_16261) );
na02f80 g775772 ( .a(n_5028), .b(FE_OCPN846_n_4046), .o(n_5159) );
na02f80 g746406 ( .a(n_35020), .b(n_34760), .o(n_34778) );
in01f80 g775207 ( .a(n_5955), .o(n_5962) );
no02f80 g749708 ( .a(n_29970), .b(n_29930), .o(n_29931) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_24_ ( .ck(newNet_1310), .d(n_1260), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_) );
in01f80 FE_OCP_RBC3611_FE_OCPN1797_n_20333 ( .a(FE_OCP_RBN3610_FE_OCPN1797_n_20333), .o(FE_OCP_RBN3611_FE_OCPN1797_n_20333) );
in01f80 FE_OCP_RBC2739_n_20432 ( .a(n_20432), .o(FE_OCP_RBN2739_n_20432) );
na02f80 FE_RC_2127_0 ( .a(FE_RN_741_0), .b(n_25455), .o(FE_RN_742_0) );
no02f80 g769770 ( .a(FE_OCP_RBN3005_n_11087), .b(n_44516), .o(n_11148) );
no02f80 g751594 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .o(n_28678) );
in01f80 g756860 ( .a(n_23348), .o(n_23349) );
na02f80 g738668 ( .a(n_41684), .b(n_41715), .o(n_41779) );
na02f80 g749830 ( .a(n_31311), .b(n_30968), .o(n_31528) );
in01f80 newInst_2319 ( .a(newNet_2318), .o(newNet_2319) );
in01f80 g762008 ( .a(n_19913), .o(n_18886) );
in01f80 g747400 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .o(n_32389) );
oa12f80 g780035 ( .a(n_891), .b(n_1245), .c(n_844), .o(n_1253) );
in01f80 newInst_2155 ( .a(newNet_669), .o(newNet_2155) );
in01f80 fopt783804 ( .a(n_45488), .o(n_45487) );
na02f80 g776618 ( .a(n_4240), .b(n_4134), .o(n_4241) );
in01f80 g753533 ( .a(n_26783), .o(n_26784) );
in01f80 g758835 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_7_), .o(n_21785) );
na02f80 g752280 ( .a(n_28098), .b(n_27865), .o(n_27867) );
na02f80 g738489 ( .a(n_41387), .b(n_41433), .o(n_41523) );
in01f80 g752154 ( .a(n_28062), .o(n_28063) );
na02f80 g768331 ( .a(n_12465), .b(n_12349), .o(n_12531) );
no02f80 g771199 ( .a(n_9091), .b(n_8189), .o(n_9145) );
no02f80 g751033 ( .a(n_28853), .b(n_28832), .o(n_28833) );
na02f80 g748980 ( .a(n_30948), .b(n_31011), .o(n_31054) );
in01f80 g773651 ( .a(n_7351), .o(n_7352) );
in01f80 FE_OCPC927_n_26231 ( .a(n_26231), .o(FE_OCPN927_n_26231) );
na02f80 g756000 ( .a(n_25188), .b(n_24275), .o(n_25407) );
ao12f80 g773629 ( .a(n_6858), .b(n_47180), .c(n_6887), .o(n_7409) );
na02f80 g754127 ( .a(n_26834), .b(n_26382), .o(n_26974) );
in01f80 g748361 ( .a(n_31825), .o(n_31826) );
in01f80 g744479 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_2_), .o(n_35497) );
in01f80 g773647 ( .a(n_7368), .o(n_7369) );
na02f80 g758165 ( .a(n_44268), .b(n_21367), .o(n_22219) );
in01f80 g760052 ( .a(n_20672), .o(n_20673) );
no02f80 g766014 ( .a(n_47256), .b(n_14709), .o(n_14745) );
na02f80 g756617 ( .a(n_23545), .b(n_23519), .o(n_23520) );
in01f80 g750919 ( .a(n_28977), .o(n_28978) );
no02f80 g741276 ( .a(FE_OCP_RBN2552_n_44921), .b(n_38514), .o(n_39041) );
in01f80 g761702 ( .a(n_18887), .o(n_18888) );
in01f80 newInst_1627 ( .a(newNet_385), .o(newNet_1627) );
in01f80 g772767 ( .a(n_9304), .o(n_8147) );
in01f80 g752589 ( .a(n_27602), .o(n_27595) );
na02f80 g740875 ( .a(n_39168), .b(n_39111), .o(n_39264) );
no02f80 g763527 ( .a(FE_OCP_RBN3082_n_16977), .b(n_16117), .o(n_17165) );
in01f80 g770168 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_), .o(n_12452) );
ao12f80 g756506 ( .a(n_23854), .b(n_23843), .c(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n_23919) );
in01f80 fopt782729 ( .a(n_34066), .o(n_44100) );
in01f80 newInst_1515 ( .a(newNet_1514), .o(newNet_1515) );
na02f80 g776644 ( .a(n_4229), .b(n_4228), .o(n_4296) );
in01f80 g760593 ( .a(n_19915), .o(n_19916) );
na02f80 g749006 ( .a(n_31096), .b(n_31078), .o(n_31198) );
in01f80 FE_OCP_RBC2163_n_12312 ( .a(n_12312), .o(FE_OCP_RBN2163_n_12312) );
na02f80 g743680 ( .a(n_36329), .b(n_35864), .o(n_36349) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_20_ ( .ck(newNet_3533), .d(n_22701), .o(delay_add_ln22_unr14_stage6_stallmux_q_20_) );
na02f80 g742844 ( .a(n_37200), .b(n_37197), .o(n_37198) );
in01f80 newInst_1744 ( .a(newNet_1743), .o(newNet_1744) );
no02f80 g738042 ( .a(n_42120), .b(n_42111), .o(n_42309) );
oa12f80 g747855 ( .a(n_33392), .b(n_33552), .c(n_33027), .o(n_33553) );
na02f80 g765666 ( .a(n_15036), .b(n_15035), .o(n_15071) );
in01f80 g750159 ( .a(n_30210), .o(n_30211) );
in01f80 g736419 ( .a(n_43798), .o(n_43799) );
no02f80 g745516 ( .a(n_34565), .b(n_34564), .o(n_34566) );
no02f80 g762260 ( .a(n_18523), .b(n_18497), .o(n_18615) );
in01f80 g739149 ( .a(n_40964), .o(n_40925) );
na02f80 g736720 ( .a(n_43103), .b(n_43141), .o(n_43282) );
in01f80 g741760 ( .a(n_38457), .o(n_38458) );
in01f80 g765252 ( .a(n_15884), .o(n_15634) );
in01f80 g754340 ( .a(n_25826), .o(n_27142) );
na02f80 g755278 ( .a(n_25010), .b(n_24985), .o(n_25095) );
in01f80 g768623 ( .a(n_12321), .o(n_12322) );
no02f80 g741172 ( .a(FE_OCP_RBN2635_n_38806), .b(n_38859), .o(n_38885) );
oa22f80 FE_RC_1474_0 ( .a(n_24059), .b(n_27784), .c(n_27845), .d(n_27757), .o(n_27846) );
oa12f80 g778247 ( .a(n_2947), .b(n_2946), .c(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n_2948) );
na02f80 g761697 ( .a(n_18852), .b(n_18481), .o(n_18889) );
in01f80 g777301 ( .a(n_4576), .o(n_4577) );
no02f80 g752793 ( .a(n_28198), .b(n_28199), .o(n_28214) );
in01f80 g768094 ( .a(n_12627), .o(n_12628) );
in01f80 FE_RC_4206_0 ( .a(n_18140), .o(FE_RN_1841_0) );
na02f80 g761260 ( .a(n_19055), .b(n_17783), .o(n_19056) );
oa22f80 g775380 ( .a(n_5757), .b(n_5563), .c(n_5756), .d(n_5564), .o(n_5913) );
in01f80 g773556 ( .a(n_7422), .o(n_7435) );
oa22f80 FE_RC_717_0 ( .a(n_7361), .b(n_8074), .c(n_7362), .d(n_8075), .o(n_8187) );
in01f80 g764016 ( .a(n_18032), .o(n_19418) );
no02f80 g762967 ( .a(FE_OCP_RBN2141_FE_OCPN861_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_10_), .o(n_17765) );
in01f80 g758790 ( .a(n_21684), .o(n_21618) );
na02f80 g763159 ( .a(n_17009), .b(n_16879), .o(n_17146) );
in01f80 g738107 ( .a(n_42100), .o(n_42099) );
in01f80 g758901 ( .a(n_21761), .o(n_21762) );
in01f80 g771319 ( .a(n_9091), .o(n_9148) );
in01f80 g753170 ( .a(n_27519), .o(n_27520) );
oa12f80 g750771 ( .a(n_29156), .b(n_29313), .c(n_29158), .o(n_29436) );
in01f80 g750451 ( .a(n_31223), .o(n_30615) );
in01f80 g768979 ( .a(n_11734), .o(n_11735) );
na02f80 g754102 ( .a(n_25999), .b(FE_OFN737_n_22641), .o(n_26032) );
na02f80 g743452 ( .a(n_36539), .b(n_36521), .o(n_36583) );
in01f80 newInst_2587 ( .a(newNet_2229), .o(newNet_2587) );
in01f80 FE_OCP_RBC3521_n_19663 ( .a(n_19663), .o(FE_OCP_RBN3521_n_19663) );
na02f80 g772234 ( .a(n_8609), .b(FE_OCP_RBN3467_n_7886), .o(n_8678) );
in01f80 g769758 ( .a(n_11200), .o(n_11201) );
ao12f80 g745772 ( .a(n_34178), .b(n_44102), .c(n_33632), .o(n_34662) );
in01f80 newInst_270 ( .a(newNet_269), .o(newNet_270) );
in01f80 g746807 ( .a(n_33267), .o(n_33268) );
ao12f80 g752458 ( .a(n_27507), .b(n_27672), .c(n_27326), .o(n_27673) );
in01f80 newInst_766 ( .a(newNet_239), .o(newNet_766) );
no02f80 g771835 ( .a(n_9219), .b(n_9324), .o(n_9263) );
no02f80 g748047 ( .a(n_32026), .b(n_31952), .o(n_32107) );
ao12f80 g752415 ( .a(n_28380), .b(n_28401), .c(n_28379), .o(n_28879) );
no02f80 g784412 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n_46224) );
in01f80 newInst_2715 ( .a(newNet_2714), .o(newNet_2715) );
no02f80 g745129 ( .a(n_34749), .b(n_34435), .o(n_34790) );
na02f80 g776473 ( .a(n_4385), .b(n_4358), .o(n_4398) );
in01f80 g749885 ( .a(n_30176), .o(n_30177) );
no02f80 g774493 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .o(n_6696) );
oa12f80 g767444 ( .a(n_12563), .b(n_13009), .c(n_12549), .o(n_13139) );
in01f80 g773796 ( .a(n_7218), .o(n_7203) );
in01f80 newInst_501 ( .a(newNet_500), .o(newNet_501) );
no02f80 g756550 ( .a(n_23572), .b(n_22859), .o(n_23884) );
no02f80 g770240 ( .a(n_10363), .b(n_10518), .o(n_10595) );
oa22f80 FE_RC_1377_0 ( .a(FE_OCP_RBN3606_n_8981), .b(n_10865), .c(n_10712), .d(n_10863), .o(n_11008) );
no02f80 g741135 ( .a(n_38943), .b(n_39043), .o(n_39072) );
na02f80 g767803 ( .a(n_12925), .b(n_13248), .o(n_13088) );
in01f80 newInst_3649 ( .a(newNet_3648), .o(newNet_3649) );
in01f80 g749669 ( .a(FE_RN_1594_0), .o(n_31795) );
ao22s80 FE_RC_1084_0 ( .a(n_6908), .b(n_6731), .c(n_6909), .d(n_6732), .o(n_7020) );
no02f80 g756420 ( .a(n_25002), .b(n_24275), .o(n_24276) );
in01f80 newInst_3237 ( .a(newNet_3236), .o(newNet_3237) );
in01f80 g749040 ( .a(n_32292), .o(n_32293) );
na02f80 FE_RC_838_0 ( .a(n_9261), .b(FE_RN_251_0), .o(n_9362) );
in01f80 g755406 ( .a(n_24830), .o(n_24831) );
in01f80 g773194 ( .a(n_7917), .o(n_7918) );
in01f80 newInst_3669 ( .a(newNet_1922), .o(newNet_3669) );
ao12f80 g749600 ( .a(n_30462), .b(n_30461), .c(n_30460), .o(n_31773) );
no02f80 g748397 ( .a(n_31518), .b(n_31599), .o(n_31601) );
na02f80 g740505 ( .a(n_39684), .b(n_39677), .o(n_39710) );
no02f80 g756596 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .o(n_23872) );
no02f80 g756472 ( .a(n_23639), .b(n_23613), .o(n_23661) );
in01f80 g749545 ( .a(n_30409), .o(n_30389) );
oa22f80 g779894 ( .a(n_44659), .b(n_1092), .c(n_44623), .d(n_1050), .o(n_1292) );
no02f80 FE_RC_998_0 ( .a(FE_RN_287_0), .b(n_22889), .o(n_23066) );
in01f80 fopt783137 ( .a(n_44623), .o(n_44626) );
na02f80 g765574 ( .a(n_15103), .b(n_14465), .o(n_15402) );
na02f80 FE_RC_2305_0 ( .a(FE_RN_872_0), .b(n_25254), .o(FE_RN_873_0) );
na02f80 g772567 ( .a(n_8372), .b(n_8371), .o(n_8373) );
no02f80 g766366 ( .a(n_14177), .b(n_13469), .o(n_14333) );
in01f80 g761671 ( .a(n_20345), .o(n_20797) );
no02f80 g741601 ( .a(n_38587), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38604) );
na02f80 g772497 ( .a(n_8401), .b(n_8291), .o(n_8464) );
na02f80 g765523 ( .a(n_15565), .b(n_15865), .o(n_16018) );
ao22s80 g736306 ( .a(n_43855), .b(n_43394), .c(n_43854), .d(n_43395), .o(n_43887) );
in01f80 g752379 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_3_), .o(n_27823) );
na02f80 g762289 ( .a(n_18808), .b(n_18575), .o(n_19488) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_20_ ( .ck(newNet_2561), .d(n_27653), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_) );
no02f80 g743264 ( .a(n_36789), .b(n_36777), .o(n_36831) );
no02f80 g761658 ( .a(n_19489), .b(n_19488), .o(n_19490) );
oa12f80 g763620 ( .a(n_17470), .b(n_17469), .c(n_17262), .o(n_17502) );
in01f80 newInst_3470 ( .a(newNet_3469), .o(newNet_3470) );
in01f80 newInst_934 ( .a(newNet_933), .o(newNet_934) );
na02f80 g756193 ( .a(n_24164), .b(n_23733), .o(n_24200) );
in01f80 g743360 ( .a(n_36673), .o(n_36674) );
oa22f80 FE_RC_1410_0 ( .a(n_32180), .b(n_32214), .c(n_32181), .d(n_32215), .o(n_32263) );
na02f80 g775724 ( .a(n_5490), .b(n_3867), .o(n_5565) );
in01f80 newInst_3185 ( .a(newNet_3184), .o(newNet_3185) );
in01f80 g770244 ( .a(n_10914), .o(n_10923) );
in01f80 g768291 ( .a(n_12659), .o(n_12660) );
in01f80 FE_OCP_RBC2583_n_3734 ( .a(FE_OCP_RBN2579_n_3734), .o(FE_OCP_RBN2583_n_3734) );
no02f80 g774016 ( .a(n_6949), .b(n_6948), .o(n_6950) );
oa12f80 g778963 ( .a(n_1890), .b(FE_OCP_RBN2195_n_2103), .c(n_1856), .o(n_2160) );
no02f80 g775122 ( .a(n_5819), .b(n_5943), .o(n_5968) );
na02f80 g778316 ( .a(n_2874), .b(FE_OCP_RBN2460_n_2818), .o(n_2904) );
oa12f80 g772629 ( .a(n_8224), .b(n_8255), .c(n_8123), .o(n_8256) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_14_ ( .ck(newNet_1251), .d(n_5578), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_) );
oa12f80 g767721 ( .a(n_13101), .b(n_12823), .c(n_13086), .o(n_13087) );
no02f80 g775606 ( .a(n_5388), .b(n_5370), .o(n_5484) );
na02f80 g757621 ( .a(n_22584), .b(n_22314), .o(n_22639) );
oa12f80 g738458 ( .a(n_41443), .b(n_41397), .c(n_41405), .o(n_41551) );
in01f80 FE_RC_2041_0 ( .a(n_25542), .o(FE_RN_683_0) );
no02f80 g778063 ( .a(n_3626), .b(FE_OCP_RBN2294_n_2438), .o(n_2953) );
no02f80 g763894 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .o(n_17260) );
in01f80 g736467 ( .a(n_43728), .o(n_43729) );
na02f80 g765645 ( .a(n_15325), .b(n_14423), .o(n_15397) );
in01f80 newInst_2921 ( .a(newNet_2920), .o(newNet_2921) );
na02f80 g776548 ( .a(n_4432), .b(n_4419), .o(n_4420) );
oa12f80 g762704 ( .a(n_17917), .b(n_17875), .c(FE_OCP_RBN2144_FE_OCPN861_n_45450), .o(n_18018) );
in01f80 newInst_86 ( .a(newNet_85), .o(newNet_86) );
na02f80 g753330 ( .a(n_27057), .b(n_27068), .o(n_27056) );
na02f80 g773460 ( .a(n_7503), .b(n_7536), .o(n_7545) );
in01f80 newInst_591 ( .a(newNet_570), .o(newNet_591) );
na02f80 g755473 ( .a(n_24581), .b(n_24267), .o(n_24604) );
in01f80 fopt783446 ( .a(n_45012), .o(n_45050) );
in01f80 g763591 ( .a(n_17192), .o(n_17020) );
in01f80 g750748 ( .a(n_29265), .o(n_29266) );
na02f80 g760642 ( .a(n_19975), .b(n_19744), .o(n_19803) );
in01f80 FE_RC_2802_0 ( .a(n_38862), .o(FE_RN_1199_0) );
in01f80 g769958 ( .a(n_11072), .o(n_11073) );
in01f80 g746952 ( .a(n_33079), .o(n_33033) );
in01f80 newInst_555 ( .a(newNet_346), .o(newNet_555) );
in01f80 newInst_2009 ( .a(newNet_2008), .o(newNet_2009) );
in01f80 g758312 ( .a(n_22330), .o(n_22370) );
in01f80 g745863 ( .a(n_34219), .o(n_34193) );
in01f80 g778870 ( .a(FE_OCP_RBN2292_n_2438), .o(n_2741) );
in01f80 g778414 ( .a(n_2786), .o(n_2787) );
no02f80 g770151 ( .a(n_10770), .b(n_10768), .o(n_10769) );
oa22f80 g779089 ( .a(n_2042), .b(n_1804), .c(n_2024), .d(n_1805), .o(n_2086) );
in01f80 FE_OCP_RBC2559_n_44576 ( .a(FE_OCP_RBN2557_n_44576), .o(FE_OCP_RBN2559_n_44576) );
oa22f80 g784341 ( .a(FE_OFN774_n_46137), .b(n_6365), .c(n_46195), .d(n_6376), .o(n_46147) );
oa22f80 FE_RC_3962_0 ( .a(n_23760), .b(n_24224), .c(FE_OCPN1462_n_23759), .d(n_24225), .o(n_24305) );
in01f80 g748194 ( .a(n_31774), .o(n_31775) );
no02f80 g768010 ( .a(n_12634), .b(n_13412), .o(n_12682) );
no02f80 g740402 ( .a(FE_OCP_RBN3027_n_39942), .b(n_39932), .o(n_40032) );
na02f80 g776901 ( .a(n_3633), .b(n_2895), .o(n_3684) );
in01f80 g753308 ( .a(n_27291), .o(n_27292) );
in01f80 fopt783247 ( .a(n_36669), .o(n_44809) );
in01f80 g740084 ( .a(n_40038), .o(n_40068) );
in01f80 FE_OCPC1488_n_23447 ( .a(FE_OCPN1487_n_23447), .o(FE_OCPN1488_n_23447) );
na02f80 g766382 ( .a(n_14191), .b(n_14190), .o(n_14238) );
no02f80 g761097 ( .a(n_19087), .b(n_19115), .o(n_19206) );
na02f80 g756078 ( .a(n_24183), .b(n_23734), .o(n_24208) );
na02f80 g776567 ( .a(n_4283), .b(FE_OCP_RBN2692_FE_OCPN843_n_3912), .o(n_4447) );
na02f80 FE_RC_2176_0 ( .a(FE_RN_775_0), .b(n_26445), .o(FE_RN_776_0) );
in01f80 g752059 ( .a(n_28690), .o(n_28691) );
oa12f80 g757063 ( .a(n_23743), .b(n_23897), .c(n_23294), .o(n_23898) );
na02f80 g777149 ( .a(n_4873), .b(n_4852), .o(n_4874) );
in01f80 g752623 ( .a(n_27569), .o(n_27570) );
ao12f80 g746460 ( .a(n_34666), .b(n_34942), .c(n_34891), .o(n_34892) );
in01f80 newInst_1142 ( .a(newNet_1141), .o(newNet_1142) );
na02f80 g762325 ( .a(n_18072), .b(n_18109), .o(n_18128) );
in01f80 g749021 ( .a(n_31079), .o(n_31097) );
no02f80 g767934 ( .a(n_12635), .b(n_12658), .o(n_12705) );
in01f80 g765133 ( .a(n_15237), .o(n_15238) );
no02f80 g763387 ( .a(n_16919), .b(n_15939), .o(n_16957) );
na02f80 g769015 ( .a(n_11498), .b(n_11604), .o(n_11661) );
in01f80 newInst_1851 ( .a(newNet_320), .o(newNet_1851) );
in01f80 FE_OCP_RBC2851_n_46982 ( .a(FE_OCP_RBN2849_n_46982), .o(FE_OCP_RBN2851_n_46982) );
ao22s80 g737336 ( .a(n_42813), .b(n_42615), .c(n_42814), .d(n_42614), .o(n_42856) );
oa22f80 g779658 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .c(FE_OCPN946_n_1780), .d(n_1392), .o(n_1545) );
in01f80 newInst_857 ( .a(newNet_856), .o(newNet_857) );
no02f80 g751535 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_26_), .o(n_28673) );
oa12f80 g756797 ( .a(n_23045), .b(n_23379), .c(n_23378), .o(n_23380) );
in01f80 g741666 ( .a(n_38596), .o(n_38609) );
no02f80 g781305 ( .a(beta_31), .b(beta_16), .o(n_68) );
in01f80 g763901 ( .a(n_17106), .o(n_17056) );
ao12f80 g738047 ( .a(n_42134), .b(n_42133), .c(n_42132), .o(n_42148) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_6_ ( .ck(newNet_3583), .d(n_15751), .o(delay_add_ln22_unr11_stage5_stallmux_q_6_) );
na02f80 g740837 ( .a(n_39434), .b(n_39433), .o(n_39435) );
no02f80 g745816 ( .a(n_44102), .b(n_33580), .o(n_34162) );
no02f80 g752652 ( .a(n_28159), .b(n_27987), .o(n_28242) );
na02f80 g779159 ( .a(n_2606), .b(FE_OFN810_n_1941), .o(n_1942) );
na02f80 FE_RC_147_0 ( .a(FE_RN_44_0), .b(n_12040), .o(n_12232) );
no02f80 g742765 ( .a(n_37291), .b(n_37214), .o(n_37302) );
in01f80 g753322 ( .a(n_27101), .o(n_27102) );
in01f80 g747474 ( .a(n_32433), .o(n_32602) );
na02f80 g761875 ( .a(n_18915), .b(n_18914), .o(n_18936) );
na02f80 g756575 ( .a(n_23574), .b(n_22562), .o(n_23608) );
in01f80 g760148 ( .a(n_20665), .o(n_20666) );
no02f80 g764394 ( .a(n_16128), .b(n_16094), .o(n_16230) );
in01f80 g756397 ( .a(n_24277), .o(n_24330) );
in01f80 g749491 ( .a(n_30453), .o(n_30454) );
no02f80 g741492 ( .a(n_38775), .b(n_38774), .o(n_38776) );
in01f80 g747786 ( .a(n_32111), .o(n_32112) );
no02f80 g751340 ( .a(n_29460), .b(n_29459), .o(n_29461) );
na02f80 g740607 ( .a(n_39633), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39678) );
na02f80 FE_RC_2197_0 ( .a(FE_RN_788_0), .b(n_26100), .o(n_26140) );
na02f80 g781234 ( .a(n_101), .b(n_38), .o(n_80) );
na02f80 g770673 ( .a(n_10109), .b(n_44463), .o(n_10313) );
na02f80 g772995 ( .a(n_7803), .b(n_7786), .o(n_7787) );
in01f80 g757377 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .o(n_22873) );
in01f80 g736564 ( .a(n_43651), .o(n_43659) );
no02f80 g749446 ( .a(n_30558), .b(n_45744), .o(n_30562) );
no02f80 g748517 ( .a(n_32675), .b(n_32606), .o(n_32748) );
in01f80 g760108 ( .a(n_20374), .o(n_20407) );
in01f80 g740392 ( .a(n_40242), .o(n_40243) );
in01f80 g739165 ( .a(n_40992), .o(n_40990) );
in01f80 g750966 ( .a(n_30185), .o(n_30186) );
na02f80 g766266 ( .a(n_14249), .b(n_13437), .o(n_14250) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_16_ ( .ck(newNet_578), .d(n_17750), .o(delay_xor_ln22_unr12_stage5_stallmux_q_16_) );
in01f80 newInst_67 ( .a(newNet_66), .o(newNet_67) );
no02f80 g749140 ( .a(n_30862), .b(n_30832), .o(n_30833) );
na02f80 g736987 ( .a(n_43120), .b(n_42997), .o(n_43400) );
in01f80 newInst_3106 ( .a(newNet_888), .o(newNet_3106) );
no02f80 g744592 ( .a(n_36621), .b(n_36284), .o(n_36662) );
in01f80 FE_OCP_RBC2876_n_10354 ( .a(n_10354), .o(FE_OCP_RBN2876_n_10354) );
na02f80 g774184 ( .a(n_6656), .b(n_6619), .o(n_6635) );
in01f80 newInst_2305 ( .a(newNet_2304), .o(newNet_2305) );
no03m80 g748002 ( .a(n_44042), .b(n_33006), .c(n_32406), .o(n_33125) );
na02f80 g772012 ( .a(FE_OFN754_n_44461), .b(n_9381), .o(n_9431) );
in01f80 g761144 ( .a(n_19201), .o(n_19202) );
in01f80 FE_RC_3597_0 ( .a(n_13272), .o(FE_RN_1571_0) );
in01f80 g756532 ( .a(n_24048), .o(n_24049) );
na02f80 g770955 ( .a(FE_OCP_RBN3634_n_47260), .b(n_9985), .o(n_9987) );
in01f80 g744954 ( .a(FE_OCP_RBN2645_n_34980), .o(n_35023) );
na02f80 g780479 ( .a(n_1002), .b(n_736), .o(n_763) );
na02f80 g768641 ( .a(n_12106), .b(n_12105), .o(n_12107) );
na02f80 g751800 ( .a(n_28911), .b(n_28909), .o(n_28910) );
na02f80 g761863 ( .a(n_18343), .b(n_18301), .o(n_18374) );
no02f80 g758275 ( .a(n_22288), .b(FE_OCP_RBN1716_n_20734), .o(n_22554) );
in01f80 g753088 ( .a(n_27267), .o(n_27268) );
na02f80 g749879 ( .a(n_29902), .b(n_29968), .o(n_29969) );
na02f80 g766281 ( .a(n_14241), .b(n_14091), .o(n_14336) );
na02f80 g749515 ( .a(n_31857), .b(n_31351), .o(n_31939) );
in01f80 FE_OCP_RBC3473_n_7886 ( .a(FE_OCP_RBN3470_n_7886), .o(FE_OCP_RBN3473_n_7886) );
in01f80 fopt783175 ( .a(n_35221), .o(n_44713) );
na02f80 FE_RC_2490_0 ( .a(FE_RN_1006_0), .b(FE_RN_1007_0), .o(FE_RN_1008_0) );
na02f80 g747152 ( .a(n_32856), .b(n_32855), .o(n_32870) );
na02f80 g758848 ( .a(n_21475), .b(n_45081), .o(n_21506) );
in01f80 FE_OCP_RBC2006_n_45209 ( .a(n_45209), .o(FE_OCP_RBN2006_n_45209) );
in01f80 g736920 ( .a(n_43023), .o(n_43024) );
in01f80 g784704 ( .a(n_6749), .o(n_47177) );
na02f80 g763892 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_24_), .o(n_17353) );
oa12f80 g763618 ( .a(n_17430), .b(n_17208), .c(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17471) );
na02f80 g737422 ( .a(n_42733), .b(n_42749), .o(n_42802) );
in01f80 g762779 ( .a(n_17825), .o(n_17802) );
no02f80 g763821 ( .a(n_17309), .b(n_17304), .o(n_17356) );
no02f80 g741322 ( .a(FE_OCP_RBN3582_n_44944), .b(n_38598), .o(n_39149) );
na02f80 g766922 ( .a(n_13864), .b(n_13863), .o(n_13865) );
in01f80 g751807 ( .a(n_28268), .o(n_28301) );
na02f80 g758145 ( .a(n_22330), .b(n_22293), .o(n_22413) );
in01f80 g751166 ( .a(n_29943), .o(n_30037) );
in01f80 newInst_3403 ( .a(newNet_3402), .o(newNet_3403) );
na02f80 g766495 ( .a(n_14494), .b(n_14493), .o(n_14495) );
na02f80 g781033 ( .a(sin_out_0), .b(FE_OFN5_n_43918), .o(n_334) );
oa12f80 g778209 ( .a(n_2123), .b(FE_OCP_RBN2322_n_2638), .c(n_2097), .o(n_2747) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_13_ ( .ck(newNet_2878), .d(n_11098), .o(delay_add_ln22_unr8_stage4_stallmux_q_13_) );
in01f80 g748913 ( .a(n_32408), .o(n_32490) );
in01f80 newInst_3428 ( .a(newNet_3422), .o(newNet_3428) );
na02f80 g777926 ( .a(n_3132), .b(n_3145), .o(n_3214) );
na02f80 g745239 ( .a(n_35853), .b(n_35795), .o(n_36419) );
na02f80 g745425 ( .a(FE_OCP_RBN2993_n_35539), .b(n_35675), .o(n_35717) );
in01f80 g776734 ( .a(n_3963), .o(n_3964) );
no02f80 g773527 ( .a(n_7440), .b(delay_add_ln22_unr5_stage3_stallmux_q_22_), .o(n_8405) );
no03m80 g743810 ( .a(n_37224), .b(n_37191), .c(n_37167), .o(n_37225) );
no02f80 g772048 ( .a(n_8824), .b(n_8772), .o(n_8773) );
na02f80 g762426 ( .a(n_18089), .b(n_18073), .o(n_18163) );
no02f80 g775974 ( .a(n_5325), .b(n_5227), .o(n_5481) );
in01f80 newInst_377 ( .a(newNet_376), .o(newNet_377) );
na02f80 g780167 ( .a(n_1170), .b(n_797), .o(n_1147) );
na02f80 g779748 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .o(n_1527) );
in01f80 FE_OCPC1016_n_23307 ( .a(n_23307), .o(FE_OCPN1016_n_23307) );
no02f80 g759453 ( .a(FE_OCP_RBN1727_FE_RN_1583_0), .b(n_20774), .o(n_20823) );
na02f80 g763271 ( .a(n_17233), .b(n_17134), .o(n_17234) );
no02f80 g736577 ( .a(n_43528), .b(n_43224), .o(n_43567) );
na02f80 g738993 ( .a(n_41149), .b(n_40910), .o(n_41154) );
in01f80 g772891 ( .a(n_7798), .o(n_7821) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_2_ ( .ck(newNet_1583), .d(n_26996), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_2_) );
in01f80 drc ( .a(n_45809), .o(n_45812) );
na02f80 g778743 ( .a(n_2207), .b(n_2006), .o(n_2303) );
in01f80 g766919 ( .a(n_13906), .o(n_13976) );
no02f80 g765494 ( .a(FE_OFN764_n_15670), .b(n_15833), .o(n_15829) );
no02f80 g737029 ( .a(n_43020), .b(n_43019), .o(n_43033) );
na02f80 g773531 ( .a(n_7507), .b(n_7505), .o(n_7506) );
oa12f80 g756224 ( .a(n_24771), .b(n_24770), .c(n_24769), .o(n_25124) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_0_ ( .ck(newNet_894), .d(n_32289), .o(delay_xor_ln21_unr21_stage8_stallmux_q_0_) );
na02f80 g766933 ( .a(n_13863), .b(n_13822), .o(n_14010) );
in01f80 g768712 ( .a(n_12134), .o(n_12135) );
na02f80 FE_RC_1955_0 ( .a(n_19218), .b(n_19219), .o(FE_RN_629_0) );
in01f80 g737657 ( .a(n_42756), .o(n_42757) );
in01f80 g742565 ( .a(n_37581), .o(n_37575) );
oa22f80 FE_RC_38_0 ( .a(FE_OFN806_n_46196), .b(FE_OCP_RBN3124_n_6557), .c(FE_OFN84_n_46137), .d(n_6557), .o(n_46185) );
na02f80 g742003 ( .a(n_38316), .b(n_38256), .o(n_38362) );
in01f80 newInst_1343 ( .a(newNet_1342), .o(newNet_1343) );
na02f80 g775044 ( .a(n_6012), .b(n_6086), .o(n_6114) );
oa22f80 g772274 ( .a(n_8630), .b(n_8685), .c(n_8629), .d(n_8647), .o(n_8809) );
no02f80 g763168 ( .a(n_17288), .b(n_17118), .o(n_17404) );
in01f80 g770117 ( .a(n_10833), .o(n_10806) );
na02f80 g771774 ( .a(n_9035), .b(FE_OCP_RBN3548_n_44575), .o(n_9229) );
in01f80 fopt782966 ( .a(n_44429), .o(n_44428) );
na02f80 g755832 ( .a(n_25004), .b(n_24994), .o(n_25112) );
ao12f80 g750790 ( .a(n_29379), .b(n_29115), .c(n_29033), .o(n_29192) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_14_ ( .ck(newNet_1539), .d(n_32064), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_) );
no02f80 g770470 ( .a(n_10559), .b(FE_OCP_RBN3592_n_8902), .o(n_10584) );
in01f80 FE_OCP_RBC2229_n_7598 ( .a(FE_OCP_RBN2228_n_7598), .o(FE_OCP_RBN2229_n_7598) );
oa22f80 FE_RC_158_0 ( .a(n_17382), .b(n_17689), .c(n_17383), .d(n_45205), .o(n_17834) );
no02f80 g736447 ( .a(n_43768), .b(n_43524), .o(n_43822) );
na02f80 g768792 ( .a(n_11956), .b(n_11955), .o(n_11994) );
no02f80 g743469 ( .a(n_36515), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36538) );
in01f80 g769315 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .o(n_11528) );
na03f80 FE_RC_638_0 ( .a(n_6889), .b(FE_RN_200_0), .c(n_6634), .o(n_6980) );
na02f80 g749771 ( .a(n_31287), .b(n_31285), .o(n_31286) );
in01f80 g772346 ( .a(n_8434), .o(n_8435) );
ao12f80 g774271 ( .a(n_6425), .b(n_6491), .c(n_6362), .o(n_6565) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_23_ ( .ck(newNet_2846), .d(n_11873), .o(delay_add_ln22_unr8_stage4_stallmux_q_23_) );
na02f80 g779082 ( .a(n_2035), .b(delay_add_ln22_unr2_stage2_stallmux_q_14_), .o(n_2085) );
na02f80 g749714 ( .a(n_31325), .b(n_31374), .o(n_31395) );
in01f80 FE_RC_1600_0 ( .a(n_27432), .o(FE_RN_448_0) );
in01f80 g770900 ( .a(n_9807), .o(n_9808) );
na02f80 g766027 ( .a(n_14687), .b(n_14719), .o(n_14720) );
in01f80 newInst_1792 ( .a(newNet_1390), .o(newNet_1792) );
oa12f80 g760195 ( .a(n_20896), .b(n_20834), .c(n_20055), .o(n_20897) );
na02f80 g750827 ( .a(n_29210), .b(n_29094), .o(n_29258) );
in01f80 newInst_1254 ( .a(newNet_376), .o(newNet_1254) );
in01f80 FE_OCP_RBC1173_n_13858 ( .a(FE_OCP_RBN2353_n_13858), .o(FE_OCP_RBN1173_n_13858) );
no02f80 g765363 ( .a(n_15447), .b(n_14082), .o(n_15569) );
in01f80 g765113 ( .a(n_15163), .o(n_15164) );
no02f80 g743699 ( .a(n_36346), .b(n_36331), .o(n_36376) );
na02f80 g766436 ( .a(n_14621), .b(n_14620), .o(n_14622) );
in01f80 g769956 ( .a(n_10946), .o(n_10947) );
in01f80 g745163 ( .a(n_36252), .o(n_36253) );
ao12f80 g783820 ( .a(n_2424), .b(n_2575), .c(n_2349), .o(n_45505) );
ao12f80 g752727 ( .a(n_44046), .b(n_27814), .c(n_27899), .o(n_28054) );
no02f80 g755884 ( .a(n_25055), .b(n_25083), .o(n_25084) );
na02f80 g784594 ( .a(n_38453), .b(n_38486), .o(n_46417) );
na02f80 g779273 ( .a(n_1736), .b(n_1559), .o(n_1755) );
oa12f80 g744531 ( .a(n_35398), .b(n_35397), .c(n_35396), .o(n_35419) );
na02f80 g744935 ( .a(n_34903), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34936) );
in01f80 g770198 ( .a(n_10676), .o(n_11502) );
in01f80 g742124 ( .a(n_37906), .o(n_37941) );
na02f80 g745793 ( .a(n_44102), .b(FE_OCP_RBN2323_n_33942), .o(n_34303) );
no02f80 g765303 ( .a(n_15826), .b(n_15834), .o(n_15871) );
no02f80 g743118 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n_37091) );
na02f80 g763616 ( .a(n_16758), .b(n_16832), .o(n_16864) );
in01f80 newInst_2523 ( .a(newNet_1033), .o(newNet_2523) );
oa22f80 FE_RC_782_0 ( .a(FE_OFN803_n_46285), .b(n_12212), .c(FE_OFN771_n_46337), .d(n_12194), .o(n_46345) );
in01f80 g763077 ( .a(n_17617), .o(n_17618) );
in01f80 g738231 ( .a(n_41939), .o(n_41977) );
in01f80 g761176 ( .a(n_19064), .o(n_19641) );
ao12f80 g747201 ( .a(n_33796), .b(n_33795), .c(n_33794), .o(n_34585) );
na02f80 g749791 ( .a(FE_OCP_RBN3010_n_31117), .b(n_31281), .o(n_31393) );
no02f80 FE_RC_2527_0 ( .a(FE_RN_1029_0), .b(FE_RN_1030_0), .o(FE_RN_1031_0) );
in01f80 FE_RC_3623_0 ( .a(FE_RN_1587_0), .o(n_20890) );
na02f80 g750614 ( .a(FE_OCP_RBN1690_n_29491), .b(n_28350), .o(n_29633) );
no02f80 g780778 ( .a(n_455), .b(n_454), .o(n_540) );
no02f80 g758321 ( .a(FE_OCPN991_n_22249), .b(n_21393), .o(n_22366) );
in01f80 FE_RC_176_0 ( .a(beta_0), .o(FE_RN_55_0) );
na02f80 g759014 ( .a(n_22011), .b(n_21995), .o(n_21996) );
ao12f80 g754962 ( .a(n_25804), .b(n_25803), .c(n_25802), .o(n_26605) );
in01f80 g767888 ( .a(n_12865), .o(n_12754) );
na02f80 FE_RC_2818_0 ( .a(n_34343), .b(n_34344), .o(FE_RN_1207_0) );
in01f80 newInst_3041 ( .a(newNet_3040), .o(newNet_3041) );
in01f80 FE_OCP_RBC3616_n_20249 ( .a(FE_OCP_RBN2670_n_20249), .o(FE_OCP_RBN3616_n_20249) );
na02f80 g751446 ( .a(n_28632), .b(n_28548), .o(n_28576) );
in01f80 g772241 ( .a(n_8856), .o(n_8893) );
in01f80 g763732 ( .a(n_17536), .o(n_17604) );
na02f80 g751491 ( .a(n_29177), .b(n_29201), .o(n_29255) );
in01f80 g751605 ( .a(n_28463), .o(n_28464) );
na02f80 g739205 ( .a(n_40869), .b(n_40790), .o(n_40791) );
no02f80 g764964 ( .a(n_15423), .b(n_15469), .o(n_15542) );
na02f80 g738423 ( .a(n_41694), .b(n_41699), .o(n_42001) );
ao12f80 g738872 ( .a(n_41305), .b(n_41304), .c(n_41303), .o(n_41634) );
no02f80 g742589 ( .a(n_37432), .b(n_37431), .o(n_37433) );
no02f80 g742375 ( .a(n_37809), .b(n_37808), .o(n_37845) );
no02f80 g750017 ( .a(n_30198), .b(n_30212), .o(n_30273) );
in01f80 FE_OCP_RBC3365_n_44722 ( .a(FE_OCP_RBN3306_n_44722), .o(FE_OCP_RBN3365_n_44722) );
no02f80 g738360 ( .a(n_41733), .b(n_41692), .o(n_41734) );
na02f80 g772354 ( .a(n_8717), .b(n_8716), .o(n_8718) );
in01f80 g761475 ( .a(n_19903), .o(n_19871) );
na02f80 g748429 ( .a(n_31476), .b(n_31655), .o(n_31681) );
no02f80 g772022 ( .a(FE_OCPN903_n_44581), .b(n_9220), .o(n_9309) );
in01f80 g750134 ( .a(n_29890), .o(n_29916) );
na02f80 g775736 ( .a(n_5549), .b(n_47013), .o(n_5727) );
no02f80 g761187 ( .a(n_18986), .b(n_17732), .o(n_19017) );
oa22f80 FE_RC_3152_0 ( .a(FE_RN_761_0), .b(n_15231), .c(n_15175), .d(FE_OCP_RBN2825_n_15231), .o(n_15459) );
na02f80 g776916 ( .a(n_3897), .b(n_3980), .o(n_4064) );
oa12f80 g772738 ( .a(n_7830), .b(n_8169), .c(n_7740), .o(n_8480) );
na02f80 g776661 ( .a(n_3860), .b(n_2982), .o(n_4131) );
in01f80 newInst_1155 ( .a(newNet_1154), .o(newNet_1155) );
no02f80 g774343 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .o(n_7029) );
na02f80 g771231 ( .a(n_9794), .b(n_9737), .o(n_9738) );
oa12f80 g750492 ( .a(n_29544), .b(n_29543), .c(n_29542), .o(n_31125) );
no02f80 g750994 ( .a(n_28918), .b(n_28576), .o(n_28963) );
no02f80 g749142 ( .a(FE_OCP_RBN2888_n_46957), .b(n_30759), .o(n_31943) );
in01f80 g776143 ( .a(n_5114), .o(n_5115) );
in01f80 g748099 ( .a(n_33310), .o(n_33316) );
na02f80 g741263 ( .a(FE_OCP_RBN2550_n_44944), .b(n_38436), .o(n_39271) );
in01f80 g762951 ( .a(n_17687), .o(n_17649) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_19_ ( .ck(newNet_1237), .d(n_5915), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_) );
in01f80 FE_OCP_DRV_C1569_n_29777 ( .a(n_29777), .o(FE_OCP_DRV_N1569_n_29777) );
in01f80 g778710 ( .a(n_2389), .o(n_2448) );
oa12f80 g762934 ( .a(n_17619), .b(n_17678), .c(n_17548), .o(n_17771) );
no02f80 g773874 ( .a(n_7052), .b(n_6880), .o(n_7073) );
ao22s80 g780853 ( .a(n_521), .b(n_476), .c(n_420), .d(n_261), .o(n_621) );
no02f80 g742235 ( .a(FE_OCP_RBN3425_n_44881), .b(n_37654), .o(n_38131) );
na02f80 g763708 ( .a(n_16733), .b(n_16778), .o(n_16998) );
oa22f80 g763967 ( .a(n_16889), .b(n_16064), .c(n_16890), .d(n_16063), .o(n_17017) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_26_ ( .ck(newNet_1597), .d(n_27574), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_) );
na02f80 g748120 ( .a(n_31948), .b(n_31930), .o(n_31970) );
no02f80 g746624 ( .a(n_34473), .b(n_34523), .o(n_34544) );
no02f80 g769575 ( .a(n_11335), .b(n_11353), .o(n_11379) );
no02f80 g784762 ( .a(FE_OCP_RBN2203_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n_47248) );
in01f80 newInst_2393 ( .a(newNet_785), .o(newNet_2393) );
na02f80 FE_RC_2756_0 ( .a(FE_RN_1171_0), .b(FE_RN_1172_0), .o(n_2938) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_14_ ( .ck(newNet_972), .d(n_22962), .o(delay_xor_ln21_unr15_stage6_stallmux_q_14_) );
oa12f80 g771635 ( .a(n_9430), .b(n_9482), .c(n_9429), .o(n_9518) );
in01f80 FE_OCPC1236_n_32791 ( .a(FE_OCPN1235_n_32791), .o(FE_OCPN1236_n_32791) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_13_ ( .ck(newNet_3168), .d(n_40459), .o(delay_add_ln22_unr27_stage10_stallmux_q_13_) );
no02f80 g776349 ( .a(n_4347), .b(n_3106), .o(n_4568) );
no02f80 g738911 ( .a(n_41265), .b(n_41251), .o(n_41298) );
in01f80 g747154 ( .a(n_32925), .o(n_32926) );
in01f80 FE_OCP_RBC2713_n_14982 ( .a(n_14982), .o(FE_OCP_RBN2713_n_14982) );
na02f80 FE_RC_4256_0 ( .a(n_21283), .b(n_22294), .o(FE_RN_1874_0) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_17_ ( .ck(newNet_1756), .d(n_22362), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_7_ ( .ck(newNet_2435), .d(n_31673), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_) );
in01f80 g745849 ( .a(n_34157), .o(n_34158) );
na02f80 g752535 ( .a(n_27600), .b(n_27551), .o(n_27639) );
no02f80 g769226 ( .a(n_11627), .b(n_45301), .o(n_11628) );
in01f80 g736529 ( .a(n_43699), .o(n_43700) );
na02f80 g769723 ( .a(n_11172), .b(n_11159), .o(n_11225) );
no02f80 g780935 ( .a(n_420), .b(n_240), .o(n_433) );
na02f80 g767283 ( .a(n_13541), .b(n_13540), .o(n_13542) );
ao22s80 FE_RC_1591_0 ( .a(n_2218), .b(n_2293), .c(n_2622), .d(n_2245), .o(n_2342) );
oa22f80 g745785 ( .a(n_44102), .b(n_34200), .c(n_44112), .d(n_33686), .o(n_34716) );
na02f80 g775538 ( .a(n_5581), .b(n_5451), .o(n_5465) );
na02f80 g748926 ( .a(n_30967), .b(n_30913), .o(n_31061) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_13_ ( .ck(newNet_3444), .d(n_27360), .o(delay_add_ln22_unr17_stage7_stallmux_q_13_) );
in01f80 g742516 ( .a(n_37604), .o(n_37605) );
ao12f80 g769876 ( .a(n_10903), .b(n_11032), .c(n_10872), .o(n_11129) );
in01f80 FE_RC_1401_0 ( .a(FE_RN_410_0), .o(n_45331) );
in01f80 FE_OCP_RBC2430_n_14018 ( .a(n_14018), .o(FE_OCP_RBN2430_n_14018) );
in01f80 FE_OCP_RBC3658_n_15314 ( .a(FE_OCP_RBN3657_n_15314), .o(FE_OCP_RBN3658_n_15314) );
in01f80 g765014 ( .a(n_16263), .o(n_16264) );
in01f80 FE_OCP_RBC3286_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3286_n_44365) );
no02f80 g777213 ( .a(n_3612), .b(n_3567), .o(n_3755) );
no02f80 g742105 ( .a(n_37886), .b(n_37883), .o(n_37943) );
oa22f80 g743779 ( .a(n_36324), .b(n_36320), .c(n_36073), .d(n_36321), .o(n_36388) );
in01f80 FE_OCP_RBC2603_n_39126 ( .a(n_39126), .o(FE_OCP_RBN2603_n_39126) );
na02f80 g766183 ( .a(n_14544), .b(n_14543), .o(n_14573) );
na02f80 g756083 ( .a(n_24904), .b(n_24903), .o(n_24905) );
no02f80 g779620 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_21_), .o(n_1990) );
na02f80 g758980 ( .a(n_21195), .b(n_21191), .o(n_21332) );
in01f80 FE_OCPC1049_n_4459 ( .a(n_4459), .o(FE_OCPN1049_n_4459) );
na02f80 g750462 ( .a(n_29500), .b(n_25738), .o(n_29596) );
no02f80 g737696 ( .a(n_42216), .b(n_41916), .o(n_42260) );
na02f80 FE_RC_813_0 ( .a(FE_RN_243_0), .b(FE_RN_244_0), .o(FE_RN_245_0) );
in01f80 g747611 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_), .o(n_32381) );
no02f80 g737575 ( .a(n_42288), .b(n_42260), .o(n_42289) );
in01f80 g738936 ( .a(n_41290), .o(n_41291) );
no02f80 g779538 ( .a(n_1553), .b(n_1603), .o(n_1884) );
in01f80 g763774 ( .a(n_17365), .o(n_17366) );
oa22f80 g744668 ( .a(n_35262), .b(FE_OCPN1434_n_30614), .c(n_35281), .d(n_30633), .o(n_35340) );
oa12f80 g746745 ( .a(n_34170), .b(n_34169), .c(n_34168), .o(n_34227) );
no03m80 FE_RC_1530_0 ( .a(n_27929), .b(n_28280), .c(n_28298), .o(n_28328) );
na02f80 g773152 ( .a(FE_OCPN940_n_7712), .b(n_7812), .o(n_7824) );
in01f80 newInst_2555 ( .a(newNet_1444), .o(newNet_2555) );
na02f80 g746556 ( .a(n_34638), .b(n_34606), .o(n_34639) );
in01f80 g763803 ( .a(n_17358), .o(n_17468) );
no02f80 g742081 ( .a(FE_OCP_RBN3445_n_37945), .b(n_38279), .o(n_38311) );
na02f80 g767309 ( .a(n_13496), .b(n_13495), .o(n_13538) );
in01f80 g759794 ( .a(n_20417), .o(n_20418) );
in01f80 FE_OCP_RBC2718_n_9182 ( .a(n_9182), .o(FE_OCP_RBN2718_n_9182) );
oa12f80 g744712 ( .a(n_36122), .b(n_36494), .c(n_35848), .o(n_36571) );
na02f80 g763296 ( .a(n_17037), .b(n_17135), .o(n_17136) );
no02f80 g740149 ( .a(n_39816), .b(n_39506), .o(n_39921) );
in01f80 g769313 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_20_), .o(n_12693) );
na02f80 g777169 ( .a(n_4201), .b(n_4193), .o(n_4695) );
no02f80 g746916 ( .a(FE_OCP_RBN3385_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_20_), .o(n_33151) );
na02f80 g738688 ( .a(n_41716), .b(n_41340), .o(n_41717) );
ao12f80 g757310 ( .a(n_23131), .b(n_44068), .c(delay_xor_ln21_unr15_stage6_stallmux_q_15_), .o(n_23165) );
na02f80 g742176 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37620), .o(n_38306) );
in01f80 g773250 ( .a(n_7631), .o(n_7632) );
na02f80 g748796 ( .a(n_32407), .b(n_32357), .o(n_32453) );
in01f80 g744625 ( .a(n_36638), .o(n_36639) );
in01f80 g763499 ( .a(n_16904), .o(n_16905) );
oa22f80 FE_RC_1289_0 ( .a(n_38778), .b(n_38681), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .d(n_38655), .o(n_38693) );
in01f80 g770469 ( .a(n_10584), .o(n_10653) );
in01f80 newInst_2226 ( .a(newNet_2225), .o(newNet_2226) );
no02f80 g771258 ( .a(n_9353), .b(FE_OCP_RBN2564_FE_RN_1125_0), .o(n_9489) );
no02f80 g757674 ( .a(n_22542), .b(n_22273), .o(n_22601) );
no02f80 g776438 ( .a(n_4103), .b(n_4007), .o(n_4161) );
in01f80 FE_OCPUNCOC3146_n_21058 ( .a(FE_OCPUNCON3145_n_21058), .o(FE_OCPUNCON3146_n_21058) );
na02f80 g770106 ( .a(n_10807), .b(n_10782), .o(n_10922) );
in01f80 FE_OFC507_n_25938 ( .a(FE_OFN792_n_25938), .o(FE_OFN507_n_25938) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_13_ ( .ck(newNet_516), .d(n_22834), .o(delay_xor_ln22_unr15_stage6_stallmux_q_13_) );
na02f80 g742832 ( .a(n_37268), .b(n_37271), .o(n_37311) );
in01f80 g744210 ( .a(n_36238), .o(n_36239) );
na02f80 g757211 ( .a(n_23193), .b(n_23192), .o(n_23249) );
in01f80 g761163 ( .a(n_19140), .o(n_19141) );
ms00f80 sin_out_reg_1_ ( .ck(newNet_60), .d(n_43237), .o(sin_out_1) );
in01f80 g768869 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n_11886) );
no02f80 g740359 ( .a(n_39741), .b(n_39740), .o(n_39772) );
na02f80 g770875 ( .a(n_9852), .b(n_44819), .o(n_9932) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_20_ ( .ck(newNet_2656), .d(n_22635), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_) );
na02f80 g770628 ( .a(n_10423), .b(n_10350), .o(n_10560) );
oa12f80 g760759 ( .a(n_19465), .b(n_19602), .c(n_19532), .o(n_19719) );
na02f80 g746093 ( .a(n_35109), .b(n_34634), .o(n_35191) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_18_ ( .ck(newNet_178), .d(n_46344), .o(delay_xor_ln22_unr9_stage4_stallmux_q_18_) );
no02f80 g778177 ( .a(n_2727), .b(n_2526), .o(n_2783) );
na02f80 g766891 ( .a(n_14259), .b(n_14758), .o(n_14381) );
no02f80 g780707 ( .a(n_634), .b(n_475), .o(n_635) );
in01f80 g746356 ( .a(n_33523), .o(n_33616) );
in01f80 newInst_3346 ( .a(newNet_2677), .o(newNet_3346) );
in01f80 newInst_2415 ( .a(newNet_2414), .o(newNet_2415) );
ao12f80 g747764 ( .a(n_33950), .b(n_33372), .c(n_33626), .o(n_34103) );
no02f80 g753761 ( .a(FE_OCP_RBN3694_n_26409), .b(n_26407), .o(n_26500) );
na02f80 g750719 ( .a(n_29198), .b(n_29219), .o(n_29298) );
in01f80 g753632 ( .a(n_27321), .o(n_27322) );
oa22f80 g746501 ( .a(n_33306), .b(n_33101), .c(n_33272), .d(n_33100), .o(n_33341) );
na02f80 g743871 ( .a(n_35671), .b(n_35670), .o(n_35672) );
oa12f80 g780122 ( .a(n_1161), .b(n_1160), .c(n_1159), .o(n_1188) );
no02f80 g739795 ( .a(n_40467), .b(n_40499), .o(n_40500) );
ao22s80 g742959 ( .a(n_36995), .b(n_36913), .c(n_36921), .d(n_36912), .o(n_37741) );
in01f80 g746475 ( .a(n_35809), .o(n_34671) );
oa12f80 g755363 ( .a(n_25031), .b(n_25494), .c(n_25436), .o(n_25577) );
in01f80 newInst_2211 ( .a(newNet_2210), .o(newNet_2211) );
na02f80 g749524 ( .a(n_30498), .b(n_30071), .o(n_30530) );
no02f80 g771684 ( .a(n_9169), .b(n_9168), .o(n_9238) );
na02f80 g753569 ( .a(n_26698), .b(n_26672), .o(n_26802) );
na02f80 g773763 ( .a(n_7201), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_), .o(n_7234) );
in01f80 FE_RC_2375_0 ( .a(n_12278), .o(FE_RN_923_0) );
in01f80 g739599 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_1_), .o(n_40604) );
in01f80 g743390 ( .a(n_36748), .o(n_36749) );
oa22f80 FE_RC_3877_0 ( .a(n_23963), .b(FE_OCP_RBN2417_n_24720), .c(n_23962), .d(n_24720), .o(n_24857) );
in01f80 g737060 ( .a(n_43125), .o(n_43166) );
na02f80 g776925 ( .a(n_4014), .b(n_3938), .o(n_4172) );
na02f80 g742927 ( .a(n_44038), .b(n_44037), .o(n_37115) );
in01f80 g746852 ( .a(n_33017), .o(n_33018) );
na02f80 g750986 ( .a(n_30100), .b(n_30036), .o(n_30811) );
in01f80 FE_OCP_RBC3433_n_33664 ( .a(FE_OCP_RBN3432_n_33664), .o(FE_OCP_RBN3433_n_33664) );
in01f80 g770753 ( .a(n_9896), .o(n_9897) );
in01f80 FE_RC_32_0 ( .a(n_6081), .o(FE_RN_6_0) );
oa22f80 g770782 ( .a(n_9859), .b(FE_OCP_RBN3597_FE_OCPN1243_n_44460), .c(FE_OCP_RBN2783_n_9859), .d(FE_RN_1433_0), .o(n_10057) );
na02f80 g753424 ( .a(n_26967), .b(n_26966), .o(n_27026) );
no02f80 g760818 ( .a(n_19533), .b(FE_OCP_RBN1838_n_19528), .o(n_19617) );
na03f80 FE_RC_576_0 ( .a(n_23515), .b(n_23500), .c(n_23104), .o(n_23516) );
na02f80 g742386 ( .a(n_37780), .b(FE_OCP_RBN2187_n_37686), .o(n_37781) );
in01f80 g767484 ( .a(FE_OCP_RBN3430_n_13245), .o(n_14555) );
no02f80 g749855 ( .a(FE_OCP_RBN3016_n_31117), .b(n_31253), .o(n_31321) );
in01f80 FE_OCP_RBC2218_FE_OCPN950_n_28595 ( .a(FE_OCP_RBN2217_FE_OCPN950_n_28595), .o(FE_OCP_RBN2218_FE_OCPN950_n_28595) );
ao22s80 FE_RC_3958_0 ( .a(n_28572), .b(n_28951), .c(n_28573), .d(n_28950), .o(n_29033) );
in01f80 g766220 ( .a(n_14379), .o(n_14416) );
ao12f80 g738966 ( .a(n_40996), .b(n_41155), .c(n_40872), .o(n_41213) );
oa12f80 g739708 ( .a(n_40338), .b(n_40505), .c(n_40117), .o(n_40519) );
in01f80 g761484 ( .a(n_19676), .o(n_19731) );
no03m80 FE_RC_1175_0 ( .a(n_2448), .b(n_2435), .c(n_2390), .o(n_2510) );
in01f80 FE_OFC627_n_34445 ( .a(FE_OFN626_n_34445), .o(FE_OFN627_n_34445) );
na02f80 g780832 ( .a(n_415), .b(n_438), .o(n_593) );
no02f80 g777811 ( .a(n_3362), .b(n_3361), .o(n_3556) );
in01f80 g778937 ( .a(n_2898), .o(n_2206) );
ao12f80 g752169 ( .a(n_28038), .b(n_28037), .c(n_28036), .o(n_28143) );
in01f80 g774459 ( .a(n_6864), .o(n_6865) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_10_ ( .ck(newNet_1348), .d(n_1082), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_) );
na02f80 g755584 ( .a(n_45635), .b(n_22089), .o(n_24571) );
no02f80 g775667 ( .a(n_5340), .b(n_5440), .o(n_5442) );
na02f80 g738606 ( .a(n_41759), .b(n_41717), .o(n_41782) );
no02f80 g778606 ( .a(n_2266), .b(n_2359), .o(n_2267) );
in01f80 FE_OCP_RBC2148_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2144_FE_OCPN861_n_45450), .o(FE_OCP_RBN2148_FE_OCPN861_n_45450) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_5_ ( .ck(newNet_439), .d(n_27741), .o(delay_xor_ln22_unr18_stage7_stallmux_q_5_) );
oa12f80 g742631 ( .a(n_37316), .b(n_37399), .c(n_37426), .o(n_37449) );
na02f80 g770841 ( .a(n_9908), .b(n_9741), .o(n_9970) );
no02f80 g756268 ( .a(n_24080), .b(n_23775), .o(n_24094) );
na02f80 g759466 ( .a(n_20966), .b(n_20911), .o(n_20991) );
na02f80 g755242 ( .a(n_25018), .b(FE_OCP_RBN3843_n_24972), .o(n_25073) );
oa12f80 g754833 ( .a(n_25906), .b(n_25923), .c(n_25905), .o(n_26542) );
oa22f80 g748200 ( .a(FE_OCP_RBN3731_n_31819), .b(n_30573), .c(FE_OCPN880_n_31944), .d(n_30593), .o(n_32180) );
in01f80 g758526 ( .a(n_21951), .o(n_21968) );
no02f80 g758163 ( .a(n_44277), .b(n_21339), .o(n_22127) );
na02f80 g775949 ( .a(n_4807), .b(n_4717), .o(n_4808) );
na02f80 g770729 ( .a(n_10180), .b(n_10176), .o(n_10258) );
na02f80 g768360 ( .a(n_12523), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .o(n_12554) );
in01f80 g751818 ( .a(n_28928), .o(n_28929) );
in01f80 g758643 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_18_), .o(n_22455) );
na02f80 g742231 ( .a(n_44867), .b(n_37929), .o(n_37930) );
in01f80 FE_OCP_RBC3412_n_2100 ( .a(n_2100), .o(FE_OCP_RBN3412_n_2100) );
oa12f80 g745957 ( .a(n_33927), .b(n_33926), .c(n_33925), .o(n_35420) );
na02f80 g746724 ( .a(n_33234), .b(n_33189), .o(n_33270) );
in01f80 FE_OCP_RBC2413_n_13960 ( .a(FE_OCP_RBN3514_n_13960), .o(FE_OCP_RBN2413_n_13960) );
na02f80 g766162 ( .a(n_14443), .b(n_13515), .o(n_14513) );
no02f80 g763392 ( .a(FE_OCP_RBN1134_n_16041), .b(FE_OCP_RBN3725_n_16975), .o(n_17220) );
no02f80 g760488 ( .a(n_18676), .b(n_19922), .o(n_20005) );
oa12f80 g741227 ( .a(n_38941), .b(FE_OCPN942_n_44925), .c(n_38550), .o(n_39509) );
na02f80 g747147 ( .a(n_32700), .b(n_31650), .o(n_32775) );
in01f80 g755781 ( .a(n_26162), .o(n_26192) );
in01f80 FE_OCP_RBC2860_n_10399 ( .a(FE_OCP_RBN2859_n_10399), .o(FE_OCP_RBN2860_n_10399) );
in01f80 g760661 ( .a(n_19774), .o(n_19799) );
no02f80 g784779 ( .a(FE_OCP_RBN2902_n_44174), .b(n_34946), .o(n_47265) );
ao12f80 g780713 ( .a(n_623), .b(n_622), .c(n_621), .o(n_783) );
ao12f80 g763842 ( .a(n_16563), .b(n_16536), .c(n_16566), .o(n_16646) );
in01f80 newInst_950 ( .a(newNet_949), .o(newNet_950) );
in01f80 g770172 ( .a(n_10789), .o(n_10790) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_24_ ( .ck(newNet_3613), .d(n_17728), .o(delay_add_ln22_unr11_stage5_stallmux_q_24_) );
na02f80 g738224 ( .a(n_41924), .b(n_41850), .o(n_41971) );
in01f80 FE_OCP_RBC3223_n_22068 ( .a(FE_OCP_RBN3222_n_22068), .o(FE_OCP_RBN3223_n_22068) );
ao12f80 g777794 ( .a(n_2821), .b(n_3225), .c(n_2730), .o(n_3367) );
na02f80 g771242 ( .a(n_9356), .b(n_9397), .o(n_9502) );
no02f80 g742458 ( .a(n_37582), .b(n_36955), .o(n_37629) );
ao12f80 g751697 ( .a(n_29205), .b(n_29125), .c(n_28919), .o(n_29249) );
no02f80 g769029 ( .a(n_11728), .b(n_11727), .o(n_11852) );
no02f80 FE_RC_4073_0 ( .a(FE_RN_1773_0), .b(n_36416), .o(FE_RN_1775_0) );
oa22f80 g739622 ( .a(n_40586), .b(delay_sub_ln23_0_unr27_stage10_stallmux_z), .c(FE_OCP_RBN3108_n_40586), .d(n_40598), .o(n_40600) );
oa22f80 FE_RC_3781_0 ( .a(n_17344), .b(n_17312), .c(n_17404), .d(n_17311), .o(n_17591) );
oa12f80 g749653 ( .a(n_29984), .b(n_30154), .c(n_29916), .o(n_30226) );
in01f80 newInst_2652 ( .a(newNet_1814), .o(newNet_2652) );
in01f80 g767205 ( .a(FE_OCPN1006_n_13962), .o(n_14419) );
in01f80 g745047 ( .a(FE_OCP_RBN2642_n_34921), .o(n_35774) );
in01f80 g741631 ( .a(n_38624), .o(n_38637) );
na02f80 g737729 ( .a(n_42392), .b(n_42094), .o(n_42520) );
na02f80 g764971 ( .a(n_15389), .b(n_13950), .o(n_15390) );
oa12f80 g780227 ( .a(n_961), .b(n_960), .c(n_1155), .o(n_1065) );
na02f80 g758227 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .o(n_22654) );
in01f80 g756489 ( .a(n_23763), .o(n_23764) );
no02f80 g741856 ( .a(n_38360), .b(n_38359), .o(n_38361) );
in01f80 g783827 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .o(n_45512) );
in01f80 g760545 ( .a(n_19945), .o(n_19965) );
no02f80 g750297 ( .a(n_30756), .b(n_30811), .o(n_30893) );
in01f80 g775427 ( .a(n_5814), .o(n_5863) );
in01f80 g780625 ( .a(n_703), .o(n_704) );
in01f80 FE_OCP_RBC3431_n_33664 ( .a(n_33664), .o(FE_OCP_RBN3431_n_33664) );
in01f80 newInst_3012 ( .a(newNet_3011), .o(newNet_3012) );
in01f80 g765739 ( .a(n_15396), .o(n_15441) );
in01f80 g753659 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_2_), .o(n_26566) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_5_ ( .ck(newNet_3105), .d(n_40161), .o(delay_add_ln22_unr27_stage10_stallmux_q_5_) );
no02f80 g746985 ( .a(n_32857), .b(n_32319), .o(n_32936) );
no02f80 g773921 ( .a(n_6980), .b(n_6772), .o(n_7007) );
na02f80 g766170 ( .a(n_14591), .b(FE_OCP_RBN2509_n_13896), .o(n_14682) );
na02f80 g777902 ( .a(n_3119), .b(n_2329), .o(n_3164) );
na02f80 g758016 ( .a(n_22216), .b(n_22258), .o(n_22385) );
na02f80 g758995 ( .a(n_21425), .b(n_21497), .o(n_21538) );
na02f80 g765039 ( .a(n_15382), .b(n_15425), .o(n_15500) );
na02f80 g754863 ( .a(n_25923), .b(n_25905), .o(n_25906) );
in01f80 g754415 ( .a(n_25733), .o(n_25758) );
in01f80 g772827 ( .a(n_8073), .o(n_8089) );
no02f80 g770833 ( .a(n_9810), .b(n_8537), .o(n_9933) );
na02f80 g759987 ( .a(n_20375), .b(n_20374), .o(n_20441) );
no02f80 g741895 ( .a(n_38338), .b(n_38337), .o(n_38339) );
oa22f80 g743640 ( .a(n_36427), .b(n_35953), .c(n_36428), .d(n_35952), .o(n_36468) );
in01f80 newInst_3059 ( .a(newNet_1120), .o(newNet_3059) );
oa12f80 g746770 ( .a(n_32863), .b(n_32879), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n_32923) );
in01f80 g779805 ( .a(n_1601), .o(n_1630) );
in01f80 g769320 ( .a(n_11794), .o(n_11895) );
no02f80 g750057 ( .a(n_29869), .b(FE_OCP_RBN1324_n_29056), .o(n_29958) );
no02f80 g776697 ( .a(n_4256), .b(n_4072), .o(n_4345) );
na02f80 g777617 ( .a(n_3338), .b(n_3506), .o(n_3552) );
na02f80 g753768 ( .a(n_26478), .b(n_26473), .o(n_26497) );
no02f80 FE_RC_3059_0 ( .a(n_23564), .b(FE_RN_1341_0), .o(FE_RN_1342_0) );
na02f80 g752241 ( .a(FE_OCP_RBN2126_n_44734), .b(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .o(n_28005) );
in01f80 FE_OCP_RBC1368_n_20763 ( .a(n_20763), .o(FE_OCP_RBN1368_n_20763) );
oa22f80 g747970 ( .a(n_32184), .b(n_32182), .c(n_32185), .d(n_32183), .o(n_32252) );
in01f80 newInst_1098 ( .a(newNet_1097), .o(newNet_1098) );
no02f80 g770393 ( .a(n_10510), .b(n_10505), .o(n_10612) );
in01f80 g740272 ( .a(n_40212), .o(n_40213) );
in01f80 g772690 ( .a(n_8191), .o(n_8211) );
in01f80 g745324 ( .a(n_35886), .o(n_35887) );
in01f80 g750380 ( .a(n_29730), .o(n_29749) );
na02f80 g766678 ( .a(n_13729), .b(n_12900), .o(n_13730) );
ao12f80 g757955 ( .a(n_22787), .b(n_22786), .c(n_22785), .o(n_22882) );
no02f80 g752747 ( .a(n_27434), .b(n_27470), .o(n_27471) );
in01f80 FE_OCPC1779_n_24097 ( .a(n_24097), .o(FE_OCPN1779_n_24097) );
na02f80 g775176 ( .a(n_5802), .b(n_4875), .o(n_5870) );
no02f80 g771221 ( .a(n_9411), .b(FE_OCP_RBN3572_n_44563), .o(n_9462) );
no02f80 g772796 ( .a(n_8175), .b(n_8174), .o(n_8234) );
na02f80 g776891 ( .a(n_3607), .b(n_3642), .o(n_3867) );
no02f80 g740591 ( .a(n_39648), .b(n_39652), .o(n_39664) );
in01f80 newInst_3220 ( .a(newNet_3134), .o(newNet_3220) );
in01f80 g747369 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_9_), .o(n_32688) );
in01f80 g746606 ( .a(n_34609), .o(n_34610) );
in01f80 g756589 ( .a(n_23817), .o(n_23922) );
na02f80 g767436 ( .a(n_13395), .b(n_13394), .o(n_13396) );
in01f80 fopt782827 ( .a(n_44221), .o(n_44223) );
in01f80 newInst_2270 ( .a(newNet_2269), .o(newNet_2270) );
in01f80 newInst_3282 ( .a(newNet_2622), .o(newNet_3282) );
na02f80 g739224 ( .a(n_40675), .b(n_40493), .o(n_40701) );
oa12f80 g775880 ( .a(n_4844), .b(n_5234), .c(n_4808), .o(n_5359) );
na02f80 g764650 ( .a(n_15774), .b(n_15742), .o(n_15911) );
in01f80 FE_OCP_RBC2616_n_44561 ( .a(FE_OCP_RBN3573_n_44563), .o(FE_OCP_RBN2616_n_44561) );
oa22f80 FE_RC_1465_0 ( .a(n_17584), .b(n_17725), .c(n_17753), .d(n_17674), .o(n_17769) );
na02f80 g745594 ( .a(n_34286), .b(n_34350), .o(n_34401) );
no02f80 g773604 ( .a(n_7347), .b(n_7328), .o(n_7329) );
oa12f80 FE_RC_2178_0 ( .a(FE_RN_776_0), .b(n_26445), .c(FE_RN_777_0), .o(n_26627) );
na02f80 g752195 ( .a(n_28035), .b(n_28034), .o(n_28059) );
in01f80 newInst_219 ( .a(newNet_218), .o(newNet_219) );
na02f80 g764174 ( .a(n_16582), .b(FE_OCP_RBN1188_n_14823), .o(n_16637) );
ao12f80 g751852 ( .a(n_29100), .b(n_28919), .c(n_29068), .o(n_29757) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_22_ ( .ck(newNet_2095), .d(n_6419), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_) );
in01f80 FE_OCP_RBC3568_n_29857 ( .a(FE_OCP_RBN3565_n_29857), .o(FE_OCP_RBN3568_n_29857) );
na02f80 g779758 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .o(n_1663) );
in01f80 g778953 ( .a(n_2243), .o(n_2244) );
no02f80 g771847 ( .a(FE_OCP_RBN3546_n_44575), .b(FE_OCP_RBN3593_n_8902), .o(n_9049) );
in01f80 g768293 ( .a(n_12623), .o(n_12604) );
oa22f80 g784355 ( .a(FE_OFN86_n_46137), .b(n_6175), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_46995), .o(n_46161) );
na02f80 g755072 ( .a(n_25413), .b(n_25444), .o(n_25533) );
in01f80 g737603 ( .a(n_42262), .o(n_42263) );
in01f80 FE_OCP_RBC2542_n_38721 ( .a(n_38721), .o(FE_OCP_RBN2542_n_38721) );
in01f80 fopt783574 ( .a(n_45202), .o(n_45200) );
no02f80 g738548 ( .a(n_41582), .b(n_41321), .o(n_41735) );
na02f80 g741022 ( .a(n_39205), .b(n_39175), .o(n_39234) );
no02f80 g777783 ( .a(n_3391), .b(FE_OCP_RBN3489_n_3390), .o(n_3425) );
oa12f80 g741886 ( .a(n_38336), .b(n_38335), .c(n_38334), .o(n_38434) );
na02f80 FE_RC_2853_0 ( .a(n_13886), .b(n_14102), .o(FE_RN_1229_0) );
no03m80 FE_RC_3319_0 ( .a(n_14104), .b(n_14051), .c(n_14121), .o(n_14122) );
oa12f80 g752639 ( .a(n_28204), .b(n_28158), .c(n_27990), .o(n_28245) );
no02f80 g746140 ( .a(FE_OCP_RBN1355_n_44259), .b(n_33663), .o(n_33755) );
na02f80 g759121 ( .a(n_21461), .b(n_45080), .o(n_21489) );
in01f80 FE_OCP_RBC3424_n_37794 ( .a(n_37794), .o(FE_OCP_RBN3424_n_37794) );
in01f80 newInst_2405 ( .a(newNet_306), .o(newNet_2405) );
na02f80 g783830 ( .a(n_32090), .b(n_31880), .o(n_45516) );
no02f80 g766427 ( .a(n_14145), .b(n_13463), .o(n_14231) );
na02f80 g770820 ( .a(n_10215), .b(n_10214), .o(n_10251) );
in01f80 FE_OCP_RBC1329_n_18866 ( .a(n_18866), .o(FE_OCP_RBN1329_n_18866) );
no02f80 g771451 ( .a(n_9441), .b(n_7978), .o(n_9563) );
in01f80 g781219 ( .a(n_169), .o(n_164) );
ao12f80 g777412 ( .a(n_2937), .b(n_3456), .c(n_2877), .o(n_3526) );
in01f80 g740807 ( .a(n_39311), .o(n_39312) );
no02f80 g748258 ( .a(FE_OCP_RBN3083_n_31819), .b(n_31864), .o(n_31929) );
na02f80 g737012 ( .a(n_43230), .b(n_43418), .o(n_43497) );
oa12f80 g756438 ( .a(n_23678), .b(n_23884), .c(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n_23928) );
no02f80 FE_RC_3482_0 ( .a(n_37017), .b(n_37004), .o(FE_RN_1497_0) );
in01f80 g738260 ( .a(n_41952), .o(n_42271) );
oa12f80 g743773 ( .a(n_35694), .b(n_36324), .c(n_35872), .o(n_36206) );
no02f80 g738700 ( .a(n_41382), .b(n_41141), .o(n_41534) );
na02f80 g778911 ( .a(n_2324), .b(n_2300), .o(n_2333) );
no02f80 g766588 ( .a(n_13924), .b(n_13470), .o(n_13954) );
na02f80 g776428 ( .a(n_4585), .b(n_4198), .o(n_4641) );
ao12f80 g751276 ( .a(n_29205), .b(n_29721), .c(n_29150), .o(n_29771) );
in01f80 g768748 ( .a(n_12180), .o(n_12181) );
ao12f80 g748515 ( .a(n_31491), .b(n_31546), .c(n_31489), .o(n_31678) );
oa12f80 g736348 ( .a(n_43526), .b(n_43814), .c(n_43351), .o(n_43825) );
oa12f80 g767459 ( .a(n_13297), .b(n_13296), .c(n_13295), .o(n_14968) );
oa12f80 g774266 ( .a(n_6341), .b(n_6487), .c(n_6382), .o(n_6488) );
no02f80 g738765 ( .a(n_41358), .b(n_40864), .o(n_41374) );
oa12f80 g773041 ( .a(n_7802), .b(n_7849), .c(n_7848), .o(n_7850) );
na02f80 g757041 ( .a(n_23803), .b(n_23801), .o(n_23909) );
no02f80 g752146 ( .a(n_28617), .b(n_28616), .o(n_28618) );
na02f80 g774954 ( .a(n_6054), .b(n_6078), .o(n_6104) );
in01f80 newInst_2481 ( .a(newNet_912), .o(newNet_2481) );
in01f80 g777860 ( .a(n_3227), .o(n_3224) );
in01f80 FE_RC_2470_0 ( .a(n_14078), .o(FE_RN_995_0) );
na02f80 g740536 ( .a(FE_OCP_RBN2944_FE_RN_1269_0), .b(n_45514), .o(n_39683) );
no02f80 g784519 ( .a(n_11365), .b(n_10386), .o(n_46337) );
na02f80 g768740 ( .a(n_11993), .b(n_11998), .o(n_12039) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_30_ ( .ck(newNet_3288), .d(n_32338), .o(delay_add_ln22_unr20_stage8_stallmux_q_30_) );
in01f80 g744490 ( .a(n_35535), .o(n_35446) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_11_ ( .ck(newNet_3173), .d(n_40452), .o(delay_add_ln22_unr27_stage10_stallmux_q_11_) );
in01f80 newInst_876 ( .a(newNet_875), .o(newNet_876) );
no02f80 g744670 ( .a(n_35254), .b(n_35271), .o(n_35324) );
no02f80 FE_RC_3964_0 ( .a(FE_RN_1716_0), .b(n_24285), .o(n_24340) );
na02f80 g769966 ( .a(n_10894), .b(n_10884), .o(n_10895) );
na02f80 g767471 ( .a(n_13296), .b(n_13295), .o(n_13297) );
no02f80 g763369 ( .a(n_16912), .b(n_15351), .o(n_17045) );
no02f80 g768539 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .o(n_12368) );
in01f80 FE_OCP_RBC3082_n_16977 ( .a(FE_OCP_RBN3080_n_16977), .o(FE_OCP_RBN3082_n_16977) );
in01f80 FE_OCP_RBC1188_n_14823 ( .a(FE_OCP_RBN1187_n_14823), .o(FE_OCP_RBN1188_n_14823) );
no02f80 g749716 ( .a(n_31417), .b(n_31311), .o(n_31455) );
na02f80 g745521 ( .a(n_34348), .b(n_34347), .o(n_34349) );
no02f80 g772584 ( .a(n_8396), .b(n_8437), .o(n_8530) );
in01f80 FE_RC_4207_0 ( .a(FE_RN_1842_0), .o(n_19867) );
ao12f80 g739108 ( .a(n_41045), .b(n_41044), .c(n_41043), .o(n_41407) );
na02f80 g779529 ( .a(n_1580), .b(n_1441), .o(n_1581) );
in01f80 FE_RC_2484_0 ( .a(n_9591), .o(FE_RN_1003_0) );
in01f80 g747998 ( .a(n_31938), .o(n_31956) );
in01f80 newInst_3572 ( .a(newNet_2047), .o(newNet_3572) );
in01f80 g755426 ( .a(n_24891), .o(n_24910) );
na02f80 g778131 ( .a(n_3494), .b(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(n_2832) );
in01f80 FE_OCP_RBC2912_n_30908 ( .a(n_30908), .o(FE_OCP_RBN2912_n_30908) );
no02f80 g771409 ( .a(n_9634), .b(n_9604), .o(n_9834) );
na02f80 g767797 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_30_), .o(n_13193) );
na02f80 g751550 ( .a(n_28450), .b(n_28449), .o(n_28504) );
in01f80 g745303 ( .a(n_36169), .o(n_36170) );
na02f80 g767695 ( .a(n_13236), .b(n_13168), .o(n_13286) );
in01f80 newInst_2114 ( .a(newNet_2113), .o(newNet_2114) );
in01f80 newInst_3442 ( .a(newNet_3441), .o(newNet_3442) );
no02f80 g771945 ( .a(n_8696), .b(FE_OCP_RBN3467_n_7886), .o(n_8697) );
in01f80 FE_OCP_RBC2463_n_3076 ( .a(n_3076), .o(FE_OCP_RBN2463_n_3076) );
no02f80 FE_RC_2275_0 ( .a(FE_RN_847_0), .b(n_17605), .o(FE_RN_848_0) );
in01f80 newInst_472 ( .a(newNet_471), .o(newNet_472) );
in01f80 FE_OCP_RBC3853_n_20848 ( .a(FE_OCP_RBN3852_n_20848), .o(FE_OCP_RBN3853_n_20848) );
in01f80 g770276 ( .a(n_10801), .o(n_10836) );
na02f80 g745809 ( .a(n_44100), .b(n_34098), .o(n_34187) );
ao12f80 g779422 ( .a(n_2030), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_23_), .o(n_2353) );
na02f80 g765314 ( .a(n_15208), .b(n_15207), .o(n_15264) );
oa22f80 FE_RC_847_0 ( .a(n_23846), .b(n_24364), .c(n_23847), .d(n_24363), .o(n_24461) );
oa12f80 g778638 ( .a(FE_OCPN850_n_2306), .b(n_3082), .c(n_2255), .o(n_3207) );
na02f80 FE_RC_1673_0 ( .a(n_28308), .b(n_28309), .o(FE_RN_465_0) );
na02f80 g743381 ( .a(n_36613), .b(n_36750), .o(n_36659) );
ao12f80 g779504 ( .a(n_1913), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_19_), .o(n_2194) );
na02f80 g775265 ( .a(n_5731), .b(n_5772), .o(n_5881) );
na02f80 g772008 ( .a(FE_OCPN903_n_44581), .b(FE_OCPN1390_n_9220), .o(n_9281) );
ao12f80 g762813 ( .a(n_17727), .b(n_17656), .c(n_17726), .o(n_17826) );
no02f80 g750787 ( .a(n_29164), .b(n_28746), .o(n_29193) );
na02f80 g739071 ( .a(n_41065), .b(n_40796), .o(n_41092) );
in01f80 newInst_146 ( .a(newNet_145), .o(newNet_146) );
na02f80 g755702 ( .a(n_24447), .b(n_24446), .o(n_24448) );
na02f80 g776506 ( .a(n_4474), .b(n_4412), .o(n_4532) );
ao12f80 g763623 ( .a(n_17373), .b(n_17372), .c(n_17371), .o(n_18417) );
no02f80 FE_RC_1343_0 ( .a(FE_RN_401_0), .b(n_4453), .o(n_47008) );
in01f80 newInst_784 ( .a(newNet_783), .o(newNet_784) );
na02f80 g769258 ( .a(n_11480), .b(n_11479), .o(n_11481) );
na02f80 g749182 ( .a(n_30806), .b(n_30348), .o(n_30830) );
in01f80 fopt783146 ( .a(n_44659), .o(n_44661) );
oa12f80 g745698 ( .a(n_34843), .b(n_35433), .c(n_34805), .o(n_35479) );
in01f80 newInst_2610 ( .a(newNet_2609), .o(newNet_2610) );
in01f80 newInst_2902 ( .a(newNet_2901), .o(newNet_2902) );
ao22s80 g736400 ( .a(n_43731), .b(n_43546), .c(n_43732), .d(n_43545), .o(n_43774) );
in01f80 newInst_1316 ( .a(newNet_799), .o(newNet_1316) );
oa12f80 g760601 ( .a(n_19852), .b(n_20301), .c(n_19824), .o(n_20385) );
in01f80 newInst_2447 ( .a(newNet_2446), .o(newNet_2447) );
ao12f80 g779497 ( .a(n_2011), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .o(n_2046) );
in01f80 g742763 ( .a(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_43012) );
in01f80 g780396 ( .a(n_916), .o(n_938) );
na02f80 g762453 ( .a(FE_OCPN854_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .o(n_18050) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_3_ ( .ck(newNet_1185), .d(n_4192), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_) );
no02f80 g757502 ( .a(n_22932), .b(n_22864), .o(n_22989) );
in01f80 newInst_3140 ( .a(newNet_250), .o(newNet_3140) );
oa12f80 g776679 ( .a(n_4270), .b(n_4297), .c(n_4269), .o(n_4380) );
na02f80 g771896 ( .a(n_8804), .b(n_8799), .o(n_8968) );
na02f80 g757243 ( .a(n_23110), .b(n_23109), .o(n_23138) );
na02f80 g776197 ( .a(n_4963), .b(n_5017), .o(n_5228) );
in01f80 fopt783238 ( .a(n_44797), .o(n_44769) );
in01f80 FE_OCPC3756_n_13889 ( .a(n_13889), .o(FE_OCPN3756_n_13889) );
na02f80 g759720 ( .a(n_21798), .b(n_21691), .o(n_21831) );
no02f80 g778009 ( .a(n_3065), .b(n_3098), .o(n_3218) );
in01f80 g745719 ( .a(n_34307), .o(n_34308) );
in01f80 FE_OCP_RBC3664_n_35326 ( .a(n_35326), .o(FE_OCP_RBN3664_n_35326) );
in01f80 g739049 ( .a(n_41175), .o(n_41176) );
no02f80 g741574 ( .a(n_38615), .b(n_38778), .o(n_38632) );
in01f80 fopt783564 ( .a(n_40662), .o(n_45145) );
in01f80 newInst_2474 ( .a(newNet_2266), .o(newNet_2474) );
oa12f80 g780329 ( .a(n_690), .b(n_739), .c(n_706), .o(n_1104) );
in01f80 g750399 ( .a(n_29660), .o(n_29661) );
in01f80 g743281 ( .a(n_36771), .o(n_36772) );
na02f80 g770333 ( .a(n_10707), .b(FE_OCP_RBN2586_n_9009), .o(n_10811) );
no02f80 g751310 ( .a(n_28685), .b(n_28660), .o(n_28661) );
no02f80 g779378 ( .a(n_1524), .b(n_1548), .o(n_1623) );
no02f80 g773787 ( .a(n_7206), .b(n_6688), .o(n_7230) );
na02f80 g773202 ( .a(n_7599), .b(n_7726), .o(n_7626) );
no02f80 g763575 ( .a(n_16814), .b(n_16866), .o(n_16867) );
na02f80 g776290 ( .a(n_4697), .b(n_4695), .o(n_4696) );
in01f80 FE_RC_397_0 ( .a(n_15187), .o(FE_RN_117_0) );
in01f80 newInst_1265 ( .a(newNet_1264), .o(newNet_1265) );
oa12f80 g736299 ( .a(n_43644), .b(n_43846), .c(n_43562), .o(n_43880) );
ao22s80 FE_RC_4062_0 ( .a(n_26500), .b(n_26465), .c(n_26501), .d(n_26466), .o(n_26657) );
na02f80 g737440 ( .a(n_42722), .b(n_42721), .o(n_42723) );
in01f80 g759902 ( .a(n_21774), .o(n_21775) );
ao22s80 FE_RC_1360_0 ( .a(n_43604), .b(n_43799), .c(n_43603), .d(n_43798), .o(n_43845) );
in01f80 g773740 ( .a(n_7287), .o(n_7261) );
ao12f80 g739400 ( .a(n_40825), .b(FE_OCPN898_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(n_41134) );
na02f80 g778475 ( .a(n_2630), .b(n_2658), .o(n_2681) );
no02f80 g763908 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n_17360) );
in01f80 g746150 ( .a(n_33735), .o(n_34560) );
oa12f80 g772787 ( .a(n_7760), .b(n_8041), .c(n_7757), .o(n_8093) );
ao12f80 g748846 ( .a(n_30947), .b(n_31011), .c(n_31053), .o(n_31138) );
no02f80 g743189 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_3_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_3_), .o(n_36878) );
in01f80 FE_OCP_RBC2576_n_47017 ( .a(n_47017), .o(FE_OCP_RBN2576_n_47017) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_16_ ( .ck(newNet_2576), .d(n_27576), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_) );
oa12f80 g741755 ( .a(n_38328), .b(n_38455), .c(n_38378), .o(n_38481) );
no02f80 g750270 ( .a(n_30812), .b(n_30230), .o(n_30840) );
in01f80 newInst_825 ( .a(newNet_824), .o(newNet_825) );
in01f80 FE_OCP_RBC2853_n_26169 ( .a(n_26169), .o(FE_OCP_RBN2853_n_26169) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_7_ ( .ck(newNet_1465), .d(n_31779), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_) );
in01f80 newInst_3083 ( .a(newNet_165), .o(newNet_3083) );
na02f80 g772950 ( .a(n_7846), .b(n_7825), .o(n_7992) );
in01f80 FE_OCP_RBC2314_n_41420 ( .a(n_41420), .o(FE_OCP_RBN2314_n_41420) );
in01f80 newInst_963 ( .a(newNet_391), .o(newNet_963) );
in01f80 g778583 ( .a(n_2530), .o(n_2608) );
in01f80 newInst_1526 ( .a(newNet_1525), .o(newNet_1526) );
oa12f80 g764813 ( .a(n_16357), .b(n_16356), .c(n_16355), .o(n_16413) );
in01f80 FE_OCP_RBC3062_FE_RN_640_0 ( .a(FE_RN_640_0), .o(FE_OCP_RBN3062_FE_RN_640_0) );
ao12f80 g745769 ( .a(n_34414), .b(n_44102), .c(n_33500), .o(n_34596) );
in01f80 g749778 ( .a(n_31317), .o(n_31318) );
na02f80 g741058 ( .a(FE_OCP_RBN3623_n_39097), .b(n_39098), .o(n_39189) );
in01f80 g775809 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .o(n_5393) );
in01f80 g765238 ( .a(n_15059), .o(n_15060) );
oa22f80 g779222 ( .a(n_1820), .b(n_1483), .c(n_1821), .d(n_1482), .o(n_2364) );
no02f80 g736588 ( .a(n_43417), .b(n_43114), .o(n_43528) );
no02f80 g751959 ( .a(n_28919), .b(n_28899), .o(n_29071) );
ao22s80 FE_RC_1706_0 ( .a(n_21438), .b(n_21512), .c(n_21511), .d(n_21439), .o(n_21656) );
no02f80 g742135 ( .a(n_38292), .b(n_38303), .o(n_38412) );
oa22f80 FE_RC_3217_0 ( .a(n_11748), .b(n_11953), .c(FE_RN_1428_0), .d(n_11952), .o(n_12145) );
no02f80 g768837 ( .a(n_11978), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .o(n_12091) );
in01f80 FE_OFC751_n_45003 ( .a(FE_OFN749_n_45003), .o(FE_OFN751_n_45003) );
no02f80 g737459 ( .a(n_42638), .b(n_42653), .o(n_43132) );
na02f80 g743030 ( .a(n_37051), .b(n_37101), .o(n_37155) );
oa22f80 FE_RC_1141_0 ( .a(n_36763), .b(n_36894), .c(n_36764), .d(n_36867), .o(n_36895) );
no02f80 g737743 ( .a(FE_OCPN885_n_42216), .b(n_42067), .o(n_42468) );
na02f80 g768918 ( .a(n_11760), .b(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n_12124) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_25_ ( .ck(newNet_807), .d(n_1346), .o(delay_xor_ln21_unr3_stage2_stallmux_q_25_) );
na02f80 FE_RC_3162_0 ( .a(FE_RN_1401_0), .b(n_27204), .o(n_27400) );
ao12f80 g770658 ( .a(n_9891), .b(FE_OCP_RBN3636_n_47260), .c(FE_OCP_RBN2823_n_10068), .o(n_10203) );
in01f80 g754187 ( .a(n_26045), .o(n_26044) );
in01f80 newInst_2127 ( .a(newNet_2126), .o(newNet_2127) );
no02f80 g780456 ( .a(FE_OFN794_n_45813), .b(n_1099), .o(n_840) );
in01f80 g758337 ( .a(n_22326), .o(n_22327) );
in01f80 FE_OCP_RBC3820_n_44061 ( .a(FE_OCP_RBN3821_n_44061), .o(FE_OCP_RBN3820_n_44061) );
no02f80 g746011 ( .a(n_35259), .b(n_35258), .o(n_35260) );
na02f80 g753824 ( .a(n_26322), .b(n_23467), .o(n_26372) );
ao12f80 g738117 ( .a(n_41722), .b(n_42031), .c(n_41657), .o(n_42062) );
ao12f80 g767328 ( .a(n_13493), .b(n_13492), .c(n_13491), .o(n_15223) );
na02f80 g764414 ( .a(n_16202), .b(n_16157), .o(n_16203) );
na02f80 g737677 ( .a(n_42392), .b(n_42049), .o(n_42801) );
na02f80 g772905 ( .a(n_7882), .b(n_7852), .o(n_8017) );
in01f80 g766880 ( .a(n_14421), .o(n_14488) );
in01f80 g740045 ( .a(n_40330), .o(n_40331) );
no02f80 g765827 ( .a(n_14873), .b(FE_OCP_RBN2506_n_13896), .o(n_14958) );
no02f80 g765773 ( .a(n_14957), .b(n_14941), .o(n_15077) );
no02f80 g770414 ( .a(n_10477), .b(n_44463), .o(n_10505) );
in01f80 FE_OFC828_n_29140 ( .a(n_29140), .o(FE_OFN828_n_29140) );
in01f80 g749376 ( .a(n_30670), .o(n_30698) );
no03m80 g742874 ( .a(n_37002), .b(n_37077), .c(n_37072), .o(n_37186) );
no02f80 g743093 ( .a(n_36950), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_36988) );
in01f80 g763263 ( .a(n_17195), .o(n_17235) );
na02f80 g737769 ( .a(n_42546), .b(n_42582), .o(n_42629) );
in01f80 newInst_3418 ( .a(newNet_3417), .o(newNet_3418) );
in01f80 g744221 ( .a(n_36289), .o(n_36290) );
in01f80 g745827 ( .a(n_34196), .o(n_34687) );
ao12f80 g762673 ( .a(n_18236), .b(n_18235), .c(n_18234), .o(n_18441) );
oa22f80 g762603 ( .a(n_18253), .b(n_17707), .c(n_18254), .d(n_17706), .o(n_18492) );
in01f80 g756147 ( .a(n_24165), .o(n_24179) );
in01f80 g742013 ( .a(n_38374), .o(n_38375) );
na02f80 g772798 ( .a(n_8125), .b(n_8124), .o(n_8126) );
in01f80 newInst_3482 ( .a(newNet_3481), .o(newNet_3482) );
in01f80 g772308 ( .a(n_8653), .o(n_8654) );
in01f80 g766655 ( .a(n_14015), .o(n_14016) );
in01f80 newInst_2040 ( .a(newNet_2039), .o(newNet_2040) );
in01f80 g754561 ( .a(n_26683), .o(n_26684) );
no02f80 g744602 ( .a(FE_OCP_RBN1373_n_35275), .b(n_35294), .o(n_35296) );
ao22s80 FE_RC_3734_0 ( .a(FE_RN_1550_0), .b(FE_RN_1551_0), .c(n_24462), .d(FE_RN_1552_0), .o(n_24614) );
in01f80 g778183 ( .a(n_2865), .o(n_2785) );
in01f80 g743637 ( .a(n_36398), .o(n_36399) );
na02f80 g772961 ( .a(n_7748), .b(n_7027), .o(n_7847) );
no02f80 FE_RC_2815_0 ( .a(n_34364), .b(FE_RN_1205_0), .o(n_34908) );
in01f80 g739617 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .o(n_40624) );
no02f80 g746488 ( .a(n_34700), .b(n_34641), .o(n_34701) );
no02f80 g763674 ( .a(n_17372), .b(n_17371), .o(n_17373) );
no02f80 g753582 ( .a(n_26622), .b(n_23590), .o(n_26673) );
na02f80 g740458 ( .a(n_39701), .b(n_39710), .o(n_39741) );
no02f80 g775870 ( .a(n_5240), .b(n_5194), .o(n_5195) );
na02f80 g765296 ( .a(n_15925), .b(n_15924), .o(n_15964) );
in01f80 newInst_920 ( .a(newNet_687), .o(newNet_920) );
oa12f80 g780699 ( .a(n_639), .b(n_638), .c(n_637), .o(n_839) );
in01f80 g760384 ( .a(n_21591), .o(n_20809) );
no02f80 g748342 ( .a(n_31733), .b(n_31764), .o(n_31833) );
in01f80 FE_OCP_RBC3726_FE_RN_1787_0 ( .a(FE_RN_1787_0), .o(FE_OCP_RBN3726_FE_RN_1787_0) );
ao22s80 FE_RC_254_0 ( .a(n_13154), .b(FE_OCP_RBN2230_n_13141), .c(FE_OCP_RBN2233_n_13141), .d(n_13185), .o(n_13331) );
in01f80 g770531 ( .a(FE_OCP_RBN2860_n_10399), .o(n_10451) );
na02f80 g760970 ( .a(n_19375), .b(n_19344), .o(n_19499) );
oa12f80 g743322 ( .a(n_37841), .b(n_37840), .c(n_37839), .o(n_38021) );
na02f80 g779175 ( .a(n_1874), .b(n_1744), .o(n_1868) );
in01f80 g757446 ( .a(n_23094), .o(n_23390) );
na02f80 g749905 ( .a(n_30196), .b(n_30138), .o(n_30202) );
in01f80 FE_OCP_RBC2913_n_30949 ( .a(n_30949), .o(FE_OCP_RBN2913_n_30949) );
no02f80 FE_RC_3089_0 ( .a(FE_RN_1363_0), .b(n_31443), .o(n_31492) );
na02f80 g762040 ( .a(n_18847), .b(n_18845), .o(n_18846) );
no02f80 g758771 ( .a(n_22210), .b(n_21669), .o(n_22246) );
in01f80 newInst_2262 ( .a(newNet_634), .o(newNet_2262) );
na02f80 g772471 ( .a(n_8416), .b(n_8404), .o(n_10214) );
oa12f80 g752772 ( .a(n_27899), .b(n_27902), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n_27928) );
no02f80 g765539 ( .a(FE_OCP_RBN1170_n_13756), .b(FE_OCP_RBN2714_n_14982), .o(n_15391) );
in01f80 g743996 ( .a(n_36032), .o(n_36033) );
in01f80 g769948 ( .a(n_11074), .o(n_11102) );
na02f80 g771666 ( .a(n_9482), .b(n_9429), .o(n_9430) );
in01f80 g771175 ( .a(n_9514), .o(n_9515) );
in01f80 g771546 ( .a(n_9083), .o(n_9084) );
in01f80 g770537 ( .a(n_10554), .o(n_10555) );
na02f80 g742226 ( .a(n_44887), .b(n_38270), .o(n_38347) );
in01f80 newInst_1982 ( .a(newNet_1981), .o(newNet_1982) );
in01f80 newInst_1224 ( .a(newNet_1223), .o(newNet_1224) );
na02f80 g756272 ( .a(n_24606), .b(n_24091), .o(n_24670) );
in01f80 g739134 ( .a(n_40979), .o(n_40993) );
na02f80 g745636 ( .a(n_35461), .b(n_35159), .o(n_35496) );
in01f80 FE_OCP_RBC3817_n_44061 ( .a(n_44061), .o(FE_OCP_RBN3817_n_44061) );
oa22f80 FE_RC_722_0 ( .a(n_22961), .b(n_22778), .c(n_22580), .d(n_22757), .o(n_22832) );
in01f80 newInst_1834 ( .a(newNet_1587), .o(newNet_1834) );
na02f80 g778349 ( .a(n_2495), .b(n_2494), .o(n_2535) );
no02f80 g773171 ( .a(n_7802), .b(n_7801), .o(n_7839) );
na02f80 g755817 ( .a(n_24342), .b(n_24341), .o(n_24343) );
in01f80 g748177 ( .a(n_32128), .o(n_32129) );
in01f80 newInst_664 ( .a(newNet_44), .o(newNet_664) );
no02f80 g743170 ( .a(n_36910), .b(n_36909), .o(n_36911) );
no02f80 g755059 ( .a(n_25554), .b(n_25553), .o(n_25555) );
na02f80 g736498 ( .a(n_43701), .b(n_43367), .o(n_43716) );
in01f80 FE_OCP_RBC3107_n_22590 ( .a(n_22590), .o(FE_OCP_RBN3107_n_22590) );
no02f80 g776517 ( .a(n_4309), .b(n_4341), .o(n_4529) );
oa12f80 g775790 ( .a(n_5295), .b(n_5339), .c(n_5294), .o(n_5399) );
na02f80 g761903 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .o(n_18741) );
na02f80 g766755 ( .a(n_14085), .b(n_14083), .o(n_14084) );
no02f80 g780725 ( .a(n_612), .b(n_611), .o(n_613) );
na02f80 g766414 ( .a(n_14093), .b(n_13133), .o(n_14132) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_14_ ( .ck(newNet_2876), .d(n_11177), .o(delay_add_ln22_unr8_stage4_stallmux_q_14_) );
no02f80 g747414 ( .a(FE_OCP_RBN2102_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .o(n_32704) );
na02f80 g777722 ( .a(n_3324), .b(n_2567), .o(n_3358) );
in01f80 g765495 ( .a(n_15781), .o(n_15925) );
in01f80 g758856 ( .a(n_21838), .o(n_21839) );
na02f80 FE_RC_4152_0 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_5_), .b(n_23137), .o(FE_RN_1806_0) );
in01f80 g776264 ( .a(n_4505), .o(n_4506) );
ao12f80 g751380 ( .a(n_28513), .b(n_28535), .c(n_28512), .o(n_29777) );
in01f80 FE_OCP_RBC2425_n_47023 ( .a(n_47023), .o(FE_OCP_RBN2425_n_47023) );
oa22f80 FE_RC_1473_0 ( .a(FE_OFN767_n_15670), .b(n_17591), .c(n_17753), .d(FE_OCP_RBN3130_n_17591), .o(n_17647) );
na02f80 g780867 ( .a(n_354), .b(beta_2), .o(n_363) );
no02f80 g772743 ( .a(n_8093), .b(n_7767), .o(n_8131) );
oa12f80 g761387 ( .a(n_19579), .b(n_19578), .c(n_19577), .o(n_20036) );
no02f80 g764507 ( .a(n_16216), .b(n_16215), .o(n_16266) );
na03f80 FE_RC_3226_0 ( .a(n_8439), .b(n_8506), .c(n_8528), .o(n_8579) );
in01f80 newInst_1503 ( .a(newNet_1502), .o(newNet_1503) );
in01f80 newInst_1157 ( .a(newNet_1156), .o(newNet_1157) );
ao12f80 g751712 ( .a(n_28359), .b(n_28360), .c(n_27976), .o(n_28361) );
no02f80 g762290 ( .a(n_18607), .b(n_18694), .o(n_19367) );
ao12f80 g751920 ( .a(n_29000), .b(n_28919), .c(n_28982), .o(n_29637) );
ao12f80 g751335 ( .a(n_29461), .b(n_29460), .c(n_29459), .o(n_29999) );
oa12f80 g738318 ( .a(n_41541), .b(n_41818), .c(n_41683), .o(n_41737) );
in01f80 g778351 ( .a(n_2633), .o(n_2676) );
no02f80 FE_RC_2846_0 ( .a(n_38698), .b(n_38766), .o(FE_RN_1225_0) );
ao12f80 g749556 ( .a(n_30490), .b(n_30489), .c(n_30488), .o(n_31502) );
in01f80 g736616 ( .a(n_43334), .o(n_43376) );
oa12f80 g742614 ( .a(n_37466), .b(n_37465), .c(n_37464), .o(n_38269) );
no02f80 g759132 ( .a(n_21160), .b(n_21187), .o(n_21354) );
na02f80 g749931 ( .a(n_30372), .b(n_30371), .o(n_30373) );
na02f80 g777883 ( .a(n_3275), .b(n_3274), .o(n_3356) );
no02f80 g777263 ( .a(n_3577), .b(n_3645), .o(n_3646) );
in01f80 g749948 ( .a(n_30143), .o(n_30144) );
in01f80 g751295 ( .a(n_29709), .o(n_29710) );
in01f80 FE_OCPC1454_n_18559 ( .a(FE_OCPN1453_n_18559), .o(FE_OCPN1454_n_18559) );
ao12f80 g780782 ( .a(n_520), .b(n_519), .c(n_518), .o(n_545) );
in01f80 g750664 ( .a(n_29343), .o(n_29344) );
no02f80 g756065 ( .a(n_24247), .b(n_24263), .o(n_24362) );
no02f80 g769046 ( .a(FE_OCP_RBN3271_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .o(n_11844) );
in01f80 FE_OCP_RBC2380_n_3502 ( .a(n_3502), .o(FE_OCP_RBN2380_n_3502) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_5_ ( .ck(newNet_1927), .d(n_36866), .o(delay_sub_ln21_unr24_stage9_stallmux_q_5_) );
in01f80 FE_OCP_RBC2279_n_24199 ( .a(n_24199), .o(FE_OCP_RBN2279_n_24199) );
ao12f80 g768350 ( .a(n_12472), .b(n_12471), .c(n_12470), .o(n_12840) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_14_ ( .ck(newNet_3644), .d(n_16686), .o(delay_add_ln22_unr11_stage5_stallmux_q_14_) );
in01f80 g756211 ( .a(n_24161), .o(n_24176) );
in01f80 g745288 ( .a(n_35966), .o(n_35967) );
in01f80 g751829 ( .a(n_28271), .o(n_28251) );
no02f80 g753942 ( .a(n_26152), .b(FE_OCPN1508_n_23414), .o(n_26191) );
na02f80 g742259 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37415), .o(n_38208) );
in01f80 g755802 ( .a(n_24367), .o(n_24368) );
na02f80 g766764 ( .a(n_13722), .b(n_13721), .o(n_13753) );
na02f80 g752043 ( .a(n_28164), .b(n_28163), .o(n_28165) );
na02f80 g738014 ( .a(n_42173), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42174) );
ao12f80 g778751 ( .a(n_2355), .b(n_2354), .c(n_2353), .o(n_2420) );
no02f80 g752396 ( .a(n_28399), .b(FE_RN_520_0), .o(n_28457) );
ao12f80 g765808 ( .a(n_14697), .b(n_14775), .c(n_14754), .o(n_14830) );
no02f80 g756451 ( .a(n_23736), .b(n_23735), .o(n_23771) );
no02f80 g747738 ( .a(n_33414), .b(n_33462), .o(n_33463) );
no02f80 g777151 ( .a(n_4901), .b(n_4834), .o(n_4885) );
oa22f80 g743296 ( .a(n_36708), .b(delay_add_ln22_unr23_stage9_stallmux_q_0_), .c(n_35362), .d(delay_sub_ln22_unr24_stage9_stallmux_q_0_), .o(n_37504) );
in01f80 newInst_3017 ( .a(newNet_3016), .o(newNet_3017) );
ao12f80 g740996 ( .a(n_38831), .b(n_38968), .c(n_38894), .o(n_38934) );
na02f80 g769719 ( .a(n_11199), .b(n_11218), .o(n_11244) );
na02f80 g742468 ( .a(n_37606), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37628) );
in01f80 FE_RC_177_0 ( .a(beta_1), .o(FE_RN_56_0) );
in01f80 g750889 ( .a(n_29157), .o(n_29135) );
in01f80 FE_RC_1184_0 ( .a(n_13017), .o(FE_RN_357_0) );
oa12f80 g742422 ( .a(n_37709), .b(n_37703), .c(n_37667), .o(n_37753) );
oa22f80 g753701 ( .a(n_27108), .b(n_26683), .c(n_27109), .d(n_26684), .o(n_27200) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_16_ ( .ck(newNet_2208), .d(n_1022), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_) );
in01f80 g745557 ( .a(n_34702), .o(n_34703) );
in01f80 g761251 ( .a(n_19075), .o(n_19076) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_9_ ( .ck(newNet_1161), .d(n_5151), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_) );
in01f80 newInst_917 ( .a(newNet_916), .o(newNet_917) );
in01f80 FE_RC_4185_0 ( .a(FE_RN_1831_0), .o(FE_RN_1830_0) );
oa22f80 g784363 ( .a(FE_OFN805_n_46196), .b(n_5363), .c(FE_OFN775_n_46137), .d(n_5324), .o(n_46169) );
na02f80 g767408 ( .a(n_13334), .b(n_12914), .o(n_13405) );
in01f80 g766213 ( .a(n_14380), .o(n_14417) );
in01f80 g765875 ( .a(n_14881), .o(n_14882) );
in01f80 newInst_2148 ( .a(newNet_586), .o(newNet_2148) );
in01f80 g736895 ( .a(n_43585), .o(n_43586) );
in01f80 g745583 ( .a(n_34316), .o(n_34317) );
no02f80 g753255 ( .a(n_27110), .b(n_25873), .o(n_27141) );
na02f80 g748584 ( .a(n_31383), .b(n_31244), .o(n_31384) );
no02f80 g739124 ( .a(n_41044), .b(n_41043), .o(n_41045) );
na02f80 g749751 ( .a(n_31120), .b(n_31119), .o(n_31121) );
in01f80 FE_OCP_RBC2730_n_4219 ( .a(FE_OCP_RBN2726_n_4219), .o(FE_OCP_RBN2730_n_4219) );
na02f80 g759487 ( .a(n_20619), .b(n_20596), .o(n_20734) );
na02f80 g767053 ( .a(n_14215), .b(n_14207), .o(n_14561) );
na02f80 g776022 ( .a(FE_OCP_RBN2819_n_4872), .b(n_4879), .o(n_4937) );
in01f80 FE_OCPC996_n_44460 ( .a(FE_OCP_RBN3573_n_44563), .o(FE_OCPN996_n_44460) );
in01f80 FE_OCP_RBC3434_n_2224 ( .a(n_2224), .o(FE_OCP_RBN3434_n_2224) );
no02f80 g754025 ( .a(n_26139), .b(n_23414), .o(n_26205) );
ao22s80 FE_RC_59_0 ( .a(n_18219), .b(n_18289), .c(n_18218), .d(n_18290), .o(n_18375) );
in01f80 newInst_1752 ( .a(newNet_1249), .o(newNet_1752) );
in01f80 FE_OCP_RBC2302_n_7817 ( .a(FE_OCP_RBN2300_n_7817), .o(FE_OCP_RBN2302_n_7817) );
no02f80 g763054 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_17555) );
no02f80 g748153 ( .a(n_31772), .b(n_31871), .o(n_31850) );
in01f80 g736457 ( .a(n_43744), .o(n_43745) );
in01f80 g742300 ( .a(FE_OCP_RBN2256_n_37844), .o(n_37900) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_6_ ( .ck(newNet_293), .d(n_1360), .o(delay_xor_ln22_unr3_stage2_stallmux_q_6_) );
na02f80 g766133 ( .a(n_14556), .b(n_14555), .o(n_14636) );
in01f80 newInst_9 ( .a(newNet_8), .o(newNet_9) );
in01f80 FE_OFC806_n_46196 ( .a(FE_OFN804_n_46196), .o(FE_OFN806_n_46196) );
na02f80 g740456 ( .a(n_39774), .b(n_39759), .o(n_39788) );
no02f80 g742046 ( .a(FE_OCP_RBN3444_n_37945), .b(FE_OCP_RBN2174_n_37559), .o(n_38088) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_30_ ( .ck(newNet_1482), .d(n_32378), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_) );
no03m80 FE_RC_3055_0 ( .a(n_16171), .b(n_16166), .c(n_16236), .o(n_16237) );
oa12f80 g773719 ( .a(n_6938), .b(n_7270), .c(n_6878), .o(n_7303) );
oa12f80 g761681 ( .a(n_18749), .b(n_18795), .c(n_18748), .o(n_18895) );
in01f80 g739433 ( .a(n_40723), .o(n_40841) );
in01f80 newInst_417 ( .a(newNet_416), .o(newNet_417) );
no02f80 g743517 ( .a(n_36545), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36561) );
no02f80 g749827 ( .a(FE_OCP_RBN3013_n_31117), .b(n_31172), .o(n_31509) );
in01f80 FE_OCP_RBC2899_n_44853 ( .a(n_44853), .o(FE_OCP_RBN2899_n_44853) );
na02f80 g748404 ( .a(FE_OCP_RBN3712_n_31466), .b(FE_OCP_RBN1198_n_30619), .o(n_31553) );
na02f80 g766827 ( .a(n_14422), .b(n_14306), .o(n_15361) );
in01f80 FE_OCPC3164_n_24117 ( .a(FE_OCPN3163_n_24117), .o(FE_OCPN3164_n_24117) );
in01f80 newInst_1261 ( .a(newNet_227), .o(newNet_1261) );
ao12f80 g742852 ( .a(n_37089), .b(n_37193), .c(n_37209), .o(n_37251) );
na02f80 g743319 ( .a(n_36786), .b(n_36765), .o(n_36796) );
oa12f80 g782639 ( .a(n_44877), .b(n_37965), .c(n_38290), .o(n_44032) );
na02f80 g774086 ( .a(n_6832), .b(delay_add_ln22_unr5_stage3_stallmux_q_2_), .o(n_6847) );
in01f80 g761168 ( .a(n_21105), .o(n_21134) );
na02f80 FE_RC_3983_0 ( .a(FE_RN_1726_0), .b(n_13980), .o(n_14115) );
na02f80 g769566 ( .a(n_11392), .b(n_11479), .o(n_11398) );
no02f80 g765930 ( .a(n_14798), .b(FE_OCP_RBN3528_n_13765), .o(n_14800) );
in01f80 g745612 ( .a(n_34509), .o(n_34857) );
in01f80 FE_OCP_RBC2319_n_2367 ( .a(FE_OCP_RBN2318_n_2367), .o(FE_OCP_RBN2319_n_2367) );
oa12f80 g753857 ( .a(n_26295), .b(n_26294), .c(n_26293), .o(n_26365) );
no02f80 g756001 ( .a(n_24994), .b(n_25001), .o(n_25056) );
no02f80 g771679 ( .a(n_9028), .b(n_44516), .o(n_10341) );
na02f80 g757260 ( .a(n_23069), .b(delay_add_ln22_unr14_stage6_stallmux_q_4_), .o(n_23197) );
no02f80 g772672 ( .a(n_8315), .b(n_8343), .o(n_8445) );
no02f80 g775210 ( .a(n_5945), .b(n_5148), .o(n_6062) );
na02f80 g773894 ( .a(n_7020), .b(n_5430), .o(n_7085) );
in01f80 g749225 ( .a(n_32201), .o(n_32202) );
no02f80 g771870 ( .a(n_44575), .b(n_8902), .o(n_8988) );
in01f80 g773802 ( .a(n_7715), .o(n_7215) );
in01f80 g749469 ( .a(FE_OCP_RBN2804_n_30534), .o(n_30557) );
in01f80 newInst_1422 ( .a(newNet_1421), .o(newNet_1422) );
no02f80 g741931 ( .a(n_38092), .b(n_38069), .o(n_38070) );
in01f80 g766202 ( .a(n_14539), .o(n_14540) );
oa22f80 FE_RC_1653_0 ( .a(n_16530), .b(n_16390), .c(n_16391), .d(n_16531), .o(n_16622) );
na02f80 g739159 ( .a(n_40896), .b(n_40792), .o(n_40913) );
no02f80 g780926 ( .a(n_457), .b(n_495), .o(n_498) );
oa12f80 g771027 ( .a(n_9925), .b(n_9924), .c(n_9923), .o(n_10000) );
ao12f80 g745781 ( .a(n_34813), .b(n_35408), .c(n_34804), .o(n_35433) );
in01f80 FE_OCP_DRV_C1544_n_18854 ( .a(FE_OCP_DRV_N1543_n_18854), .o(FE_OCP_DRV_N1544_n_18854) );
ao12f80 g780940 ( .a(n_56), .b(n_284), .c(n_128), .o(n_285) );
na02f80 g748037 ( .a(n_31708), .b(n_31751), .o(n_31813) );
in01f80 g776806 ( .a(n_4275), .o(n_4276) );
in01f80 g781270 ( .a(n_113), .o(n_114) );
ao12f80 g772839 ( .a(n_7936), .b(n_8066), .c(n_7984), .o(n_8057) );
na02f80 g776108 ( .a(n_5015), .b(n_3697), .o(n_5145) );
no02f80 g755032 ( .a(n_25103), .b(n_23888), .o(n_25182) );
no02f80 g757258 ( .a(n_23136), .b(n_23135), .o(n_23169) );
in01f80 FE_OCPC1517_n_26752 ( .a(n_26752), .o(FE_OCPN1517_n_26752) );
no02f80 g767944 ( .a(n_12885), .b(n_12911), .o(n_12920) );
ao12f80 g762752 ( .a(n_17825), .b(FE_OCP_RBN2140_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .o(n_17847) );
in01f80 g761490 ( .a(n_19822), .o(n_19823) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_15_ ( .ck(newNet_3549), .d(n_22392), .o(delay_add_ln22_unr14_stage6_stallmux_q_15_) );
na02f80 g759512 ( .a(FE_OCP_RBN1366_n_20879), .b(n_20912), .o(n_20963) );
ao12f80 g778492 ( .a(n_2061), .b(n_2369), .c(n_2032), .o(n_2428) );
in01f80 FE_RC_2692_0 ( .a(FE_RN_1128_0), .o(n_4134) );
no02f80 g742991 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n_37003) );
na02f80 FE_RC_3584_0 ( .a(FE_RN_1558_0), .b(FE_RN_1562_0), .o(n_14672) );
no02f80 g769352 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_13_), .o(n_11796) );
na02f80 g767652 ( .a(n_13284), .b(n_13242), .o(n_13379) );
in01f80 g738761 ( .a(n_41364), .o(n_41365) );
in01f80 FE_OCP_RBC3115_n_6379 ( .a(n_6379), .o(FE_OCP_RBN3115_n_6379) );
in01f80 fopt782960 ( .a(n_44422), .o(n_44420) );
na02f80 g744701 ( .a(n_35199), .b(n_34056), .o(n_35266) );
no02f80 g746537 ( .a(n_35069), .b(n_34586), .o(n_35160) );
no02f80 g752133 ( .a(n_46961), .b(delay_add_ln22_unr17_stage7_stallmux_q_3_), .o(n_28093) );
na02f80 g749318 ( .a(n_32008), .b(n_31390), .o(n_32094) );
ao22s80 FE_RC_1799_0 ( .a(FE_RN_531_0), .b(FE_RN_530_0), .c(n_33984), .d(n_46955), .o(n_34066) );
in01f80 g773389 ( .a(n_7660), .o(n_7661) );
in01f80 g744315 ( .a(n_35519), .o(n_35520) );
no02f80 g744234 ( .a(n_36811), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n_36860) );
ao22s80 FE_RC_3873_0 ( .a(n_33267), .b(n_33687), .c(n_33268), .d(n_33688), .o(n_33771) );
in01f80 g772900 ( .a(n_7967), .o(n_7968) );
in01f80 g764024 ( .a(n_18099), .o(n_18117) );
no02f80 g751734 ( .a(n_28347), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .o(n_28355) );
in01f80 g737466 ( .a(n_42669), .o(n_42670) );
in01f80 g771181 ( .a(n_9510), .o(n_9511) );
in01f80 g742662 ( .a(n_37554), .o(n_37569) );
no02f80 g753875 ( .a(n_26221), .b(n_26251), .o(n_26299) );
ao12f80 g777665 ( .a(n_2541), .b(n_3313), .c(n_2582), .o(n_3386) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_2_ ( .ck(newNet_889), .d(n_32352), .o(delay_xor_ln21_unr21_stage8_stallmux_q_2_) );
no02f80 g736731 ( .a(n_43255), .b(n_43280), .o(n_43433) );
in01f80 g768416 ( .a(n_12414), .o(n_12415) );
na02f80 g739667 ( .a(n_40532), .b(n_40221), .o(n_40546) );
ao12f80 g761369 ( .a(n_19787), .b(n_19927), .c(n_19873), .o(n_19988) );
no02f80 g747542 ( .a(n_33397), .b(n_33759), .o(n_33814) );
in01f80 FE_RC_2432_0 ( .a(n_6940), .o(FE_RN_968_0) );
in01f80 FE_OCP_RBC3621_n_15135 ( .a(FE_OCP_RBN3620_n_15135), .o(FE_OCP_RBN3621_n_15135) );
ao12f80 g755760 ( .a(n_25160), .b(n_25259), .c(n_25258), .o(n_25286) );
na02f80 g760511 ( .a(n_19973), .b(n_19814), .o(n_19974) );
in01f80 g748451 ( .a(n_31783), .o(n_31835) );
na02f80 g775653 ( .a(n_5345), .b(n_5344), .o(n_5476) );
no02f80 g754702 ( .a(n_26231), .b(n_25440), .o(n_26311) );
ao12f80 g774250 ( .a(n_7029), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_16_), .o(n_7077) );
na02f80 g764828 ( .a(n_16356), .b(n_16355), .o(n_16357) );
in01f80 g769193 ( .a(n_12218), .o(n_12219) );
in01f80 g747346 ( .a(n_32663), .o(n_32664) );
in01f80 g780525 ( .a(n_1072), .o(n_1073) );
in01f80 newInst_2936 ( .a(newNet_802), .o(newNet_2936) );
no02f80 g748759 ( .a(n_31056), .b(n_29677), .o(n_31163) );
in01f80 g769363 ( .a(n_12084), .o(n_11889) );
na02f80 g739003 ( .a(n_41158), .b(n_40884), .o(n_41185) );
oa12f80 g780747 ( .a(n_435), .b(n_590), .c(n_589), .o(n_591) );
ao12f80 g771183 ( .a(n_9135), .b(n_9354), .c(n_9212), .o(n_9496) );
na02f80 g761323 ( .a(n_20177), .b(n_20220), .o(n_20810) );
in01f80 FE_RC_558_0 ( .a(n_30644), .o(FE_RN_169_0) );
in01f80 g778572 ( .a(n_2465), .o(n_2516) );
na02f80 g762203 ( .a(n_18735), .b(n_18620), .o(n_18736) );
oa22f80 g739713 ( .a(n_40526), .b(n_40390), .c(n_40527), .d(n_40391), .o(n_40560) );
no02f80 g741470 ( .a(n_38792), .b(n_38791), .o(n_38813) );
no02f80 g745438 ( .a(FE_OCP_RBN3698_n_35543), .b(n_35260), .o(n_35796) );
na02f80 g755126 ( .a(n_25374), .b(FE_OCP_RBN2366_n_24372), .o(n_25503) );
in01f80 newInst_2094 ( .a(newNet_2093), .o(newNet_2094) );
in01f80 g770252 ( .a(n_10754), .o(n_10795) );
no02f80 g756162 ( .a(n_24146), .b(n_24128), .o(n_24231) );
in01f80 g775488 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_11_), .o(n_5671) );
na02f80 g764826 ( .a(n_15598), .b(n_14524), .o(n_15695) );
in01f80 FE_RC_2602_0 ( .a(n_18052), .o(FE_RN_1080_0) );
in01f80 FE_OCPC3163_n_24117 ( .a(n_24117), .o(FE_OCPN3163_n_24117) );
no02f80 g755120 ( .a(n_25315), .b(n_24310), .o(n_25482) );
ao12f80 g772540 ( .a(n_7411), .b(n_8261), .c(n_7444), .o(n_8354) );
ao12f80 g766482 ( .a(n_14532), .b(n_14531), .c(n_14530), .o(n_15663) );
in01f80 g752381 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .o(n_27822) );
no02f80 g758259 ( .a(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n_22690) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_25_ ( .ck(newNet_2460), .d(n_32517), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_) );
no02f80 g760877 ( .a(n_19437), .b(n_19436), .o(n_19532) );
no02f80 g753735 ( .a(n_26449), .b(n_23353), .o(n_26596) );
na02f80 g738726 ( .a(n_41382), .b(n_41121), .o(n_41499) );
in01f80 newInst_780 ( .a(newNet_779), .o(newNet_780) );
na02f80 g775284 ( .a(n_5717), .b(n_4675), .o(n_5731) );
ao22s80 FE_RC_45_0 ( .a(n_2702), .b(n_2249), .c(n_2230), .d(n_1978), .o(n_2344) );
in01f80 g776578 ( .a(n_4411), .o(n_4412) );
in01f80 g768737 ( .a(n_12204), .o(n_12205) );
in01f80 FE_OCP_RBC2797_n_10106 ( .a(FE_OCP_RBN2796_n_10106), .o(FE_OCP_RBN2797_n_10106) );
na02f80 g752710 ( .a(n_28054), .b(n_28053), .o(n_28055) );
in01f80 g747679 ( .a(n_32190), .o(n_32191) );
in01f80 g773017 ( .a(n_7813), .o(n_7814) );
na02f80 g759310 ( .a(n_20862), .b(FE_OCP_RBN1715_n_20734), .o(n_20868) );
na02f80 g778981 ( .a(n_2187), .b(delay_add_ln22_unr2_stage2_stallmux_q_18_), .o(n_2232) );
na02f80 g780512 ( .a(n_1006), .b(n_882), .o(n_1074) );
no02f80 g764628 ( .a(n_15983), .b(n_15762), .o(n_15995) );
na02f80 g777154 ( .a(n_5368), .b(n_5330), .o(n_5331) );
in01f80 newInst_1483 ( .a(newNet_228), .o(newNet_1483) );
oa12f80 g758177 ( .a(n_21485), .b(n_21484), .c(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22785) );
na02f80 g755342 ( .a(n_24936), .b(n_24960), .o(n_25065) );
oa12f80 g767528 ( .a(n_12617), .b(n_12983), .c(n_12975), .o(n_13008) );
na02f80 g761342 ( .a(n_19909), .b(n_19930), .o(n_20558) );
in01f80 newInst_1561 ( .a(newNet_1560), .o(newNet_1561) );
oa12f80 g736453 ( .a(n_348), .b(n_43737), .c(FE_OFN2_n_43918), .o(n_43776) );
no02f80 g776817 ( .a(n_3978), .b(n_3891), .o(n_4152) );
no02f80 g771673 ( .a(n_9029), .b(n_44511), .o(n_10284) );
in01f80 g765897 ( .a(n_14854), .o(n_14875) );
no02f80 g750142 ( .a(n_29845), .b(n_29844), .o(n_29862) );
oa12f80 g772559 ( .a(n_8353), .b(n_8352), .c(n_8351), .o(n_8428) );
na02f80 g756742 ( .a(n_23479), .b(n_23444), .o(n_23693) );
na02f80 g741517 ( .a(n_38717), .b(n_38696), .o(n_38728) );
ao12f80 g739068 ( .a(n_40708), .b(n_41064), .c(n_40698), .o(n_41100) );
in01f80 FE_OCP_RBC1708_n_22150 ( .a(n_22150), .o(FE_OCP_RBN1708_n_22150) );
oa12f80 g775848 ( .a(n_4823), .b(n_5240), .c(n_4919), .o(n_5367) );
ao12f80 g743353 ( .a(n_37805), .b(n_37830), .c(n_46243), .o(n_37856) );
in01f80 g773829 ( .a(n_7101), .o(n_7072) );
oa22f80 g775843 ( .a(n_4903), .b(n_4182), .c(n_4858), .d(FE_OCP_RBN2727_n_4219), .o(n_5028) );
in01f80 g744372 ( .a(n_46215), .o(n_36854) );
oa22f80 FE_RC_3192_0 ( .a(n_10409), .b(FE_OCP_RBN3542_n_44575), .c(n_8732), .d(n_44563), .o(n_9020) );
in01f80 newInst_670 ( .a(newNet_669), .o(newNet_670) );
in01f80 g740437 ( .a(n_39804), .o(n_39805) );
no02f80 g741605 ( .a(n_38616), .b(n_38778), .o(n_38629) );
in01f80 FE_RC_4094_0 ( .a(n_22187), .o(FE_RN_1790_0) );
no02f80 g736954 ( .a(FE_OCPN1246_n_43120), .b(n_42953), .o(n_43510) );
oa22f80 g743567 ( .a(n_36398), .b(n_36238), .c(n_36399), .d(n_36239), .o(n_36449) );
ao12f80 g745220 ( .a(n_34571), .b(n_34570), .c(n_34569), .o(n_35644) );
no02f80 g766739 ( .a(n_13805), .b(n_13754), .o(n_13854) );
na02f80 g776689 ( .a(FE_OCP_RBN2584_n_3858), .b(n_2962), .o(n_3935) );
no02f80 g744026 ( .a(n_44256), .b(n_35598), .o(n_35625) );
na02f80 g771758 ( .a(n_10247), .b(n_10209), .o(n_10381) );
in01f80 g737299 ( .a(n_42922), .o(n_42923) );
in01f80 g746111 ( .a(n_35312), .o(n_35310) );
no02f80 g771741 ( .a(n_8969), .b(n_8968), .o(n_9006) );
ao22s80 FE_RC_1266_0 ( .a(delay_sub_ln23_0_unr25_stage9_stallmux_q), .b(n_38515), .c(n_38778), .d(FE_OCP_RBN2350_n_38515), .o(n_38579) );
in01f80 FE_OCP_RBC1365_n_29444 ( .a(n_29444), .o(FE_OCP_RBN1365_n_29444) );
in01f80 g779570 ( .a(n_1809), .o(n_1810) );
na02f80 g739117 ( .a(n_40979), .b(n_40805), .o(n_40996) );
no02f80 g755179 ( .a(n_25114), .b(n_23892), .o(n_25268) );
na02f80 g745244 ( .a(n_35725), .b(n_36049), .o(n_36124) );
no02f80 g742974 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n_37005) );
no02f80 g742311 ( .a(n_37822), .b(n_37821), .o(n_37833) );
no02f80 g743528 ( .a(n_36473), .b(n_36063), .o(n_36516) );
na02f80 g750103 ( .a(FE_OCP_RBN3566_n_29857), .b(FE_OCP_RBN1153_n_29053), .o(n_30051) );
na02f80 g761933 ( .a(n_19050), .b(n_18839), .o(n_19096) );
no02f80 g739447 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n_40770) );
na02f80 FE_RC_1232_0 ( .a(n_6513), .b(n_6380), .o(FE_RN_369_0) );
na02f80 g769693 ( .a(n_11316), .b(n_11187), .o(n_11361) );
na02f80 g762794 ( .a(n_18158), .b(n_18141), .o(n_18142) );
in01f80 FE_OCP_RBC2763_n_25732 ( .a(n_25732), .o(FE_OCP_RBN2763_n_25732) );
na02f80 g743158 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_5_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .o(n_36934) );
ao22s80 g751090 ( .a(n_30156), .b(n_29797), .c(n_30303), .d(n_30095), .o(n_30972) );
in01f80 fopt784014 ( .a(n_45748), .o(n_45747) );
ao12f80 g769008 ( .a(n_11840), .b(FE_OCP_RBN2120_n_45224), .c(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .o(n_12105) );
in01f80 FE_OCPC1754_n_7225 ( .a(FE_OCPN1753_n_7225), .o(FE_OCPN1754_n_7225) );
in01f80 g771613 ( .a(n_9243), .o(n_9338) );
in01f80 g775198 ( .a(n_6032), .o(n_6033) );
na02f80 g748991 ( .a(n_31031), .b(n_31007), .o(n_31103) );
in01f80 g764465 ( .a(n_16632), .o(n_16653) );
na02f80 g761190 ( .a(n_20051), .b(n_19991), .o(n_20052) );
no02f80 g770624 ( .a(n_10410), .b(n_10409), .o(n_10523) );
in01f80 g739980 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_), .o(n_40714) );
no02f80 g758247 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n_22842) );
in01f80 g746594 ( .a(n_34699), .o(n_34637) );
ao12f80 g768704 ( .a(n_12136), .b(FE_OCPN858_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .o(n_12416) );
no02f80 g751846 ( .a(n_29077), .b(n_28919), .o(n_29131) );
na02f80 g774826 ( .a(n_6228), .b(n_5790), .o(n_6338) );
na02f80 g757752 ( .a(n_22591), .b(n_22470), .o(n_22705) );
in01f80 newInst_2997 ( .a(newNet_2996), .o(newNet_2997) );
no02f80 g780824 ( .a(n_442), .b(n_452), .o(n_453) );
ao12f80 g751028 ( .a(n_28833), .b(n_28853), .c(n_28832), .o(n_28891) );
ao12f80 g775542 ( .a(n_5248), .b(n_5232), .c(n_5185), .o(n_5375) );
na02f80 g750161 ( .a(FE_OCP_RBN3567_n_29857), .b(n_29139), .o(n_30046) );
in01f80 g741094 ( .a(n_39364), .o(n_39365) );
no02f80 g759229 ( .a(n_21242), .b(n_45026), .o(n_21268) );
ao22s80 FE_RC_1300_0 ( .a(FE_OCP_RBN2863_n_39523), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .c(n_45840), .d(n_39523), .o(n_39592) );
oa22f80 g744010 ( .a(n_44223), .b(n_34593), .c(FE_OCPN3751_n_44222), .d(n_35648), .o(n_36316) );
ao12f80 g745132 ( .a(n_34377), .b(n_34725), .c(n_34344), .o(n_34824) );
in01f80 newInst_2957 ( .a(newNet_2956), .o(newNet_2957) );
no02f80 g754085 ( .a(n_26060), .b(n_26015), .o(n_26124) );
no02f80 g777291 ( .a(n_3564), .b(n_4662), .o(n_3612) );
ao12f80 g741699 ( .a(n_38102), .b(n_38506), .c(n_46416), .o(n_38519) );
in01f80 g775791 ( .a(FE_OCP_RBN2930_n_5221), .o(n_5265) );
na02f80 g768001 ( .a(n_12761), .b(n_12760), .o(n_12762) );
na02f80 g767643 ( .a(n_12938), .b(n_12937), .o(n_12939) );
in01f80 g751281 ( .a(n_30030), .o(n_29781) );
in01f80 g767153 ( .a(FE_OCPN1006_n_13962), .o(n_14420) );
in01f80 FE_OCP_RBC1377_n_20889 ( .a(FE_OCP_RBN1376_n_20889), .o(FE_OCP_RBN1377_n_20889) );
in01f80 g779118 ( .a(n_1976), .o(n_1977) );
no02f80 g763208 ( .a(n_17283), .b(n_17131), .o(n_17284) );
in01f80 g769079 ( .a(n_11754), .o(n_11755) );
in01f80 g740885 ( .a(n_39869), .o(n_39506) );
no02f80 g784600 ( .a(n_11118), .b(n_44498), .o(n_46423) );
ao22s80 g736323 ( .a(n_43812), .b(n_43318), .c(n_43811), .d(n_43319), .o(n_43857) );
in01f80 g768631 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_27_), .o(n_13013) );
in01f80 g743285 ( .a(n_36759), .o(n_36760) );
oa12f80 g775325 ( .a(n_5701), .b(n_5876), .c(n_5877), .o(n_5883) );
no02f80 g766815 ( .a(n_14349), .b(n_14382), .o(n_14430) );
in01f80 newInst_2548 ( .a(newNet_1082), .o(newNet_2548) );
na02f80 g771272 ( .a(n_9194), .b(n_9149), .o(n_9299) );
no02f80 g739281 ( .a(n_40811), .b(n_40777), .o(n_40778) );
in01f80 FE_OCP_RBC3857_FE_RN_779_0 ( .a(FE_RN_779_0), .o(FE_OCP_RBN3857_FE_RN_779_0) );
in01f80 g740336 ( .a(n_40407), .o(n_40408) );
in01f80 FE_OCPC1421_n_35611 ( .a(n_35611), .o(FE_OCPN1421_n_35611) );
ao22s80 g739128 ( .a(n_40964), .b(n_40955), .c(n_40925), .d(n_40954), .o(n_41028) );
oa22f80 g753657 ( .a(n_27132), .b(n_26926), .c(n_27133), .d(n_26927), .o(n_27247) );
na02f80 g743215 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .b(delay_add_ln22_unr23_stage9_stallmux_q_2_), .o(n_36886) );
no02f80 g758944 ( .a(n_21285), .b(FE_OCPN1414_n_19715), .o(n_21433) );
in01f80 g760216 ( .a(n_20311), .o(n_20269) );
no02f80 g747793 ( .a(n_33315), .b(n_33354), .o(n_33418) );
oa22f80 g740101 ( .a(FE_OCP_RBN3055_n_39913), .b(n_39508), .c(FE_OCP_RBN3722_n_39913), .d(n_39535), .o(n_40324) );
no02f80 g747724 ( .a(n_33625), .b(n_33671), .o(n_34042) );
in01f80 newInst_256 ( .a(newNet_255), .o(newNet_256) );
in01f80 g757216 ( .a(n_23140), .o(n_23141) );
in01f80 FE_OCP_RBC2281_n_29111 ( .a(n_29111), .o(FE_OCP_RBN2281_n_29111) );
no02f80 g748614 ( .a(n_31444), .b(n_31465), .o(n_31584) );
ao22s80 FE_RC_3786_0 ( .a(n_21619), .b(n_21686), .c(n_21588), .d(n_21710), .o(n_21816) );
na02f80 FE_RC_3261_0 ( .a(FE_RN_1306_0), .b(FE_RN_1439_0), .o(n_10215) );
na02f80 g784399 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .o(n_46211) );
in01f80 FE_OCP_RBC2791_n_9910 ( .a(n_9910), .o(FE_OCP_RBN2791_n_9910) );
in01f80 g777997 ( .a(n_3123), .o(n_3124) );
oa12f80 g746497 ( .a(n_33079), .b(n_33306), .c(n_33032), .o(n_33344) );
in01f80 g748890 ( .a(n_32459), .o(n_32412) );
no02f80 g763118 ( .a(n_17250), .b(n_17249), .o(n_17414) );
na02f80 g761479 ( .a(n_19647), .b(n_19793), .o(n_19826) );
in01f80 g738972 ( .a(n_41163), .o(n_41164) );
in01f80 FE_RC_672_0 ( .a(n_28291), .o(FE_RN_214_0) );
ao12f80 g778551 ( .a(FE_OCPN1234_n_2414), .b(n_2710), .c(n_2577), .o(n_3229) );
na02f80 g770692 ( .a(n_10181), .b(n_10112), .o(n_10307) );
na02f80 g750626 ( .a(n_29330), .b(n_29352), .o(n_29417) );
in01f80 g738809 ( .a(n_41382), .o(n_41478) );
in01f80 g764175 ( .a(n_16553), .o(n_16554) );
na02f80 g743907 ( .a(n_46249), .b(n_46211), .o(n_36941) );
in01f80 g767603 ( .a(n_13005), .o(n_12987) );
na02f80 g755813 ( .a(n_24426), .b(FE_OCP_DRV_N3154_n_24425), .o(n_24443) );
in01f80 FE_OCP_DRV_C1563_n_19665 ( .a(n_19665), .o(FE_OCP_DRV_N1563_n_19665) );
no02f80 g776253 ( .a(n_4824), .b(n_4919), .o(n_5194) );
in01f80 newInst_1220 ( .a(newNet_1219), .o(newNet_1220) );
in01f80 g740494 ( .a(n_39793), .o(n_39787) );
in01f80 g742371 ( .a(n_37810), .o(n_37811) );
na02f80 g747654 ( .a(n_33443), .b(n_33463), .o(n_33497) );
in01f80 g759015 ( .a(n_21285), .o(n_21286) );
na02f80 g745798 ( .a(n_34066), .b(FE_OCPN1856_n_33341), .o(n_34119) );
in01f80 g763088 ( .a(n_17292), .o(n_17349) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_4_ ( .ck(newNet_444), .d(n_27731), .o(delay_xor_ln22_unr18_stage7_stallmux_q_4_) );
na02f80 g740663 ( .a(n_39475), .b(n_39502), .o(n_39545) );
in01f80 g738692 ( .a(n_41560), .o(n_41602) );
oa12f80 g738304 ( .a(n_41522), .b(n_41648), .c(n_41524), .o(n_41888) );
in01f80 g778841 ( .a(n_3029), .o(n_3082) );
oa12f80 g741823 ( .a(n_38439), .b(n_38438), .c(n_38437), .o(n_38930) );
in01f80 FE_OCP_RBC2048_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2048_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01f80 FE_OCPC3185_FE_OCP_RBN1140_n_25816 ( .a(FE_OCP_RBN1140_n_25816), .o(FE_OCPN3185_FE_OCP_RBN1140_n_25816) );
na02f80 g755388 ( .a(n_24697), .b(n_24395), .o(n_24766) );
na02f80 g769234 ( .a(n_11556), .b(n_10542), .o(n_11753) );
na02f80 g750814 ( .a(n_30335), .b(n_30334), .o(n_30336) );
in01f80 FE_OCP_RBC3014_n_31117 ( .a(FE_OCP_RBN3009_n_31117), .o(FE_OCP_RBN3014_n_31117) );
na02f80 g769925 ( .a(n_11107), .b(n_11106), .o(n_11108) );
na02f80 g759445 ( .a(n_20939), .b(n_20968), .o(n_21121) );
in01f80 g739883 ( .a(n_40234), .o(n_40235) );
oa12f80 g736381 ( .a(n_338), .b(n_43815), .c(n_43918), .o(n_43860) );
in01f80 g748588 ( .a(n_31546), .o(n_31585) );
in01f80 FE_OCP_RBC2166_n_32892 ( .a(n_32892), .o(FE_OCP_RBN2166_n_32892) );
in01f80 newInst_3569 ( .a(newNet_1226), .o(newNet_3569) );
no02f80 g746903 ( .a(n_33015), .b(n_32082), .o(n_33061) );
in01f80 g762331 ( .a(n_18025), .o(n_18026) );
in01f80 newInst_3493 ( .a(newNet_3492), .o(newNet_3493) );
in01f80 newInst_2144 ( .a(newNet_2143), .o(newNet_2144) );
in01f80 g775304 ( .a(n_5980), .o(n_5981) );
no02f80 g766036 ( .a(n_14782), .b(n_14759), .o(n_14841) );
na02f80 g753946 ( .a(n_26221), .b(n_26220), .o(n_26298) );
no02f80 g755801 ( .a(n_24293), .b(n_22111), .o(n_24318) );
ao12f80 g754444 ( .a(n_25457), .b(n_25631), .c(n_25458), .o(n_25732) );
no02f80 g737383 ( .a(n_42784), .b(n_42444), .o(n_42821) );
na02f80 g773945 ( .a(n_6915), .b(delay_add_ln22_unr5_stage3_stallmux_q_6_), .o(n_7017) );
na02f80 g748121 ( .a(n_31807), .b(n_31783), .o(n_31875) );
na02f80 g737644 ( .a(n_42503), .b(n_42460), .o(n_42504) );
na02f80 g737774 ( .a(n_42558), .b(n_42581), .o(n_42627) );
na02f80 g737353 ( .a(n_42830), .b(n_42414), .o(n_42831) );
in01f80 fopt783451 ( .a(FE_OFN751_n_45003), .o(n_45012) );
no02f80 g774976 ( .a(n_6091), .b(n_6028), .o(n_6130) );
na02f80 g761495 ( .a(n_20086), .b(n_19758), .o(n_20082) );
no02f80 g769034 ( .a(FE_OCPN867_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .o(n_11975) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_12_ ( .ck(newNet_3078), .d(n_1137), .o(delay_add_ln22_unr2_stage2_stallmux_q_12_) );
no02f80 g743726 ( .a(n_37405), .b(n_46235), .o(n_37361) );
na02f80 g770496 ( .a(n_10319), .b(n_10096), .o(n_10330) );
no02f80 g737553 ( .a(n_42504), .b(n_42549), .o(n_42592) );
na02f80 g756562 ( .a(n_23636), .b(n_23635), .o(n_23637) );
in01f80 FE_RC_1616_0 ( .a(n_30882), .o(FE_RN_451_0) );
na02f80 FE_RC_511_0 ( .a(FE_RN_158_0), .b(n_28190), .o(n_28273) );
na02f80 g755698 ( .a(n_24485), .b(n_23283), .o(n_24592) );
in01f80 g753799 ( .a(n_26464), .o(n_26492) );
na02f80 g751167 ( .a(n_29909), .b(n_30082), .o(n_29943) );
in01f80 newInst_3031 ( .a(newNet_3030), .o(newNet_3031) );
na02f80 g746233 ( .a(n_33549), .b(n_33156), .o(n_33622) );
no02f80 g756903 ( .a(n_23367), .b(n_23366), .o(n_23368) );
in01f80 FE_OCP_RBC3091_n_11475 ( .a(n_11475), .o(FE_OCP_RBN3091_n_11475) );
na02f80 g740913 ( .a(n_39261), .b(n_39260), .o(n_39262) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_9_ ( .ck(newNet_1462), .d(n_31960), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_) );
no02f80 g759937 ( .a(n_21406), .b(n_21251), .o(n_21795) );
no02f80 g738244 ( .a(n_41940), .b(n_41925), .o(n_41926) );
in01f80 newInst_279 ( .a(newNet_278), .o(newNet_279) );
no02f80 g784790 ( .a(n_44268), .b(FE_OCPN3787_n_22156), .o(n_47278) );
oa22f80 FE_RC_1251_0 ( .a(FE_OCP_RBN2253_n_13017), .b(n_14157), .c(n_13469), .d(FE_OCP_RBN2454_n_14157), .o(n_14323) );
na02f80 g775361 ( .a(n_5528), .b(n_5480), .o(n_5609) );
no02f80 g759630 ( .a(n_20721), .b(n_20681), .o(n_20759) );
in01f80 FE_OCP_RBC2429_n_14018 ( .a(n_14018), .o(FE_OCP_RBN2429_n_14018) );
no02f80 g755435 ( .a(n_24802), .b(n_24752), .o(n_24805) );
na02f80 g770440 ( .a(n_10531), .b(n_10550), .o(n_10712) );
ao22s80 FE_RC_4121_0 ( .a(n_33250), .b(n_33656), .c(n_33251), .d(n_33655), .o(n_33728) );
in01f80 FE_OCP_RBC2481_n_14270 ( .a(n_14270), .o(FE_OCP_RBN2481_n_14270) );
na03f80 g740222 ( .a(n_39995), .b(n_39994), .c(n_39967), .o(n_40066) );
na02f80 g744459 ( .a(n_35455), .b(n_35341), .o(n_35486) );
in01f80 g739367 ( .a(n_41036), .o(n_41037) );
no02f80 g772860 ( .a(n_8017), .b(n_8016), .o(n_8052) );
in01f80 g746961 ( .a(n_32893), .o(n_32894) );
no02f80 g749742 ( .a(n_31317), .b(n_31345), .o(n_31390) );
in01f80 FE_OCP_RBC2375_n_8221 ( .a(FE_OCP_RBN2372_n_8221), .o(FE_OCP_RBN2375_n_8221) );
na02f80 g744872 ( .a(n_35115), .b(n_35094), .o(n_35192) );
ao12f80 g761624 ( .a(n_19096), .b(n_19496), .c(n_18623), .o(n_19613) );
oa12f80 g754466 ( .a(n_26793), .b(n_26713), .c(n_26541), .o(n_26794) );
in01f80 FE_OCP_RBC1152_n_29053 ( .a(n_29053), .o(FE_OCP_RBN1152_n_29053) );
in01f80 FE_OCPC936_n_42192 ( .a(FE_OCPN935_n_42192), .o(FE_OCPN936_n_42192) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_2_ ( .ck(newNet_626), .d(n_46373), .o(delay_xor_ln21_unr9_stage4_stallmux_q_2_) );
in01f80 FE_OCP_DRV_C1609_n_20146 ( .a(n_20146), .o(FE_OCP_DRV_N1609_n_20146) );
no02f80 g768024 ( .a(n_12914), .b(n_12965), .o(n_13080) );
in01f80 g742076 ( .a(n_38313), .o(n_38314) );
in01f80 FE_OCP_RBC2402_n_24638 ( .a(n_24638), .o(FE_OCP_RBN2402_n_24638) );
na02f80 g757996 ( .a(n_22763), .b(n_22696), .o(n_22764) );
in01f80 g745602 ( .a(n_34380), .o(n_34372) );
ao22s80 FE_RC_3774_0 ( .a(FE_RN_1656_0), .b(FE_OCP_RBN2367_n_24408), .c(n_23920), .d(n_24408), .o(n_24510) );
in01f80 g771587 ( .a(n_9077), .o(n_9078) );
no02f80 g749963 ( .a(n_29827), .b(n_29816), .o(n_29871) );
ao22s80 g736579 ( .a(n_43378), .b(n_43555), .c(n_43379), .d(n_43554), .o(n_43650) );
in01f80 g770179 ( .a(n_10845), .o(n_10846) );
in01f80 g761236 ( .a(FE_OCP_RBN1351_n_19148), .o(n_19164) );
ms00f80 cos_out_reg_27_ ( .ck(newNet_3706), .d(n_43909), .o(cos_out_27) );
in01f80 g777220 ( .a(n_3824), .o(n_3825) );
in01f80 g781327 ( .a(n_84), .o(n_152) );
no02f80 g740800 ( .a(n_39406), .b(n_39129), .o(n_39469) );
na02f80 g754828 ( .a(n_25948), .b(n_25341), .o(n_26007) );
in01f80 newInst_3555 ( .a(newNet_3554), .o(newNet_3555) );
na02f80 g757088 ( .a(n_23248), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_), .o(n_23290) );
in01f80 newInst_1045 ( .a(newNet_1044), .o(newNet_1045) );
in01f80 newInst_2905 ( .a(newNet_2904), .o(newNet_2905) );
in01f80 g751701 ( .a(n_28389), .o(n_28390) );
na02f80 g750646 ( .a(n_29376), .b(FE_OCPUNCON1802_n_29375), .o(n_29396) );
no02f80 g774961 ( .a(n_6135), .b(FE_OCP_RBN2924_n_5130), .o(n_6149) );
oa12f80 g751306 ( .a(FE_OCPN1034_n_28420), .b(n_28685), .c(n_28389), .o(n_28748) );
na02f80 g760481 ( .a(n_20516), .b(n_20515), .o(n_20517) );
ao12f80 g748987 ( .a(n_31454), .b(n_32295), .c(n_31511), .o(n_32316) );
in01f80 g765811 ( .a(n_15066), .o(n_15067) );
in01f80 g764342 ( .a(n_16394), .o(n_16424) );
na02f80 g741523 ( .a(n_38676), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38695) );
no02f80 g768921 ( .a(n_11761), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n_12121) );
na02f80 g752740 ( .a(n_27909), .b(n_27882), .o(n_27883) );
na02f80 g777308 ( .a(n_4182), .b(n_4537), .o(n_4612) );
in01f80 g759575 ( .a(n_20649), .o(n_20688) );
no02f80 FE_RC_1332_0 ( .a(FE_RN_393_0), .b(FE_RN_394_0), .o(FE_RN_395_0) );
in01f80 newInst_1818 ( .a(newNet_1817), .o(newNet_1818) );
in01f80 FE_OCP_RBC1208_n_16814 ( .a(FE_OCP_RBN1206_n_16814), .o(FE_OCP_RBN1208_n_16814) );
na02f80 g736829 ( .a(n_43515), .b(n_43126), .o(n_43551) );
in01f80 g739087 ( .a(n_41081), .o(n_41082) );
na02f80 g748819 ( .a(n_32482), .b(n_32481), .o(n_32725) );
in01f80 FE_OCP_RBC2738_n_15300 ( .a(n_15300), .o(FE_OCP_RBN2738_n_15300) );
in01f80 g756595 ( .a(n_23872), .o(n_23873) );
in01f80 g754392 ( .a(n_25812), .o(n_25843) );
in01f80 FE_OCP_RBC1842_n_20910 ( .a(n_20910), .o(FE_OCP_RBN1842_n_20910) );
no02f80 g755797 ( .a(n_24322), .b(n_21975), .o(n_24344) );
in01f80 g776147 ( .a(n_4942), .o(n_4986) );
in01f80 g747492 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n_32336) );
no02f80 g780896 ( .a(n_403), .b(n_402), .o(n_589) );
no02f80 g766794 ( .a(n_13661), .b(FE_OCPN860_n_12880), .o(n_13781) );
in01f80 FE_OCP_RBC3405_n_28597 ( .a(FE_OCP_RBN3404_n_28597), .o(FE_OCP_RBN3405_n_28597) );
na02f80 g737666 ( .a(FE_OCPN888_n_42367), .b(n_41992), .o(n_42659) );
no02f80 g776352 ( .a(n_4346), .b(n_4093), .o(n_4475) );
in01f80 FE_OCP_RBC3641_n_44490 ( .a(FE_OCP_RBN3637_n_44490), .o(FE_OCP_RBN3641_n_44490) );
no02f80 g744643 ( .a(n_35326), .b(n_35281), .o(n_35327) );
in01f80 g757588 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .o(n_23605) );
in01f80 g753166 ( .a(n_27542), .o(n_27543) );
in01f80 newInst_207 ( .a(newNet_206), .o(newNet_207) );
oa12f80 g768349 ( .a(n_12054), .b(n_12460), .c(n_11896), .o(n_12545) );
oa12f80 g740814 ( .a(n_39435), .b(n_39434), .c(n_39433), .o(n_39917) );
na02f80 g757247 ( .a(n_23494), .b(n_23183), .o(n_23533) );
in01f80 FE_OCPC979_n_21973 ( .a(FE_OCPN978_n_21973), .o(FE_OCPN979_n_21973) );
in01f80 FE_OCP_RBC2364_n_24372 ( .a(n_24372), .o(FE_OCP_RBN2364_n_24372) );
in01f80 FE_OCP_RBC2156_n_1602 ( .a(n_1602), .o(FE_OCP_RBN2156_n_1602) );
in01f80 g759655 ( .a(n_20555), .o(n_20614) );
no02f80 g765044 ( .a(n_16103), .b(n_15972), .o(n_16104) );
in01f80 g737568 ( .a(n_42290), .o(n_42264) );
ao12f80 g752008 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .b(n_28044), .c(FE_OCPN878_n_44734), .o(n_28045) );
na02f80 g774002 ( .a(n_6845), .b(n_6596), .o(n_6913) );
no02f80 g772760 ( .a(n_8095), .b(n_8177), .o(n_8259) );
in01f80 g767674 ( .a(n_13351), .o(n_13352) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_4_ ( .ck(newNet_1003), .d(n_16873), .o(delay_xor_ln21_unr12_stage5_stallmux_q_4_) );
ao22s80 g784420 ( .a(n_36762), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_46232) );
in01f80 g753990 ( .a(n_27031), .o(n_27032) );
no02f80 g763071 ( .a(n_17414), .b(n_17132), .o(n_17489) );
in01f80 g745775 ( .a(n_34394), .o(n_34395) );
in01f80 newInst_2184 ( .a(newNet_2183), .o(newNet_2184) );
in01f80 g765225 ( .a(n_15836), .o(n_15932) );
no02f80 g767548 ( .a(n_12983), .b(n_12638), .o(n_12984) );
no02f80 g763190 ( .a(n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(n_17436) );
na02f80 g758609 ( .a(n_21816), .b(n_20205), .o(n_21905) );
na02f80 FE_RC_4147_0 ( .a(n_16900), .b(FE_RN_1802_0), .o(FE_RN_1803_0) );
in01f80 newInst_1662 ( .a(newNet_1661), .o(newNet_1662) );
na02f80 g761439 ( .a(n_18797), .b(FE_OFN778_n_17093), .o(n_18831) );
in01f80 g743581 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(n_36951) );
in01f80 newInst_2480 ( .a(newNet_1517), .o(newNet_2480) );
no02f80 g774356 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_10_), .o(n_6747) );
na02f80 g755165 ( .a(n_25551), .b(n_24639), .o(n_25618) );
in01f80 g738684 ( .a(n_41614), .o(n_41561) );
in01f80 FE_OCPC1736_n_37877 ( .a(FE_OCPN1735_n_37877), .o(FE_OCPN1736_n_37877) );
in01f80 g777697 ( .a(n_3535), .o(n_3536) );
in01f80 g763956 ( .a(n_16609), .o(n_16626) );
in01f80 g752601 ( .a(n_27622), .o(n_27607) );
in01f80 g744905 ( .a(n_34960), .o(n_34983) );
in01f80 newInst_817 ( .a(newNet_804), .o(newNet_817) );
in01f80 g766979 ( .a(n_13577), .o(n_13593) );
in01f80 FE_RC_1056_0 ( .a(n_24099), .o(FE_RN_310_0) );
oa12f80 g755229 ( .a(n_25041), .b(n_25067), .c(n_24933), .o(n_25178) );
oa12f80 g781119 ( .a(n_161), .b(n_224), .c(n_111), .o(n_233) );
in01f80 g760563 ( .a(n_19891), .o(n_19892) );
in01f80 newInst_301 ( .a(newNet_300), .o(newNet_301) );
na02f80 g775293 ( .a(n_5810), .b(n_4759), .o(n_5857) );
na02f80 g767794 ( .a(n_12823), .b(n_13013), .o(n_13014) );
no02f80 g751693 ( .a(n_28382), .b(n_28006), .o(n_28437) );
na02f80 g739969 ( .a(n_40022), .b(n_40045), .o(n_40086) );
oa12f80 g748338 ( .a(n_31522), .b(FE_OCPN1052_n_31674), .c(FE_OCPN1418_n_31504), .o(n_31916) );
na02f80 g738348 ( .a(n_41753), .b(n_41645), .o(n_41754) );
ao12f80 g752702 ( .a(n_28615), .b(n_27993), .c(n_27899), .o(n_28202) );
no02f80 g780840 ( .a(n_589), .b(n_434), .o(n_587) );
ao12f80 g750734 ( .a(n_30307), .b(n_30306), .c(n_29882), .o(n_30337) );
in01f80 FE_OCP_RBC2191_n_28597 ( .a(n_28597), .o(FE_OCP_RBN2191_n_28597) );
no02f80 FE_RC_4038_0 ( .a(FE_RN_1753_0), .b(n_26442), .o(FE_RN_1754_0) );
no02f80 g774315 ( .a(n_6551), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6552) );
na02f80 g773586 ( .a(n_7348), .b(n_7250), .o(n_7383) );
no02f80 g772043 ( .a(n_8821), .b(n_8820), .o(n_8822) );
in01f80 newInst_606 ( .a(newNet_605), .o(newNet_606) );
no02f80 g756803 ( .a(n_23349), .b(n_23215), .o(n_23409) );
na02f80 g760196 ( .a(FE_OCP_RBN3617_n_20249), .b(n_20124), .o(n_20604) );
na02f80 g761270 ( .a(n_19678), .b(n_19787), .o(n_19959) );
na02f80 g752509 ( .a(n_27691), .b(n_27466), .o(n_27709) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_18_ ( .ck(newNet_571), .d(n_17769), .o(delay_xor_ln22_unr12_stage5_stallmux_q_18_) );
na02f80 FE_RC_2942_0 ( .a(FE_OCP_RBN3621_n_15135), .b(n_15341), .o(FE_RN_1283_0) );
in01f80 newInst_3275 ( .a(newNet_2960), .o(newNet_3275) );
in01f80 g738711 ( .a(n_41803), .o(n_41804) );
in01f80 g767586 ( .a(n_12983), .o(n_12944) );
na02f80 g749674 ( .a(n_31259), .b(n_31294), .o(n_31295) );
oa12f80 g780253 ( .a(n_1105), .b(n_1104), .c(n_1103), .o(n_1133) );
no02f80 g765510 ( .a(n_15441), .b(n_15482), .o(n_15483) );
in01f80 FE_OCP_RBC2757_FE_RN_722_0 ( .a(FE_RN_722_0), .o(FE_OCP_RBN2757_FE_RN_722_0) );
na02f80 g737020 ( .a(n_43230), .b(n_42750), .o(n_43488) );
in01f80 newInst_3322 ( .a(newNet_2115), .o(newNet_3322) );
no02f80 g750070 ( .a(n_29896), .b(n_29262), .o(n_30244) );
no02f80 g773178 ( .a(n_7612), .b(n_7611), .o(n_7613) );
no02f80 g750064 ( .a(n_29869), .b(n_29161), .o(n_30172) );
in01f80 newInst_3151 ( .a(newNet_118), .o(newNet_3151) );
in01f80 newInst_1325 ( .a(newNet_1324), .o(newNet_1325) );
in01f80 g752372 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_31_), .o(n_27824) );
no02f80 g754226 ( .a(n_25957), .b(FE_OFN737_n_22641), .o(n_25991) );
in01f80 FE_OCP_RBC2192_n_28597 ( .a(FE_OCP_RBN2191_n_28597), .o(FE_OCP_RBN2192_n_28597) );
in01f80 g774338 ( .a(n_7121), .o(n_7122) );
in01f80 newInst_1030 ( .a(newNet_1029), .o(newNet_1030) );
in01f80 FE_RC_3102_0 ( .a(FE_RN_1372_0), .o(n_21397) );
oa22f80 g765743 ( .a(n_14884), .b(n_14809), .c(n_14885), .d(n_14810), .o(n_14985) );
na02f80 g759046 ( .a(n_21128), .b(n_45024), .o(n_21287) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_31_ ( .ck(newNet_1695), .d(n_22550), .o(n_22641) );
in01f80 FE_OCP_RBC3021_n_39942 ( .a(n_39942), .o(FE_OCP_RBN3021_n_39942) );
in01f80 g779248 ( .a(n_1889), .o(n_1872) );
in01f80 newInst_1944 ( .a(newNet_1943), .o(newNet_1944) );
no02f80 g744684 ( .a(n_35156), .b(n_35152), .o(n_35237) );
in01f80 g767007 ( .a(n_14486), .o(n_14487) );
in01f80 FE_OCP_RBC2327_n_29378 ( .a(FE_OCP_RBN2326_n_29378), .o(FE_OCP_RBN2327_n_29378) );
in01f80 g778128 ( .a(n_2950), .o(n_2951) );
in01f80 FE_OCP_RBC2460_n_2818 ( .a(n_2818), .o(FE_OCP_RBN2460_n_2818) );
oa22f80 FE_RC_3428_0 ( .a(n_31825), .b(n_32172), .c(n_31826), .d(n_32195), .o(n_32290) );
in01f80 g741506 ( .a(n_38748), .o(n_38749) );
in01f80 g746100 ( .a(n_33833), .o(n_33828) );
no02f80 g758235 ( .a(n_22608), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22693) );
in01f80 g745397 ( .a(n_35958), .o(n_36021) );
in01f80 g740411 ( .a(n_40054), .o(n_40132) );
in01f80 newInst_2596 ( .a(newNet_2595), .o(newNet_2596) );
in01f80 g759964 ( .a(n_21334), .o(n_21407) );
ao12f80 g761886 ( .a(n_18820), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n_18848) );
na02f80 g759906 ( .a(n_21406), .b(n_20894), .o(n_21622) );
no03m80 FE_RC_2456_0 ( .a(n_13700), .b(n_13349), .c(n_13286), .o(FE_RN_984_0) );
na02f80 g737274 ( .a(n_42881), .b(n_42760), .o(n_42904) );
no02f80 g754439 ( .a(n_25654), .b(FE_OCPN1259_n_25353), .o(n_25704) );
no02f80 FE_RC_1618_0 ( .a(FE_RN_452_0), .b(n_30884), .o(n_46956) );
na03f80 g742409 ( .a(n_37754), .b(n_37717), .c(n_37622), .o(n_37724) );
no02f80 g746541 ( .a(n_34805), .b(n_34809), .o(n_34841) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_19_ ( .ck(newNet_3150), .d(n_40488), .o(delay_add_ln22_unr27_stage10_stallmux_q_19_) );
in01f80 newInst_1402 ( .a(newNet_1401), .o(newNet_1402) );
na02f80 g767448 ( .a(n_13494), .b(n_13201), .o(n_13503) );
oa12f80 g745052 ( .a(n_34718), .b(n_34717), .c(n_34716), .o(n_35785) );
in01f80 g743048 ( .a(n_36954), .o(n_37067) );
no02f80 g739099 ( .a(n_41060), .b(n_40918), .o(n_41061) );
no02f80 g738599 ( .a(n_41364), .b(n_40929), .o(n_41379) );
in01f80 g770400 ( .a(n_10537), .o(n_10538) );
na02f80 g775341 ( .a(n_6001), .b(n_5930), .o(n_5966) );
oa12f80 g765072 ( .a(n_15528), .b(n_15527), .c(n_15526), .o(n_15603) );
no02f80 g756736 ( .a(n_23500), .b(FE_RN_142_0), .o(n_23501) );
in01f80 g758105 ( .a(n_22300), .o(n_22301) );
na02f80 g738397 ( .a(n_41622), .b(n_41674), .o(n_41675) );
oa12f80 g747263 ( .a(n_33296), .b(n_45753), .c(n_33840), .o(n_33913) );
ao22s80 g774245 ( .a(n_6506), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .o(n_6601) );
in01f80 FE_RC_1744_0 ( .a(n_12275), .o(FE_RN_489_0) );
na02f80 g780503 ( .a(n_842), .b(n_768), .o(n_799) );
in01f80 g772434 ( .a(n_8594), .o(n_8652) );
na02f80 g769083 ( .a(n_11753), .b(n_11675), .o(n_11810) );
oa22f80 g742034 ( .a(FE_OCP_RBN3441_n_37945), .b(n_37589), .c(FE_OCP_RBN3445_n_37945), .d(n_37619), .o(n_38349) );
in01f80 FE_RC_4219_0 ( .a(FE_OCP_RBN1324_n_29056), .o(FE_RN_1848_0) );
na02f80 g753154 ( .a(n_27298), .b(n_27413), .o(n_27525) );
no02f80 g774288 ( .a(n_6765), .b(n_6764), .o(n_6766) );
in01f80 FE_OCP_RBC3061_FE_RN_640_0 ( .a(FE_RN_640_0), .o(FE_OCP_RBN3061_FE_RN_640_0) );
oa12f80 g746402 ( .a(n_33289), .b(n_33429), .c(n_33246), .o(n_33471) );
oa12f80 g779352 ( .a(n_1707), .b(n_1585), .c(delay_add_ln22_unr2_stage2_stallmux_q_1_), .o(n_2343) );
no02f80 g770701 ( .a(n_10223), .b(n_10031), .o(n_10261) );
no02f80 g746779 ( .a(n_32948), .b(n_33252), .o(n_33274) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_27_ ( .ck(newNet_1208), .d(n_6286), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_) );
na02f80 g769345 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .o(n_11601) );
na02f80 g760233 ( .a(FE_OCPN1261_n_20242), .b(FE_OCP_RBN3831_n_19204), .o(n_20433) );
no02f80 g756033 ( .a(FE_OCP_RBN2525_n_24902), .b(n_24957), .o(n_25029) );
na02f80 g774041 ( .a(n_7172), .b(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .o(n_7179) );
oa22f80 g751520 ( .a(n_28817), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .c(FE_OCP_RBN2218_FE_OCPN950_n_28595), .d(n_27623), .o(n_28970) );
na02f80 g756626 ( .a(n_23572), .b(n_22773), .o(n_23707) );
na02f80 g743345 ( .a(n_36656), .b(n_36750), .o(n_36695) );
no02f80 g751461 ( .a(n_28565), .b(n_28645), .o(n_28679) );
na02f80 FE_RC_2524_0 ( .a(FE_RN_1028_0), .b(n_40893), .o(n_41120) );
na02f80 g766537 ( .a(n_13954), .b(n_13422), .o(n_14060) );
na02f80 g764550 ( .a(n_16044), .b(n_16079), .o(n_16220) );
na02f80 g742968 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n_37010) );
no02f80 g746738 ( .a(n_33203), .b(n_33109), .o(n_33234) );
ao12f80 g756329 ( .a(n_23577), .b(n_23930), .c(n_23631), .o(n_23949) );
no02f80 g767556 ( .a(n_13005), .b(n_13004), .o(n_13006) );
na02f80 g764102 ( .a(FE_OCP_RBN3798_delay_xor_ln22_unr12_stage5_stallmux_q_0_), .b(n_44365), .o(n_16745) );
na02f80 g771238 ( .a(n_9659), .b(n_9613), .o(n_9660) );
na02f80 g754909 ( .a(n_25542), .b(n_24717), .o(n_25591) );
na02f80 g765147 ( .a(n_15189), .b(n_15236), .o(n_15310) );
in01f80 newInst_1847 ( .a(newNet_1846), .o(newNet_1847) );
no02f80 g753201 ( .a(n_27087), .b(n_46962), .o(n_27145) );
na02f80 g754931 ( .a(n_24245), .b(n_25270), .o(n_25357) );
no02f80 g769783 ( .a(n_11208), .b(n_11047), .o(n_11240) );
na02f80 g765137 ( .a(n_15311), .b(FE_OCP_RBN3660_n_15233), .o(n_15344) );
oa12f80 g738091 ( .a(n_41677), .b(n_42071), .c(n_41586), .o(n_42091) );
in01f80 g739595 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_2_), .o(n_40615) );
in01f80 g773147 ( .a(n_7716), .o(n_7697) );
in01f80 FE_OCPC1050_n_4459 ( .a(FE_OCPN1049_n_4459), .o(FE_OCPN1050_n_4459) );
in01f80 g771354 ( .a(n_9351), .o(n_9352) );
na02f80 g764261 ( .a(n_16424), .b(n_16364), .o(n_16462) );
in01f80 FE_OCPC3794_FE_RN_1789_0 ( .a(FE_RN_1789_0), .o(FE_OCPN3794_FE_RN_1789_0) );
no03m80 FE_RC_4171_0 ( .a(n_18343), .b(n_18319), .c(n_18759), .o(n_18760) );
na02f80 g743058 ( .a(n_37171), .b(n_37175), .o(n_37204) );
oa22f80 g773227 ( .a(n_44828), .b(n_45889), .c(n_44829), .d(n_7193), .o(n_7957) );
na02f80 g776576 ( .a(n_4434), .b(n_4433), .o(n_4480) );
na02f80 g777273 ( .a(n_4759), .b(n_3265), .o(n_4873) );
in01f80 g766099 ( .a(n_14659), .o(n_14660) );
in01f80 g760381 ( .a(n_20205), .o(n_20206) );
no02f80 g767479 ( .a(n_13462), .b(n_13166), .o(n_13494) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_3_ ( .ck(newNet_2250), .d(n_39848), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_3_) );
in01f80 fopt782738 ( .a(n_17685), .o(n_44147) );
in01f80 g775247 ( .a(n_6116), .o(n_6117) );
in01f80 g749772 ( .a(n_31369), .o(n_31370) );
no02f80 g743104 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .o(n_37048) );
na02f80 g776186 ( .a(n_4887), .b(n_4886), .o(n_4966) );
in01f80 FE_RC_2763_0 ( .a(FE_RN_1177_0), .o(n_9182) );
in01f80 g740530 ( .a(n_39674), .o(n_39687) );
no02f80 g746001 ( .a(n_35246), .b(n_35245), .o(n_35247) );
na02f80 g773840 ( .a(n_7125), .b(n_7011), .o(n_7209) );
in01f80 g775445 ( .a(n_5679), .o(n_5680) );
in01f80 newInst_3009 ( .a(newNet_2576), .o(newNet_3009) );
no02f80 g768289 ( .a(n_12518), .b(n_12396), .o(n_12571) );
in01f80 newInst_708 ( .a(newNet_371), .o(newNet_708) );
oa12f80 g778148 ( .a(n_2823), .b(FE_OCP_RBN3490_n_3390), .c(FE_OCP_RBN2292_n_2438), .o(n_2850) );
oa12f80 g773117 ( .a(n_7891), .b(n_8362), .c(n_7828), .o(n_8648) );
in01f80 g767616 ( .a(n_13136), .o(n_13137) );
no02f80 g737436 ( .a(n_42705), .b(n_42494), .o(n_42738) );
oa12f80 g761626 ( .a(n_19522), .b(n_19521), .c(n_19520), .o(n_19844) );
in01f80 g737699 ( .a(n_42222), .o(n_42253) );
na02f80 g749364 ( .a(n_30349), .b(n_30582), .o(n_30655) );
in01f80 FE_OCP_RBC2321_n_2638 ( .a(n_2638), .o(FE_OCP_RBN2321_n_2638) );
na02f80 g741592 ( .a(n_38626), .b(n_38623), .o(n_38651) );
in01f80 newInst_115 ( .a(newNet_114), .o(newNet_115) );
oa12f80 g756958 ( .a(n_23327), .b(n_23324), .c(n_23326), .o(n_23404) );
in01f80 g740705 ( .a(n_39584), .o(n_40005) );
na02f80 g769839 ( .a(n_11150), .b(n_11102), .o(n_11191) );
na02f80 g773187 ( .a(n_7817), .b(n_7888), .o(n_7854) );
no02f80 g759521 ( .a(n_20958), .b(n_20931), .o(n_21110) );
na02f80 g763797 ( .a(FE_OCP_RBN1678_n_44847), .b(n_44365), .o(n_16988) );
in01f80 g749245 ( .a(n_30806), .o(n_30807) );
na02f80 g743172 ( .a(n_36943), .b(n_36944), .o(n_36945) );
na02f80 g744469 ( .a(n_35483), .b(FE_OCP_DRV_N1580_n_35482), .o(n_35515) );
na02f80 g754953 ( .a(FE_OCPN985_n_25210), .b(n_24420), .o(n_25383) );
in01f80 FE_RC_3840_0 ( .a(n_17040), .o(FE_RN_1673_0) );
ms00f80 cos_out_reg_25_ ( .ck(newNet_3710), .d(n_43886), .o(cos_out_25) );
no02f80 g763007 ( .a(FE_OCP_RBN3213_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .o(n_17684) );
no02f80 g784067 ( .a(n_45812), .b(n_831), .o(n_45813) );
no02f80 g773685 ( .a(n_7311), .b(n_7788), .o(n_7312) );
in01f80 g768589 ( .a(n_12262), .o(n_12263) );
ao12f80 g766107 ( .a(n_14407), .b(n_14483), .c(n_14368), .o(n_14582) );
na02f80 g761158 ( .a(n_19143), .b(n_19142), .o(n_19144) );
in01f80 g769243 ( .a(n_11658), .o(n_11647) );
na02f80 FE_RC_3313_0 ( .a(FE_RN_553_0), .b(FE_RN_1458_0), .o(n_14092) );
no02f80 g750783 ( .a(n_29144), .b(n_28680), .o(n_29166) );
in01f80 g739626 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n_40607) );
oa12f80 g751018 ( .a(n_29909), .b(n_30037), .c(n_30083), .o(n_30100) );
na02f80 g759190 ( .a(n_21416), .b(n_21415), .o(n_21417) );
oa12f80 g775938 ( .a(n_4474), .b(n_4605), .c(n_4411), .o(n_4776) );
no02f80 g752999 ( .a(n_27299), .b(n_27294), .o(n_27427) );
oa12f80 g745030 ( .a(n_34537), .b(n_34858), .c(n_34857), .o(n_34875) );
in01f80 g753502 ( .a(n_27559), .o(n_27560) );
oa12f80 g741777 ( .a(n_38323), .b(n_38389), .c(n_38373), .o(n_38502) );
in01f80 g775051 ( .a(n_6171), .o(n_6172) );
in01f80 FE_OCP_RBC2365_n_24372 ( .a(n_24372), .o(FE_OCP_RBN2365_n_24372) );
no02f80 FE_RC_2719_0 ( .a(FE_RN_1146_0), .b(n_8410), .o(FE_RN_1148_0) );
na02f80 g764364 ( .a(n_16200), .b(n_16226), .o(n_16287) );
na02f80 g780184 ( .a(n_1128), .b(n_848), .o(n_1170) );
ao12f80 g763161 ( .a(n_17289), .b(FE_OCP_RBN3210_n_44365), .c(delay_xor_ln21_unr12_stage5_stallmux_q_5_), .o(n_17345) );
in01f80 g776198 ( .a(n_4938), .o(n_4939) );
in01f80 FE_OCP_RBC2987_n_35539 ( .a(FE_OCP_RBN3698_n_35543), .o(FE_OCP_RBN2987_n_35539) );
no02f80 g760934 ( .a(n_19457), .b(n_19456), .o(n_19458) );
na02f80 g780561 ( .a(n_779), .b(n_828), .o(n_869) );
no02f80 g752805 ( .a(n_27992), .b(n_27789), .o(n_28588) );
in01f80 g750563 ( .a(n_29473), .o(n_29474) );
na02f80 FE_RC_2322_0 ( .a(n_39652), .b(n_39637), .o(FE_RN_883_0) );
no02f80 g753554 ( .a(n_26756), .b(n_26389), .o(n_26781) );
na02f80 g781040 ( .a(sin_out_11), .b(FE_OFN3_n_43918), .o(n_349) );
na02f80 g737039 ( .a(n_43230), .b(n_42804), .o(n_43486) );
no02f80 FE_RC_4045_0 ( .a(n_21319), .b(n_21540), .o(n_21573) );
oa12f80 g742262 ( .a(FE_OCP_RBN2240_n_44881), .b(n_37697), .c(n_38047), .o(n_38199) );
oa12f80 g768844 ( .a(n_11933), .b(n_12088), .c(n_12011), .o(n_12095) );
in01f80 FE_OCP_RBC3023_n_39942 ( .a(n_39942), .o(FE_OCP_RBN3023_n_39942) );
na02f80 g742709 ( .a(n_37355), .b(n_37354), .o(n_37356) );
na02f80 g762315 ( .a(n_18080), .b(n_18057), .o(n_18058) );
no02f80 g757228 ( .a(n_23175), .b(n_23176), .o(n_23177) );
in01f80 g749983 ( .a(n_31311), .o(n_31530) );
na02f80 g769985 ( .a(n_10888), .b(n_10877), .o(n_10992) );
na02f80 g749253 ( .a(n_30733), .b(FE_OCPN1486_n_27315), .o(n_30768) );
na02f80 g747731 ( .a(n_33417), .b(n_33312), .o(n_33629) );
oa22f80 FE_RC_195_0 ( .a(n_17318), .b(n_17516), .c(n_17317), .d(n_17559), .o(n_17723) );
no02f80 g778114 ( .a(n_2966), .b(n_2928), .o(n_3040) );
in01f80 g777921 ( .a(n_4211), .o(n_3226) );
na02f80 g771972 ( .a(n_44498), .b(n_9913), .o(n_9953) );
in01f80 newInst_2465 ( .a(newNet_2464), .o(newNet_2465) );
no02f80 g773161 ( .a(n_7730), .b(n_7771), .o(n_7849) );
na02f80 g751174 ( .a(n_29944), .b(n_29942), .o(n_30126) );
in01f80 FE_OCP_RBC2472_n_8664 ( .a(n_8664), .o(FE_OCP_RBN2472_n_8664) );
oa22f80 g749012 ( .a(n_32269), .b(n_31537), .c(n_32295), .d(n_31538), .o(n_32341) );
na02f80 g746489 ( .a(n_34891), .b(n_34666), .o(n_34940) );
in01f80 g777894 ( .a(n_3236), .o(n_3192) );
no02f80 g748660 ( .a(n_31462), .b(n_31439), .o(n_31486) );
in01f80 FE_OCP_RBC3386_n_33108 ( .a(FE_OCP_RBN3385_n_33108), .o(FE_OCP_RBN3386_n_33108) );
in01f80 fopt783240 ( .a(n_44800), .o(n_44798) );
no02f80 g757238 ( .a(n_23494), .b(n_23053), .o(n_23525) );
in01f80 fopt783586 ( .a(n_45216), .o(n_45217) );
in01f80 g749486 ( .a(n_31911), .o(n_31941) );
no02f80 g738544 ( .a(n_41420), .b(n_41157), .o(n_41595) );
no02f80 g763355 ( .a(n_17192), .b(n_17084), .o(n_17126) );
ao12f80 g762052 ( .a(n_18590), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n_18631) );
in01f80 FE_OCPC3793_n_31804 ( .a(FE_OCPN3792_n_31804), .o(FE_OCPN3793_n_31804) );
no02f80 g759693 ( .a(n_20546), .b(n_20589), .o(n_20727) );
in01f80 FE_OCP_RBC3127_n_43752 ( .a(n_43752), .o(FE_OCP_RBN3127_n_43752) );
in01f80 FE_OCP_RBC1722_n_21004 ( .a(n_21004), .o(FE_OCP_RBN1722_n_21004) );
in01f80 g755561 ( .a(n_24618), .o(n_24619) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_5_ ( .ck(newNet_406), .d(n_32541), .o(delay_xor_ln22_unr21_stage8_stallmux_q_5_) );
in01f80 newInst_976 ( .a(newNet_975), .o(newNet_976) );
na02f80 g771377 ( .a(n_9370), .b(FE_OCPN903_n_44581), .o(n_9447) );
ao12f80 g740726 ( .a(n_39043), .b(n_39532), .c(n_38988), .o(n_39566) );
in01f80 g748374 ( .a(n_31501), .o(n_31560) );
ao12f80 g749625 ( .a(n_29986), .b(n_30250), .c(n_29920), .o(n_30461) );
in01f80 FE_OCP_RBC3007_n_31117 ( .a(FE_OCP_RBN3701_n_31064), .o(FE_OCP_RBN3007_n_31117) );
oa12f80 g775018 ( .a(n_5287), .b(n_6076), .c(n_5186), .o(n_6160) );
no02f80 g737544 ( .a(n_42377), .b(n_42317), .o(n_42378) );
in01f80 g760721 ( .a(n_21835), .o(n_20255) );
in01f80 g747987 ( .a(n_33072), .o(n_33073) );
na02f80 FE_RC_2013_0 ( .a(FE_RN_663_0), .b(n_20184), .o(FE_RN_664_0) );
in01f80 g779068 ( .a(n_2056), .o(n_2057) );
na02f80 g767645 ( .a(n_13156), .b(n_13192), .o(n_13700) );
na02f80 g759557 ( .a(n_20873), .b(n_19099), .o(n_20957) );
no02f80 g761481 ( .a(n_19649), .b(n_19760), .o(n_19828) );
in01f80 g768421 ( .a(n_12438), .o(n_12439) );
in01f80 newInst_948 ( .a(newNet_604), .o(newNet_948) );
na02f80 g759892 ( .a(n_20295), .b(n_45065), .o(n_20319) );
in01f80 g760299 ( .a(n_20953), .o(n_20954) );
in01f80 newInst_1434 ( .a(newNet_691), .o(newNet_1434) );
in01f80 newInst_3678 ( .a(newNet_3677), .o(newNet_3678) );
na02f80 g741034 ( .a(n_39204), .b(n_39251), .o(n_39276) );
na02f80 g769828 ( .a(n_11082), .b(n_10986), .o(n_11130) );
in01f80 g743459 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .o(n_36564) );
in01f80 g766231 ( .a(n_14503), .o(n_14504) );
na02f80 g761069 ( .a(n_19153), .b(n_19044), .o(n_19181) );
ao12f80 g765102 ( .a(n_15233), .b(n_15243), .c(n_15311), .o(n_15382) );
ao12f80 g738451 ( .a(n_41623), .b(n_41660), .c(n_41180), .o(n_41968) );
in01f80 newInst_1825 ( .a(newNet_1824), .o(newNet_1825) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_18_ ( .ck(newNet_1326), .d(n_1234), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_) );
na02f80 g768371 ( .a(n_12506), .b(n_12480), .o(n_12520) );
no02f80 g771362 ( .a(FE_OCP_RBN2564_FE_RN_1125_0), .b(n_9163), .o(n_9348) );
na02f80 g769843 ( .a(n_11128), .b(FE_OCP_RBN2769_n_9892), .o(n_11195) );
no02f80 g742904 ( .a(n_37126), .b(n_37471), .o(n_37124) );
na02f80 g775237 ( .a(n_5950), .b(n_5949), .o(n_5951) );
no02f80 g754565 ( .a(n_26548), .b(n_26604), .o(n_26573) );
oa12f80 g764769 ( .a(n_16360), .b(n_16359), .c(n_16358), .o(n_16414) );
oa12f80 g742163 ( .a(n_38300), .b(FE_OCP_RBN2241_n_44881), .c(n_38298), .o(n_38415) );
oa22f80 FE_RC_1612_0 ( .a(n_24059), .b(n_27655), .c(n_27845), .d(FE_OCP_RBN3120_n_27655), .o(n_27700) );
in01f80 g743063 ( .a(n_37140), .o(n_37141) );
na02f80 FE_RC_2907_0 ( .a(n_9486), .b(FE_RN_1262_0), .o(n_9527) );
in01f80 FE_OCP_RBC3838_n_19513 ( .a(FE_OCP_RBN3837_n_19513), .o(FE_OCP_RBN3838_n_19513) );
na02f80 g763143 ( .a(n_17401), .b(n_17396), .o(n_17480) );
oa22f80 FE_RC_3022_0 ( .a(n_40144), .b(n_40503), .c(n_40143), .d(n_40504), .o(n_40544) );
in01f80 drc784130 ( .a(n_45878), .o(n_45879) );
no02f80 g741205 ( .a(FE_OCP_RBN2685_n_38870), .b(n_39095), .o(n_39154) );
ms00f80 cos_out_reg_7_ ( .ck(newNet_3673), .d(n_43702), .o(cos_out_7) );
na02f80 g778923 ( .a(n_2152), .b(n_1840), .o(n_2191) );
na02f80 g766011 ( .a(n_14634), .b(n_14616), .o(n_14669) );
na02f80 FE_RC_2847_0 ( .a(n_38698), .b(n_38766), .o(FE_RN_1226_0) );
in01f80 g743747 ( .a(n_36247), .o(n_36277) );
na02f80 g777317 ( .a(FE_OCP_RBN2729_n_4219), .b(FE_OFN818_n_4575), .o(n_4739) );
no02f80 g760407 ( .a(n_20126), .b(n_20149), .o(n_20184) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_16_ ( .ck(newNet_1419), .d(n_36573), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_) );
na02f80 g746307 ( .a(n_33611), .b(n_33215), .o(n_33657) );
na02f80 g747427 ( .a(n_33746), .b(n_33745), .o(n_33747) );
no02f80 g754713 ( .a(FE_OCP_RBN2958_n_26231), .b(n_25713), .o(n_26550) );
in01f80 g750127 ( .a(n_30343), .o(n_30344) );
na02f80 g759593 ( .a(n_20641), .b(n_20548), .o(n_20687) );
ao22s80 FE_RC_3694_0 ( .a(n_10468), .b(n_10731), .c(n_10467), .d(n_10764), .o(n_10878) );
oa12f80 g758564 ( .a(n_21824), .b(n_22526), .c(n_21751), .o(n_22585) );
oa22f80 FE_RC_613_0 ( .a(n_40949), .b(n_41233), .c(n_40950), .d(n_41222), .o(n_41302) );
no02f80 g784785 ( .a(FE_OCP_RBN3084_n_31819), .b(n_30759), .o(n_47271) );
in01f80 newInst_2152 ( .a(newNet_862), .o(newNet_2152) );
in01f80 g776066 ( .a(n_5095), .o(n_5096) );
in01f80 FE_OCP_RBC1914_n_20965 ( .a(FE_OCP_RBN1913_n_20965), .o(FE_OCP_RBN1914_n_20965) );
in01f80 g752002 ( .a(n_29000), .o(n_29001) );
na02f80 g778518 ( .a(n_2569), .b(n_2500), .o(n_2594) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_8_ ( .ck(newNet_897), .d(n_27818), .o(delay_xor_ln21_unr18_stage7_stallmux_q_8_) );
in01f80 newInst_1875 ( .a(newNet_1874), .o(newNet_1875) );
no02f80 g780871 ( .a(n_420), .b(n_46055), .o(n_526) );
na02f80 FE_RC_2272_0 ( .a(FE_RN_845_0), .b(n_34132), .o(n_34174) );
no02f80 g750918 ( .a(n_28952), .b(n_28627), .o(n_28979) );
na02f80 g741207 ( .a(FE_OCP_RBN3626_n_38870), .b(n_38622), .o(n_39179) );
in01f80 newInst_2898 ( .a(newNet_2897), .o(newNet_2898) );
na02f80 g773519 ( .a(n_7435), .b(n_7289), .o(n_7436) );
in01f80 FE_OCP_RBC3462_n_7886 ( .a(n_7886), .o(FE_OCP_RBN3462_n_7886) );
in01f80 FE_OCPC3753_n_1448 ( .a(FE_OCPN3752_n_1448), .o(FE_OCPN3753_n_1448) );
ao22s80 FE_RC_3993_0 ( .a(n_34536), .b(FE_OCP_RBN2574_n_34822), .c(n_34507), .d(n_34822), .o(n_34921) );
in01f80 FE_RC_3259_0 ( .a(n_9849), .o(FE_RN_1438_0) );
in01f80 g770095 ( .a(n_10959), .o(n_10928) );
na02f80 g745230 ( .a(n_36124), .b(n_36086), .o(n_36250) );
na02f80 g778380 ( .a(n_2538), .b(n_2929), .o(n_2539) );
na02f80 g763512 ( .a(FE_OCP_RBN1207_n_16814), .b(n_15993), .o(n_16943) );
in01f80 newInst_1563 ( .a(newNet_102), .o(newNet_1563) );
no02f80 g747618 ( .a(n_45517), .b(FE_OCPN977_n_31594), .o(n_32200) );
na02f80 g769733 ( .a(n_11241), .b(n_11073), .o(n_11316) );
no02f80 g778342 ( .a(n_2537), .b(n_3023), .o(n_2557) );
in01f80 newInst_2029 ( .a(newNet_2028), .o(newNet_2029) );
no02f80 g775085 ( .a(n_6074), .b(n_5049), .o(n_6106) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_25_ ( .ck(newNet_1726), .d(n_22587), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_) );
no02f80 g739029 ( .a(n_41100), .b(n_41099), .o(n_41101) );
in01f80 g775072 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_15_), .o(n_7211) );
in01f80 newInst_3171 ( .a(newNet_3170), .o(newNet_3171) );
no02f80 g747139 ( .a(n_33953), .b(n_33602), .o(n_33998) );
ao12f80 g768269 ( .a(n_12300), .b(n_12553), .c(n_12335), .o(n_12569) );
no02f80 g766432 ( .a(n_14566), .b(n_14565), .o(n_14567) );
na02f80 g742644 ( .a(n_37420), .b(n_37419), .o(n_37446) );
no02f80 g744272 ( .a(n_44180), .b(n_34926), .o(n_36132) );
in01f80 g748260 ( .a(n_32020), .o(n_32052) );
ao12f80 g747854 ( .a(n_33132), .b(n_33131), .c(n_33130), .o(n_33684) );
in01f80 newInst_3535 ( .a(newNet_3534), .o(newNet_3535) );
in01f80 g768310 ( .a(n_12549), .o(n_12550) );
in01f80 newInst_1738 ( .a(newNet_1737), .o(newNet_1738) );
na02f80 g749519 ( .a(n_31816), .b(n_31292), .o(n_31909) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_4_ ( .ck(newNet_1074), .d(n_9832), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_) );
in01f80 newInst_2846 ( .a(newNet_2845), .o(newNet_2846) );
in01f80 g780667 ( .a(n_713), .o(n_745) );
no02f80 g737935 ( .a(n_42179), .b(n_41515), .o(n_42199) );
in01f80 newInst_1060 ( .a(newNet_1059), .o(newNet_1060) );
in01f80 FE_OCP_RBC2769_n_9892 ( .a(n_9892), .o(FE_OCP_RBN2769_n_9892) );
in01f80 g737899 ( .a(n_42215), .o(n_42227) );
ao12f80 g745433 ( .a(n_34890), .b(n_35540), .c(n_34942), .o(n_35581) );
na02f80 g777237 ( .a(n_3590), .b(n_3566), .o(n_3650) );
oa12f80 g780151 ( .a(n_1076), .b(n_1075), .c(n_1074), .o(n_1112) );
na02f80 g776633 ( .a(n_4082), .b(n_3938), .o(n_4287) );
in01f80 FE_OCPC1796_n_30546 ( .a(FE_OCPN1795_n_30546), .o(FE_OCPN1796_n_30546) );
no02f80 g766580 ( .a(n_13989), .b(n_13952), .o(n_14118) );
in01f80 FE_OCP_RBC3544_n_44575 ( .a(n_44575), .o(FE_OCP_RBN3544_n_44575) );
in01f80 g755738 ( .a(n_24405), .o(n_24406) );
oa22f80 g747359 ( .a(FE_OCP_RBN2102_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .c(n_32402), .d(n_44962), .o(n_32549) );
no02f80 g747632 ( .a(n_32055), .b(n_32301), .o(n_32346) );
ao12f80 g740439 ( .a(n_39756), .b(n_39778), .c(n_39775), .o(n_39792) );
in01f80 newInst_282 ( .a(newNet_281), .o(newNet_282) );
in01f80 FE_OCP_RBC2352_n_38534 ( .a(n_38534), .o(FE_OCP_RBN2352_n_38534) );
ao12f80 g780081 ( .a(n_1191), .b(n_1198), .c(n_814), .o(n_1199) );
no02f80 FE_RC_2266_0 ( .a(n_25134), .b(n_25167), .o(FE_RN_842_0) );
ao12f80 g750283 ( .a(n_30811), .b(n_30756), .c(n_30159), .o(n_30835) );
in01f80 FE_OCP_RBC2052_delay_xor_ln22_unr15_stage6_stallmux_q_2_ ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .o(FE_OCP_RBN2052_delay_xor_ln22_unr15_stage6_stallmux_q_2_) );
in01f80 FE_OCP_RBC3420_n_12739 ( .a(FE_OCP_RBN3418_n_12739), .o(FE_OCP_RBN3420_n_12739) );
in01f80 FE_OCP_RBC1363_n_20412 ( .a(n_20412), .o(FE_OCP_RBN1363_n_20412) );
na02f80 g779815 ( .a(delay_xor_ln23_unr3_stage2_stallmux_q), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1387) );
in01f80 g741162 ( .a(n_38833), .o(n_38860) );
no02f80 g755790 ( .a(n_24274), .b(n_23815), .o(n_24325) );
in01f80 FE_OCP_RBC3833_n_19241 ( .a(n_19241), .o(FE_OCP_RBN3833_n_19241) );
in01f80 newInst_2047 ( .a(newNet_2046), .o(newNet_2047) );
na02f80 g756999 ( .a(n_23270), .b(n_23197), .o(n_23310) );
in01f80 g770295 ( .a(n_10739), .o(n_10721) );
oa22f80 FE_RC_3389_0 ( .a(FE_RN_1162_0), .b(FE_RN_1163_0), .c(FE_RN_1164_0), .d(n_37762), .o(n_37818) );
no02f80 g757486 ( .a(n_22822), .b(n_22823), .o(n_22945) );
in01f80 newInst_478 ( .a(newNet_307), .o(newNet_478) );
na02f80 g775417 ( .a(n_5821), .b(n_47008), .o(n_5930) );
in01f80 FE_OCP_RBC1176_n_18981 ( .a(FE_OCP_RBN1175_n_18981), .o(FE_OCP_RBN1176_n_18981) );
na02f80 g745226 ( .a(n_34570), .b(n_34328), .o(n_34415) );
na02f80 g745541 ( .a(n_34532), .b(n_34560), .o(n_34561) );
in01f80 g755713 ( .a(n_24590), .o(n_24591) );
oa12f80 g772895 ( .a(n_7268), .b(n_45875), .c(n_7291), .o(n_7949) );
na02f80 g764197 ( .a(n_16824), .b(n_15927), .o(n_16852) );
in01f80 FE_OFC801_n_46285 ( .a(FE_OFN799_n_46285), .o(FE_OFN801_n_46285) );
in01f80 g760918 ( .a(n_19501), .o(n_19502) );
in01f80 FE_OCP_RBC3141_n_6477 ( .a(n_6477), .o(FE_OCP_RBN3141_n_6477) );
na02f80 g756416 ( .a(n_23737), .b(n_23739), .o(n_24162) );
in01f80 g776470 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n_4621) );
no02f80 g751151 ( .a(n_29802), .b(n_29801), .o(n_29803) );
na02f80 g775528 ( .a(n_5594), .b(n_5593), .o(n_5595) );
oa22f80 g739403 ( .a(FE_OCPN898_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .c(n_44775), .d(n_40522), .o(n_41225) );
na02f80 g777074 ( .a(n_3638), .b(n_3755), .o(n_3884) );
in01f80 fopt783292 ( .a(n_44869), .o(n_44871) );
no02f80 g740548 ( .a(n_39697), .b(n_39669), .o(n_39744) );
na02f80 g746349 ( .a(n_35043), .b(n_35042), .o(n_35044) );
in01f80 FE_OCP_RBC2456_n_13765 ( .a(n_13765), .o(FE_OCP_RBN2456_n_13765) );
in01f80 g776384 ( .a(n_4271), .o(n_4272) );
in01f80 g759022 ( .a(n_21238), .o(n_21283) );
na02f80 g750677 ( .a(n_29276), .b(n_29300), .o(n_29371) );
in01f80 g747974 ( .a(n_33552), .o(n_33114) );
in01f80 g750932 ( .a(n_29031), .o(n_29032) );
in01f80 FE_OCPC1248_n_44267 ( .a(n_44267), .o(FE_OCPN1248_n_44267) );
na02f80 FE_RC_438_0 ( .a(n_17599), .b(n_17328), .o(FE_RN_124_0) );
in01f80 newInst_2704 ( .a(newNet_2703), .o(newNet_2704) );
na02f80 g760743 ( .a(n_19595), .b(n_19656), .o(n_19720) );
na02f80 g771867 ( .a(n_9827), .b(n_9874), .o(n_10775) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_2_ ( .ck(newNet_1198), .d(n_4089), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_2_) );
in01f80 FE_RC_3627_0 ( .a(n_45010), .o(FE_RN_1589_0) );
na02f80 g781068 ( .a(cos_out_29), .b(FE_OFN1_n_43918), .o(n_292) );
no02f80 g771104 ( .a(n_9575), .b(n_9577), .o(n_9764) );
ao12f80 g751203 ( .a(n_29909), .b(n_30083), .c(n_30082), .o(n_30084) );
in01f80 g777373 ( .a(n_4261), .o(n_4262) );
in01f80 FE_OCP_RBC2703_n_9411 ( .a(n_9411), .o(FE_OCP_RBN2703_n_9411) );
ao12f80 g751887 ( .a(n_44735), .b(n_27972), .c(n_27978), .o(n_28074) );
in01f80 FE_OFC615_n_36594 ( .a(FE_OFN809_n_36594), .o(FE_OFN615_n_36594) );
na02f80 g773739 ( .a(n_7252), .b(n_7234), .o(n_7628) );
na02f80 g770277 ( .a(n_10781), .b(FE_OCP_RBN2718_n_9182), .o(n_10801) );
na02f80 g761915 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_22_), .o(n_18470) );
no02f80 g756322 ( .a(n_24587), .b(n_23957), .o(n_24609) );
in01f80 FE_OCP_RBC2433_n_14018 ( .a(FE_OCP_RBN2431_n_14018), .o(FE_OCP_RBN2433_n_14018) );
ms00f80 sin_out_reg_15_ ( .ck(newNet_75), .d(n_43813), .o(sin_out_15) );
no02f80 g774113 ( .a(n_6948), .b(n_4621), .o(n_6740) );
na02f80 g764905 ( .a(n_15546), .b(n_15548), .o(n_15727) );
in01f80 g754045 ( .a(FE_OCP_RBN2892_n_26152), .o(n_26201) );
no02f80 g737046 ( .a(n_43171), .b(n_43172), .o(n_43205) );
in01f80 newInst_497 ( .a(newNet_496), .o(newNet_497) );
no02f80 g748166 ( .a(n_47273), .b(n_30955), .o(n_31987) );
no02f80 g766193 ( .a(n_14504), .b(n_14469), .o(n_14634) );
in01f80 FE_OCP_RBC3829_n_19204 ( .a(FE_OCP_RBN3828_n_19204), .o(FE_OCP_RBN3829_n_19204) );
na03f80 FE_RC_473_0 ( .a(n_28542), .b(FE_RN_140_0), .c(n_28894), .o(n_28952) );
in01f80 g741041 ( .a(n_39057), .o(n_39058) );
oa22f80 g747889 ( .a(n_31938), .b(n_31895), .c(n_31956), .d(n_31896), .o(n_32029) );
oa12f80 g777646 ( .a(n_2569), .b(n_3320), .c(n_2499), .o(n_3400) );
na02f80 g739312 ( .a(n_45181), .b(delay_add_ln22_unr27_stage10_stallmux_q_22_), .o(n_40885) );
in01f80 newInst_587 ( .a(newNet_100), .o(newNet_587) );
ao12f80 g748783 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32416), .c(n_32157), .o(n_32494) );
no02f80 g776322 ( .a(n_4766), .b(n_4765), .o(n_4767) );
na02f80 g776558 ( .a(n_4273), .b(n_4387), .o(n_4487) );
no02f80 g750999 ( .a(n_30124), .b(n_30161), .o(n_30162) );
in01f80 FE_RC_4089_0 ( .a(n_15479), .o(FE_RN_1788_0) );
no02f80 g737700 ( .a(n_42198), .b(n_42211), .o(n_42222) );
oa12f80 g772943 ( .a(n_7886), .b(n_8151), .c(n_8150), .o(n_8153) );
na02f80 g764113 ( .a(n_16588), .b(FE_OCP_RBN2697_n_14814), .o(n_16641) );
in01f80 g749829 ( .a(n_31528), .o(n_31529) );
oa12f80 g777201 ( .a(n_3483), .b(n_3533), .c(n_3532), .o(n_3560) );
in01f80 newInst_2457 ( .a(newNet_526), .o(newNet_2457) );
na02f80 g773912 ( .a(n_7002), .b(n_5393), .o(n_7082) );
na02f80 g753129 ( .a(n_27298), .b(n_27297), .o(n_27299) );
in01f80 FE_OCP_RBC2385_n_8342 ( .a(FE_OCP_RBN2383_n_8342), .o(FE_OCP_RBN2385_n_8342) );
na02f80 g736924 ( .a(n_43015), .b(n_43014), .o(n_43043) );
na02f80 g760838 ( .a(FE_OCP_RBN3495_n_19390), .b(FE_OCP_RBN1701_n_19353), .o(n_19472) );
in01f80 g736676 ( .a(n_43413), .o(n_43368) );
in01f80 g773420 ( .a(n_8840), .o(n_7549) );
no02f80 g743883 ( .a(n_35985), .b(n_35820), .o(n_36012) );
no02f80 g755579 ( .a(n_24534), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24536) );
in01f80 g772713 ( .a(n_8271), .o(n_8272) );
no02f80 g759916 ( .a(n_21051), .b(n_21249), .o(n_21378) );
in01f80 g751962 ( .a(n_29006), .o(n_28986) );
no02f80 FE_RC_1862_0 ( .a(FE_OCP_RBN2354_n_13858), .b(n_14032), .o(FE_RN_572_0) );
ao12f80 g772840 ( .a(n_7977), .b(n_7976), .c(n_7975), .o(n_9172) );
na02f80 g745743 ( .a(n_34116), .b(n_34187), .o(n_34466) );
in01f80 g763721 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .o(n_16891) );
in01f80 g742691 ( .a(n_37411), .o(n_38268) );
no02f80 g772325 ( .a(n_8512), .b(n_8575), .o(n_8631) );
oa12f80 g758324 ( .a(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n_22812) );
in01f80 g738365 ( .a(n_41773), .o(n_41774) );
ao12f80 g779453 ( .a(n_1998), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .o(n_2001) );
no02f80 g763058 ( .a(n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .o(n_17641) );
in01f80 g772650 ( .a(n_8284), .o(n_8285) );
in01f80 g757725 ( .a(n_23807), .o(n_24111) );
no02f80 g774478 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .o(n_6741) );
in01f80 g767844 ( .a(n_12986), .o(n_13043) );
na02f80 g758589 ( .a(n_22034), .b(n_21961), .o(n_22035) );
in01f80 g746897 ( .a(n_33259), .o(n_33851) );
in01f80 newInst_3507 ( .a(newNet_3506), .o(newNet_3507) );
na02f80 g756820 ( .a(n_24046), .b(n_24091), .o(n_24739) );
in01f80 g760903 ( .a(FE_OCP_RBN3495_n_19390), .o(n_19461) );
na02f80 g757903 ( .a(n_22314), .b(n_22234), .o(n_22473) );
in01f80 g776193 ( .a(n_4956), .o(n_5007) );
in01f80 FE_OCP_DRV_C3744_FE_OFN737_n_22641 ( .a(FE_OFN737_n_22641), .o(FE_OCP_DRV_N3744_FE_OFN737_n_22641) );
in01f80 FE_RC_598_0 ( .a(n_25813), .o(FE_RN_187_0) );
oa22f80 g779847 ( .a(n_44652), .b(n_1190), .c(n_44623), .d(n_1183), .o(n_1302) );
ao12f80 g752212 ( .a(n_28027), .b(n_28539), .c(n_27950), .o(n_28617) );
na02f80 g750611 ( .a(n_29380), .b(n_46960), .o(n_29382) );
no02f80 g746467 ( .a(n_33453), .b(n_33452), .o(n_33454) );
na02f80 g755187 ( .a(n_25640), .b(n_25218), .o(n_25715) );
in01f80 FE_OCP_RBC3004_n_10930 ( .a(n_10930), .o(FE_OCP_RBN3004_n_10930) );
in01f80 g764742 ( .a(n_16450), .o(n_16415) );
no02f80 g745624 ( .a(n_34286), .b(n_33594), .o(n_34484) );
no02f80 g753717 ( .a(n_27135), .b(n_26772), .o(n_27203) );
in01f80 newInst_3622 ( .a(newNet_2649), .o(newNet_3622) );
no02f80 g770944 ( .a(n_9756), .b(FE_OCP_RBN3597_FE_OCPN1243_n_44460), .o(n_9759) );
in01f80 g756378 ( .a(n_23859), .o(n_23948) );
no02f80 g736772 ( .a(n_43361), .b(n_43270), .o(n_43318) );
no02f80 g751408 ( .a(n_29224), .b(n_28959), .o(n_29363) );
ao12f80 g741455 ( .a(n_38772), .b(n_38807), .c(n_38790), .o(n_38843) );
in01f80 newInst_3207 ( .a(newNet_3206), .o(newNet_3207) );
in01f80 g755744 ( .a(n_25309), .o(n_25310) );
no02f80 g745562 ( .a(n_34565), .b(n_34531), .o(n_34622) );
in01f80 FE_OCPC1532_n_21790 ( .a(FE_OCPN1531_n_21790), .o(FE_OCPN1532_n_21790) );
na02f80 g741899 ( .a(n_38242), .b(n_38010), .o(n_38243) );
na02f80 g771396 ( .a(FE_OCP_RBN3524_n_8242), .b(n_9088), .o(n_9213) );
na02f80 g740754 ( .a(n_39353), .b(n_39362), .o(n_39412) );
in01f80 g772971 ( .a(n_7749), .o(n_7750) );
no02f80 g753560 ( .a(n_26721), .b(n_25100), .o(n_26799) );
oa12f80 g741080 ( .a(n_39009), .b(FE_OCP_RBN3628_n_38870), .c(n_38919), .o(n_39502) );
ao22s80 FE_RC_290_0 ( .a(n_20704), .b(n_21178), .c(n_20703), .d(n_21177), .o(n_21346) );
no02f80 g740746 ( .a(n_39443), .b(n_39411), .o(n_39910) );
na02f80 g780243 ( .a(n_960), .b(n_1155), .o(n_961) );
in01f80 g762830 ( .a(n_18123), .o(n_18156) );
in01f80 g744278 ( .a(n_35687), .o(n_35820) );
in01f80 newInst_2279 ( .a(newNet_2278), .o(newNet_2279) );
in01f80 g753177 ( .a(n_27421), .o(n_27422) );
in01f80 FE_RC_1558_0 ( .a(n_2621), .o(FE_RN_442_0) );
in01f80 g751454 ( .a(n_28628), .o(n_28629) );
na02f80 g746550 ( .a(n_34889), .b(n_34666), .o(n_35159) );
oa12f80 g784661 ( .a(n_7868), .b(n_45875), .c(n_7318), .o(n_46991) );
na02f80 g762127 ( .a(n_18172), .b(n_18202), .o(n_18218) );
na02f80 g745464 ( .a(n_34369), .b(n_34510), .o(n_34568) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_22_ ( .ck(newNet_165), .d(n_46349), .o(delay_xor_ln22_unr9_stage4_stallmux_q_22_) );
no02f80 g776396 ( .a(n_4161), .b(n_4185), .o(n_4376) );
no02f80 g769763 ( .a(n_11087), .b(n_44463), .o(n_11121) );
ao12f80 g781225 ( .a(n_7), .b(n_116), .c(n_40), .o(n_115) );
in01f80 g773997 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .o(n_6809) );
in01f80 newInst_1373 ( .a(newNet_748), .o(newNet_1373) );
na02f80 g765980 ( .a(n_14915), .b(n_14896), .o(n_14897) );
in01f80 g743132 ( .a(n_37036), .o(n_37037) );
na02f80 g779122 ( .a(n_1950), .b(n_1949), .o(n_1951) );
in01f80 newInst_2961 ( .a(newNet_2960), .o(newNet_2961) );
oa22f80 g753314 ( .a(n_27611), .b(n_26869), .c(n_27612), .d(n_26870), .o(n_27656) );
no02f80 g743001 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_22_), .o(n_37070) );
in01f80 newInst_2696 ( .a(newNet_1652), .o(newNet_2696) );
in01f80 newInst_1361 ( .a(newNet_1360), .o(newNet_1361) );
ao12f80 g767405 ( .a(n_13358), .b(n_13448), .c(n_13403), .o(n_13548) );
na02f80 g737191 ( .a(n_42987), .b(n_42995), .o(n_43388) );
na02f80 g748939 ( .a(n_31013), .b(FE_OCP_DRV_N1588_n_31012), .o(n_31035) );
no02f80 g759357 ( .a(n_21121), .b(n_45032), .o(n_21214) );
na02f80 g740624 ( .a(n_39628), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39640) );
in01f80 g752302 ( .a(n_28479), .o(n_28480) );
na02f80 g740243 ( .a(n_39915), .b(n_39914), .o(n_39916) );
in01f80 g744285 ( .a(n_35776), .o(n_35815) );
no02f80 g753552 ( .a(n_26729), .b(n_26671), .o(n_26785) );
in01f80 g760257 ( .a(n_20428), .o(n_20429) );
no02f80 g757666 ( .a(n_22668), .b(n_22413), .o(n_22745) );
na02f80 g758754 ( .a(n_21616), .b(n_21708), .o(n_21736) );
na02f80 g753395 ( .a(n_26990), .b(n_27026), .o(n_27042) );
oa12f80 g745552 ( .a(n_34317), .b(n_34286), .c(n_34343), .o(n_34823) );
na02f80 g780934 ( .a(n_420), .b(n_242), .o(n_446) );
no02f80 g749575 ( .a(n_30377), .b(n_30376), .o(n_30378) );
na02f80 g765263 ( .a(n_15517), .b(n_15571), .o(n_15671) );
in01f80 g750424 ( .a(n_29612), .o(n_29613) );
no02f80 g757762 ( .a(n_22483), .b(n_44287), .o(n_22538) );
in01f80 g765737 ( .a(n_15514), .o(n_15565) );
na02f80 g764857 ( .a(n_15619), .b(n_47333), .o(n_15755) );
oa12f80 g736634 ( .a(n_43242), .b(n_43564), .c(n_43298), .o(n_43623) );
in01f80 g754798 ( .a(n_26163), .o(n_26160) );
in01f80 FE_RC_3187_0 ( .a(n_17847), .o(FE_RN_1415_0) );
na02f80 g770716 ( .a(n_10258), .b(n_10259), .o(n_10410) );
na02f80 g761662 ( .a(n_18759), .b(n_18718), .o(n_18719) );
oa12f80 g747768 ( .a(n_33738), .b(n_33571), .c(n_33720), .o(n_34230) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_20_ ( .ck(newNet_638), .d(n_46345), .o(delay_xor_ln21_unr9_stage4_stallmux_q_20_) );
in01f80 g739676 ( .a(n_40592), .o(n_40583) );
in01f80 g771842 ( .a(n_10156), .o(n_10157) );
no02f80 g775399 ( .a(n_5793), .b(n_5587), .o(n_5838) );
na02f80 g743706 ( .a(n_36346), .b(n_35988), .o(n_36373) );
no02f80 g760775 ( .a(n_19559), .b(FE_OCP_RBN1840_n_19528), .o(n_19629) );
in01f80 g737653 ( .a(n_42797), .o(n_42798) );
in01f80 g764611 ( .a(n_16036), .o(n_16037) );
no02f80 g770829 ( .a(n_9808), .b(n_9749), .o(n_9867) );
no02f80 g765327 ( .a(n_15135), .b(FE_OCP_RBN2433_n_14018), .o(n_15300) );
no02f80 FE_RC_1424_0 ( .a(n_22304), .b(n_22476), .o(FE_RN_415_0) );
na02f80 g738747 ( .a(n_41375), .b(n_41371), .o(n_41422) );
na02f80 FE_RC_4223_0 ( .a(n_29954), .b(FE_RN_1851_0), .o(FE_RN_1852_0) );
in01f80 g772476 ( .a(n_8380), .o(n_8379) );
no02f80 g770511 ( .a(n_10529), .b(FE_OCP_RBN2539_n_8781), .o(n_10556) );
oa22f80 FE_RC_3828_0 ( .a(n_24059), .b(n_27793), .c(n_27796), .d(n_27743), .o(n_27815) );
in01f80 newInst_1103 ( .a(newNet_1102), .o(newNet_1103) );
no02f80 g755870 ( .a(n_25195), .b(n_25216), .o(n_25196) );
no02f80 g740091 ( .a(n_40066), .b(n_40032), .o(n_40067) );
in01f80 g762682 ( .a(n_17924), .o(n_17925) );
in01f80 g772735 ( .a(n_8237), .o(n_8238) );
no02f80 g762111 ( .a(FE_OCP_RBN2205_n_18242), .b(n_17813), .o(n_18462) );
in01f80 FE_OCP_RBC2588_n_9492 ( .a(n_9492), .o(FE_OCP_RBN2588_n_9492) );
oa22f80 g774840 ( .a(n_6209), .b(n_5380), .c(n_6210), .d(n_5381), .o(n_6286) );
na02f80 g741199 ( .a(FE_OCP_RBN2636_n_38806), .b(n_38917), .o(n_39006) );
in01f80 newInst_3400 ( .a(newNet_2542), .o(newNet_3400) );
ao12f80 g772460 ( .a(n_8398), .b(n_8462), .c(FE_OCP_RBN3466_n_7886), .o(n_8515) );
in01f80 newInst_2243 ( .a(newNet_2242), .o(newNet_2243) );
na02f80 g763253 ( .a(n_17130), .b(FE_OCPN869_n_16086), .o(n_17196) );
oa12f80 g760983 ( .a(n_17881), .b(n_19278), .c(n_19273), .o(n_19330) );
in01f80 g779135 ( .a(n_2702), .o(n_1978) );
in01f80 g767614 ( .a(n_12805), .o(n_12830) );
in01f80 g736901 ( .a(n_43579), .o(n_43580) );
no02f80 g737903 ( .a(n_42189), .b(n_42188), .o(n_42220) );
in01f80 newInst_595 ( .a(newNet_594), .o(newNet_595) );
in01f80 g770371 ( .a(n_10713), .o(n_10714) );
na02f80 g772875 ( .a(n_8153), .b(n_8143), .o(n_8200) );
na02f80 g770505 ( .a(n_10292), .b(FE_OCP_RBN3601_FE_OCPN1243_n_44460), .o(n_10367) );
in01f80 g757016 ( .a(n_24234), .o(n_24235) );
no02f80 g743097 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_), .o(n_37426) );
in01f80 g767335 ( .a(n_13568), .o(n_13609) );
na02f80 g746815 ( .a(n_33247), .b(n_33289), .o(n_33303) );
ao12f80 g754273 ( .a(n_26343), .b(n_26646), .c(n_26690), .o(n_26744) );
in01f80 g779120 ( .a(n_2024), .o(n_2042) );
no02f80 g771537 ( .a(n_9337), .b(n_9338), .o(n_9398) );
no02f80 g749587 ( .a(n_30448), .b(n_30447), .o(n_30449) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_4_ ( .ck(newNet_3373), .d(n_26668), .o(delay_add_ln22_unr17_stage7_stallmux_q_4_) );
na02f80 g766370 ( .a(n_14096), .b(n_13916), .o(n_14160) );
na02f80 g764881 ( .a(n_15394), .b(n_15267), .o(n_15439) );
no02f80 g746398 ( .a(n_33388), .b(n_32995), .o(n_33411) );
in01f80 FE_OCP_RBC1350_n_19148 ( .a(n_19148), .o(FE_OCP_RBN1350_n_19148) );
in01f80 FE_RC_3508_0 ( .a(FE_RN_1515_0), .o(FE_RN_1513_0) );
oa12f80 g743689 ( .a(n_37383), .b(n_37382), .c(n_37381), .o(n_37541) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_26_ ( .ck(newNet_2458), .d(n_32512), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_26_) );
no02f80 g741187 ( .a(FE_OCP_RBN2637_n_38806), .b(n_38513), .o(n_38987) );
no02f80 FE_RC_498_0 ( .a(FE_RN_149_0), .b(n_28231), .o(n_28306) );
in01f80 fopt782889 ( .a(n_22875), .o(n_44329) );
in01f80 newInst_138 ( .a(newNet_137), .o(newNet_138) );
in01f80 g757921 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_13_), .o(n_22203) );
in01f80 g757073 ( .a(n_24088), .o(n_23641) );
in01f80 newInst_1920 ( .a(newNet_1919), .o(newNet_1920) );
in01f80 g779609 ( .a(n_1802), .o(n_1803) );
in01f80 g754185 ( .a(n_26114), .o(n_26107) );
oa22f80 FE_RC_2986_0 ( .a(n_23486), .b(n_26464), .c(n_23590), .d(n_26492), .o(n_26583) );
in01f80 newInst_2241 ( .a(newNet_2240), .o(newNet_2241) );
na02f80 g777186 ( .a(n_3757), .b(n_3726), .o(n_3903) );
na02f80 g764842 ( .a(n_15556), .b(n_45501), .o(n_15734) );
oa22f80 FE_RC_39_0 ( .a(FE_OFN84_n_46137), .b(n_6700), .c(FE_OFN806_n_46196), .d(n_6739), .o(n_46191) );
no02f80 g738084 ( .a(n_42082), .b(n_41599), .o(n_42145) );
no02f80 g765490 ( .a(n_15599), .b(n_15869), .o(n_15920) );
in01f80 g752317 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_27834) );
na02f80 g776301 ( .a(n_4472), .b(n_3029), .o(n_4666) );
na02f80 g768394 ( .a(n_12476), .b(n_12507), .o(n_12526) );
in01f80 FE_RC_2657_0 ( .a(n_8107), .o(FE_RN_1110_0) );
na02f80 g736892 ( .a(n_43488), .b(n_43186), .o(n_43589) );
oa12f80 g780196 ( .a(n_1030), .b(n_1069), .c(n_1180), .o(n_1137) );
na02f80 g741613 ( .a(n_38589), .b(n_38584), .o(n_38654) );
no02f80 g742771 ( .a(n_37514), .b(n_36957), .o(n_37561) );
na02f80 g759281 ( .a(n_20803), .b(n_20579), .o(n_20866) );
in01f80 g758889 ( .a(n_21501), .o(n_21502) );
in01f80 g776299 ( .a(n_4535), .o(n_4583) );
na02f80 g771088 ( .a(n_9924), .b(n_9923), .o(n_9925) );
no02f80 g758804 ( .a(n_21504), .b(n_19962), .o(n_21660) );
na02f80 g738671 ( .a(n_41525), .b(n_41563), .o(n_41608) );
na02f80 g740158 ( .a(FE_OCP_RBN3722_n_39913), .b(n_40183), .o(n_40292) );
na02f80 g780381 ( .a(n_907), .b(n_805), .o(n_942) );
no02f80 g777193 ( .a(n_5548), .b(n_4773), .o(n_5517) );
ao12f80 g775597 ( .a(n_5548), .b(n_5552), .c(n_4702), .o(n_5594) );
in01f80 newInst_2927 ( .a(newNet_2926), .o(newNet_2927) );
no02f80 g753839 ( .a(n_26268), .b(FE_OCPN1488_n_23447), .o(n_26336) );
na02f80 g754887 ( .a(n_25485), .b(n_25452), .o(n_25562) );
no02f80 g769213 ( .a(n_11738), .b(n_11727), .o(n_12139) );
no02f80 g769060 ( .a(FE_OCP_RBN1094_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(n_11919) );
in01f80 newInst_159 ( .a(newNet_14), .o(newNet_159) );
ao12f80 g768994 ( .a(n_11756), .b(FE_OCP_RBN2119_n_45224), .c(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .o(n_11877) );
na02f80 g742005 ( .a(n_38181), .b(n_38216), .o(n_38239) );
in01f80 g743245 ( .a(n_36801), .o(n_36832) );
in01f80 g780331 ( .a(n_957), .o(n_1022) );
na02f80 g779282 ( .a(n_1696), .b(n_1657), .o(n_1795) );
in01f80 g754742 ( .a(n_26415), .o(n_26416) );
oa12f80 g753541 ( .a(n_26703), .b(n_26702), .c(n_26701), .o(n_26761) );
oa22f80 FE_RC_867_0 ( .a(n_27490), .b(n_27701), .c(n_27491), .d(n_27702), .o(n_27799) );
na02f80 g776712 ( .a(n_4016), .b(n_3845), .o(n_4130) );
no02f80 FE_RC_2577_0 ( .a(FE_RN_1059_0), .b(FE_RN_1060_0), .o(FE_RN_1061_0) );
in01f80 g768648 ( .a(n_12146), .o(n_12233) );
na02f80 g763813 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .o(n_17428) );
in01f80 g756785 ( .a(n_23456), .o(n_23514) );
na02f80 g765331 ( .a(FE_OCP_RBN3621_n_15135), .b(FE_OCP_RBN2436_n_14072), .o(n_15335) );
na02f80 g773133 ( .a(n_7617), .b(n_7690), .o(n_7710) );
in01f80 fopt783211 ( .a(n_32316), .o(n_44764) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_10_ ( .ck(newNet_597), .d(n_17585), .o(delay_xor_ln22_unr12_stage5_stallmux_q_10_) );
no02f80 g762416 ( .a(n_18421), .b(n_18416), .o(n_18443) );
na02f80 FE_RC_3172_0 ( .a(FE_RN_1405_0), .b(n_22536), .o(n_46965) );
no02f80 g759236 ( .a(n_21125), .b(n_21045), .o(n_21184) );
na02f80 g736898 ( .a(n_43203), .b(n_43484), .o(n_43583) );
ao22s80 FE_RC_1268_0 ( .a(n_38212), .b(n_38577), .c(n_38211), .d(n_38578), .o(n_38622) );
na02f80 g781159 ( .a(n_189), .b(n_188), .o(n_190) );
in01f80 g770474 ( .a(n_10440), .o(n_10441) );
no02f80 g737349 ( .a(n_42821), .b(n_42763), .o(n_42832) );
in01f80 FE_OCP_RBC3458_n_33872 ( .a(FE_OCP_RBN3457_n_33872), .o(FE_OCP_RBN3458_n_33872) );
na03f80 g749721 ( .a(n_31394), .b(n_31314), .c(n_31393), .o(n_31456) );
in01f80 FE_RC_982_0 ( .a(n_27395), .o(FE_RN_282_0) );
in01f80 FE_OCP_RBC3847_FE_RN_1548_0 ( .a(FE_RN_1548_0), .o(FE_OCP_RBN3847_FE_RN_1548_0) );
ao12f80 g782666 ( .a(n_485), .b(n_457), .c(n_465), .o(n_44060) );
na02f80 g779250 ( .a(n_1834), .b(n_1833), .o(n_1981) );
na02f80 g764332 ( .a(n_16289), .b(n_16363), .o(n_16493) );
in01f80 g757696 ( .a(n_23221), .o(n_23244) );
oa12f80 g749174 ( .a(n_31513), .b(n_32115), .c(n_31432), .o(n_32227) );
ao12f80 g768720 ( .a(n_11617), .b(n_12024), .c(n_11752), .o(n_12025) );
in01f80 g753200 ( .a(n_27145), .o(n_27231) );
oa12f80 g738437 ( .a(n_41676), .b(FE_OCPN952_n_41540), .c(n_41634), .o(n_41906) );
na02f80 g750856 ( .a(FE_OCP_RBN1324_n_29056), .b(FE_OFN811_n_29140), .o(n_29188) );
in01f80 g752618 ( .a(n_27604), .o(n_27605) );
in01f80 g773853 ( .a(n_7108), .o(n_7109) );
no02f80 g752763 ( .a(n_27402), .b(n_27464), .o(n_27511) );
na02f80 g737450 ( .a(n_42670), .b(n_42386), .o(n_42716) );
na02f80 g738276 ( .a(n_41801), .b(n_41646), .o(n_41846) );
in01f80 g742427 ( .a(n_37719), .o(n_37734) );
ms00f80 cos_out_reg_6_ ( .ck(newNet_3678), .d(n_43688), .o(cos_out_6) );
no02f80 g770118 ( .a(n_10704), .b(n_10729), .o(n_10833) );
ao22s80 FE_RC_3240_0 ( .a(FE_OCP_RBN2792_n_9910), .b(n_10060), .c(n_10019), .d(n_9910), .o(n_10225) );
in01f80 g742510 ( .a(FE_OCP_RBN3397_n_37624), .o(n_37653) );
in01f80 g761898 ( .a(n_18544), .o(n_18545) );
no02f80 g743607 ( .a(n_36502), .b(n_36485), .o(n_36543) );
in01f80 newInst_3087 ( .a(newNet_3086), .o(newNet_3087) );
no02f80 g777679 ( .a(n_3377), .b(n_3371), .o(n_4905) );
na02f80 g741108 ( .a(n_39021), .b(n_39044), .o(n_39076) );
in01f80 g750441 ( .a(n_29634), .o(n_29591) );
oa22f80 FE_RC_3739_0 ( .a(n_21636), .b(n_21492), .c(n_21491), .d(n_21637), .o(n_21789) );
na02f80 g765971 ( .a(n_14712), .b(FE_OCP_RBN2503_n_13896), .o(n_14748) );
na02f80 g750333 ( .a(n_29716), .b(FE_OCPN1768_n_29715), .o(n_29764) );
in01f80 newInst_1320 ( .a(newNet_723), .o(newNet_1320) );
na02f80 g739410 ( .a(FE_OCPN898_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n_41022) );
na02f80 g771900 ( .a(n_8798), .b(n_8508), .o(n_8859) );
ao12f80 g760518 ( .a(n_19842), .b(n_19924), .c(n_19786), .o(n_19972) );
na02f80 g742307 ( .a(n_37815), .b(n_37778), .o(n_37835) );
in01f80 g772709 ( .a(n_8163), .o(n_8164) );
no02f80 g757045 ( .a(n_23803), .b(n_23801), .o(n_23900) );
in01f80 newInst_3637 ( .a(newNet_3636), .o(newNet_3637) );
na02f80 g773548 ( .a(n_7405), .b(n_7404), .o(n_7406) );
in01f80 FE_RC_2488_0 ( .a(n_23680), .o(FE_RN_1006_0) );
no02f80 g756468 ( .a(n_23585), .b(n_23664), .o(n_23689) );
na02f80 g758621 ( .a(n_22489), .b(n_21796), .o(n_22526) );
in01f80 g756405 ( .a(n_23826), .o(n_23777) );
na02f80 g759781 ( .a(n_21598), .b(n_21622), .o(n_21627) );
na02f80 g739368 ( .a(n_41013), .b(n_40982), .o(n_41036) );
in01f80 newInst_517 ( .a(newNet_273), .o(newNet_517) );
in01f80 FE_OCPC1482_n_22207 ( .a(FE_OCPN1481_n_22207), .o(FE_OCPN1482_n_22207) );
in01f80 g776390 ( .a(n_4323), .o(n_4363) );
no02f80 FE_RC_2829_0 ( .a(n_29586), .b(FE_RN_1215_0), .o(n_29663) );
no02f80 FE_RC_4069_0 ( .a(FE_RN_1771_0), .b(n_26802), .o(n_26822) );
ao12f80 g771154 ( .a(n_9385), .b(n_9884), .c(n_9475), .o(n_10001) );
in01f80 g766548 ( .a(n_14000), .o(n_13958) );
in01f80 g756718 ( .a(n_23626), .o(n_23594) );
ao12f80 g754586 ( .a(n_26860), .b(n_26856), .c(n_26680), .o(n_26894) );
no02f80 g750305 ( .a(n_29766), .b(n_29765), .o(n_29775) );
no03m80 FE_RC_1083_0 ( .a(n_41084), .b(n_41083), .c(n_40806), .o(n_41110) );
ao12f80 g756061 ( .a(n_24998), .b(n_25085), .c(n_25000), .o(n_24996) );
in01f80 FE_OCP_RBC2261_n_33691 ( .a(n_33691), .o(FE_OCP_RBN2261_n_33691) );
na02f80 g744014 ( .a(n_36295), .b(n_36265), .o(n_36359) );
no02f80 g770052 ( .a(n_10890), .b(n_10834), .o(n_10954) );
oa12f80 g763024 ( .a(n_17082), .b(n_17403), .c(n_17515), .o(n_17557) );
in01f80 g776702 ( .a(n_4368), .o(n_4369) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_6_ ( .ck(newNet_691), .d(n_46170), .o(delay_xor_ln21_unr6_stage3_stallmux_q_6_) );
no02f80 g772578 ( .a(n_8336), .b(n_7886), .o(n_8455) );
no02f80 FE_RC_2569_0 ( .a(n_12619), .b(n_13270), .o(FE_RN_1055_0) );
oa12f80 g745768 ( .a(n_34130), .b(n_44112), .c(n_34118), .o(n_34519) );
no02f80 g742773 ( .a(n_37346), .b(n_37345), .o(n_37347) );
in01f80 g754164 ( .a(n_26049), .o(n_26050) );
na02f80 g746430 ( .a(n_33351), .b(n_33350), .o(n_33352) );
oa22f80 g757638 ( .a(n_23244), .b(n_22762), .c(n_23220), .d(n_22761), .o(n_23746) );
na02f80 g778326 ( .a(n_2524), .b(n_2066), .o(n_2615) );
na02f80 g776943 ( .a(n_4008), .b(FE_OFN78_n_4117), .o(n_4400) );
in01f80 newInst_3126 ( .a(newNet_3125), .o(newNet_3126) );
in01f80 FE_OCP_DRV_C3155_n_15342 ( .a(n_15342), .o(FE_OCP_DRV_N3155_n_15342) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_8_ ( .ck(newNet_1941), .d(n_10524), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_) );
no02f80 FE_RC_3855_0 ( .a(FE_RN_1682_0), .b(n_20160), .o(n_20161) );
in01f80 g739762 ( .a(n_40511), .o(n_40538) );
oa12f80 g749636 ( .a(n_29965), .b(n_30283), .c(n_29899), .o(n_30458) );
no02f80 g755537 ( .a(n_24748), .b(n_24747), .o(n_24776) );
na02f80 g754281 ( .a(n_25856), .b(n_25879), .o(n_25931) );
in01f80 g738560 ( .a(n_41504), .o(n_41505) );
na02f80 g755902 ( .a(n_24232), .b(n_24269), .o(n_24320) );
oa22f80 FE_RC_1019_0 ( .a(n_20003), .b(n_19813), .c(n_19838), .d(n_20028), .o(n_20095) );
no02f80 g763907 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_), .o(n_17362) );
na02f80 g757850 ( .a(n_22279), .b(n_22084), .o(n_22356) );
na02f80 g751195 ( .a(n_29837), .b(n_29938), .o(n_29974) );
na02f80 g781301 ( .a(beta_29), .b(beta_31), .o(n_128) );
na02f80 g738189 ( .a(n_41989), .b(n_41662), .o(n_42006) );
in01f80 g759010 ( .a(n_21632), .o(n_21633) );
oa22f80 FE_RC_959_0 ( .a(n_28336), .b(n_32466), .c(n_32566), .d(n_32517), .o(n_32565) );
na02f80 g758579 ( .a(n_21875), .b(FE_OCPN856_n_20367), .o(n_21954) );
in01f80 g773559 ( .a(n_7411), .o(n_7412) );
na02f80 g764959 ( .a(n_15472), .b(n_14215), .o(n_15473) );
in01f80 g753694 ( .a(n_26583), .o(n_26664) );
ao22s80 FE_RC_1385_0 ( .a(n_26143), .b(n_25695), .c(n_25696), .d(n_26142), .o(n_26276) );
na02f80 g780488 ( .a(n_869), .b(n_868), .o(n_870) );
in01f80 newInst_3621 ( .a(newNet_3620), .o(newNet_3621) );
na02f80 g774739 ( .a(n_6239), .b(n_6169), .o(n_6277) );
in01f80 newInst_980 ( .a(newNet_979), .o(newNet_980) );
in01f80 g762381 ( .a(n_18665), .o(n_18571) );
no02f80 FE_RC_180_0 ( .a(FE_RN_58_0), .b(FE_RN_57_0), .o(FE_RN_59_0) );
na02f80 g738918 ( .a(n_41283), .b(n_41282), .o(n_41284) );
in01f80 g774039 ( .a(n_6802), .o(n_6752) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_31_ ( .ck(newNet_2623), .d(n_22835), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_) );
no02f80 g770239 ( .a(n_10618), .b(n_10306), .o(n_10648) );
oa12f80 g736440 ( .a(n_43480), .b(n_43716), .c(n_43225), .o(n_43781) );
na02f80 g754362 ( .a(n_25759), .b(n_25446), .o(n_25821) );
no02f80 g778089 ( .a(n_3003), .b(n_2981), .o(n_3076) );
no03m80 FE_RC_4272_0 ( .a(n_18870), .b(n_18513), .c(n_18871), .o(n_18901) );
in01f80 g737594 ( .a(n_42817), .o(n_42818) );
na02f80 g768055 ( .a(FE_OCPN860_n_12880), .b(n_12871), .o(n_13078) );
na02f80 g779060 ( .a(n_2086), .b(delay_add_ln22_unr2_stage2_stallmux_q_15_), .o(n_2123) );
in01f80 g762132 ( .a(n_18259), .o(n_18260) );
oa12f80 g756200 ( .a(n_23634), .b(n_24072), .c(n_23638), .o(n_24084) );
in01f80 FE_OCP_RBC2727_n_4219 ( .a(FE_OCP_RBN2724_n_4219), .o(FE_OCP_RBN2727_n_4219) );
no02f80 g740185 ( .a(FE_OCP_RBN3052_n_39913), .b(n_39531), .o(n_40112) );
in01f80 g776419 ( .a(n_4403), .o(n_4699) );
oa22f80 FE_RC_1420_0 ( .a(FE_OFN806_n_46196), .b(n_6719), .c(FE_OFN84_n_46137), .d(n_6701), .o(n_46194) );
in01f80 newInst_2507 ( .a(newNet_544), .o(newNet_2507) );
in01f80 newInst_684 ( .a(newNet_683), .o(newNet_684) );
in01f80 FE_OCP_RBC2864_n_39523 ( .a(n_39523), .o(FE_OCP_RBN2864_n_39523) );
na02f80 g748226 ( .a(n_31765), .b(n_30284), .o(n_31805) );
na02f80 g744888 ( .a(n_35000), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35056) );
na02f80 g777914 ( .a(n_3114), .b(n_2967), .o(n_3115) );
in01f80 g766626 ( .a(FE_OCP_RBN2356_n_13858), .o(n_13950) );
in01f80 g754855 ( .a(n_25695), .o(n_25696) );
in01f80 g771434 ( .a(n_9112), .o(n_9047) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_4_ ( .ck(newNet_3282), .d(n_31182), .o(delay_add_ln22_unr20_stage8_stallmux_q_4_) );
no03m80 FE_RC_148_0 ( .a(n_18051), .b(n_18052), .c(n_17971), .o(n_18047) );
na02f80 g750437 ( .a(n_29564), .b(n_29583), .o(n_29609) );
na02f80 g763378 ( .a(FE_OCP_RBN3725_n_16975), .b(FE_OCP_RBN2850_n_46982), .o(n_17223) );
na03f80 g746377 ( .a(n_33388), .b(n_33386), .c(n_33017), .o(n_33412) );
oa12f80 g774269 ( .a(n_6395), .b(n_6514), .c(n_6279), .o(n_6581) );
na02f80 g747093 ( .a(n_32889), .b(n_32683), .o(n_32908) );
na02f80 g762402 ( .a(n_18421), .b(n_18417), .o(n_18701) );
no02f80 g755173 ( .a(n_24945), .b(n_23627), .o(n_25024) );
na02f80 g750756 ( .a(n_29218), .b(n_28727), .o(n_29232) );
ao12f80 g764212 ( .a(n_15834), .b(n_16741), .c(n_15778), .o(n_16818) );
na02f80 FE_RC_3565_0 ( .a(n_18949), .b(n_20164), .o(FE_RN_1548_0) );
in01f80 g743151 ( .a(n_36947), .o(n_36948) );
in01f80 newInst_624 ( .a(newNet_623), .o(newNet_624) );
in01f80 g778472 ( .a(n_2656), .o(n_2657) );
in01f80 FE_OCP_RBC3657_n_15314 ( .a(n_15314), .o(FE_OCP_RBN3657_n_15314) );
in01f80 g776480 ( .a(n_4366), .o(n_4405) );
na02f80 g745707 ( .a(n_34223), .b(FE_OCPN3763_n_34222), .o(n_34245) );
no02f80 g765784 ( .a(n_14979), .b(n_14758), .o(n_14981) );
no02f80 g758151 ( .a(n_22667), .b(n_22331), .o(n_22376) );
in01f80 g777582 ( .a(n_3698), .o(n_3700) );
no02f80 g743022 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_30_), .o(n_36955) );
in01f80 g777404 ( .a(n_3727), .o(n_3728) );
in01f80 g742839 ( .a(n_37215), .o(n_37199) );
in01f80 g746309 ( .a(n_33527), .o(n_33528) );
na02f80 g778168 ( .a(FE_OCP_RBN3488_n_3390), .b(FE_OCP_RBN2292_n_2438), .o(n_2813) );
in01f80 g759094 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n_22657) );
na02f80 g770003 ( .a(n_10909), .b(n_10882), .o(n_10991) );
in01f80 g780607 ( .a(n_725), .o(n_726) );
na02f80 g753428 ( .a(n_27020), .b(n_26981), .o(n_27037) );
na02f80 g758204 ( .a(n_22409), .b(n_22372), .o(n_22494) );
in01f80 g772427 ( .a(n_8518), .o(n_8519) );
in01f80 g756318 ( .a(n_24042), .o(n_24068) );
in01f80 g764702 ( .a(n_16447), .o(n_16448) );
na02f80 g743987 ( .a(n_35650), .b(n_35623), .o(n_35792) );
oa22f80 FE_RC_3335_0 ( .a(n_24245), .b(FE_RN_654_0), .c(n_24222), .d(n_24281), .o(n_24426) );
oa12f80 g774897 ( .a(n_6187), .b(n_6237), .c(n_6087), .o(n_6311) );
in01f80 g771792 ( .a(n_9028), .o(n_9029) );
ao12f80 g750989 ( .a(n_30254), .b(n_30207), .c(n_30303), .o(n_31090) );
in01f80 g780284 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_3_), .o(n_1622) );
na02f80 g776993 ( .a(n_3885), .b(n_3884), .o(n_3920) );
na02f80 g770749 ( .a(FE_OCP_RBN3652_n_10100), .b(FE_OCP_RBN2468_n_8767), .o(n_10241) );
in01f80 g762047 ( .a(n_18537), .o(n_18538) );
no02f80 g736667 ( .a(n_43327), .b(n_43325), .o(n_43440) );
in01f80 g774400 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .o(n_6580) );
ao22s80 g762956 ( .a(n_17717), .b(n_17738), .c(n_17645), .d(n_17737), .o(n_17836) );
in01f80 FE_RC_2699_0 ( .a(n_7502), .o(FE_RN_1132_0) );
in01f80 newInst_5 ( .a(newNet_4), .o(newNet_5) );
in01f80 newInst_1868 ( .a(newNet_1867), .o(newNet_1868) );
in01f80 FE_OCP_RBC3011_n_31117 ( .a(FE_OCP_RBN3007_n_31117), .o(FE_OCP_RBN3011_n_31117) );
in01f80 g760646 ( .a(n_19812), .o(n_19753) );
na02f80 g781070 ( .a(cos_out_19), .b(n_43918), .o(n_309) );
ao22s80 g784147 ( .a(n_38193), .b(n_37225), .c(n_38221), .d(n_45894), .o(n_45897) );
in01f80 g743583 ( .a(n_37584), .o(n_37585) );
no02f80 g756023 ( .a(n_25032), .b(n_25122), .o(n_25167) );
na02f80 FE_RC_3009_0 ( .a(n_20459), .b(n_20489), .o(FE_RN_1318_0) );
no02f80 g770680 ( .a(n_10309), .b(FE_OCP_RBN3538_n_8597), .o(n_10349) );
oa12f80 g779519 ( .a(n_1686), .b(n_1739), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_1781) );
no02f80 FE_RC_2337_0 ( .a(FE_RN_893_0), .b(n_18661), .o(FE_RN_894_0) );
in01f80 g740619 ( .a(n_39652), .o(n_39642) );
in01f80 g761716 ( .a(n_19398), .o(n_19399) );
in01f80 g769440 ( .a(FE_OCP_RBN3093_n_11475), .o(n_11556) );
in01f80 g754884 ( .a(n_25394), .o(n_25395) );
na02f80 g767722 ( .a(n_12861), .b(n_12750), .o(n_13019) );
in01f80 g743496 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n_36563) );
no02f80 g749458 ( .a(n_30598), .b(FE_OCPN1410_n_27014), .o(n_30620) );
ao12f80 g764719 ( .a(n_15178), .b(n_15851), .c(FE_OCP_RBN2760_n_15180), .o(n_15852) );
ao12f80 g752023 ( .a(n_28712), .b(n_28711), .c(n_28710), .o(n_29041) );
in01f80 newInst_1958 ( .a(newNet_1957), .o(newNet_1958) );
na02f80 g777760 ( .a(n_3254), .b(n_3233), .o(n_5062) );
oa22f80 FE_RC_3366_0 ( .a(n_22494), .b(n_22574), .c(n_22558), .d(n_22495), .o(n_22715) );
in01f80 g750473 ( .a(n_29589), .o(n_29641) );
na02f80 FE_RC_2336_0 ( .a(FE_RN_892_0), .b(n_18620), .o(FE_RN_893_0) );
in01f80 FE_OCP_RBC2252_n_13017 ( .a(FE_OCP_RBN2251_n_13017), .o(FE_OCP_RBN2252_n_13017) );
no02f80 g763508 ( .a(n_16814), .b(n_16842), .o(n_16903) );
in01f80 FE_OCPC1259_n_25353 ( .a(FE_OCPN1258_n_25353), .o(FE_OCPN1259_n_25353) );
in01f80 newInst_1962 ( .a(newNet_1961), .o(newNet_1962) );
no02f80 g759423 ( .a(n_20991), .b(n_20963), .o(n_21034) );
ao12f80 g739256 ( .a(n_40707), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n_41102) );
na02f80 g769383 ( .a(n_11378), .b(n_10451), .o(n_11454) );
ao22s80 FE_RC_1200_0 ( .a(n_2594), .b(n_3344), .c(n_2595), .d(n_3343), .o(n_3421) );
no02f80 g779369 ( .a(n_1589), .b(n_1390), .o(n_1614) );
in01f80 g759243 ( .a(n_21094), .o(n_21095) );
in01f80 g744138 ( .a(n_35778), .o(n_35779) );
na02f80 g781055 ( .a(cos_out_16), .b(n_43918), .o(n_336) );
no02f80 g784765 ( .a(n_29231), .b(FE_RN_1513_0), .o(n_47251) );
no02f80 g779477 ( .a(n_1581), .b(n_1630), .o(n_1631) );
na02f80 g758900 ( .a(n_46966), .b(n_21728), .o(n_21803) );
in01f80 g750912 ( .a(n_29081), .o(n_29082) );
in01f80 g752496 ( .a(n_28834), .o(n_28396) );
in01f80 g771169 ( .a(n_9761), .o(n_9840) );
in01f80 g771540 ( .a(n_9135), .o(n_9136) );
in01f80 FE_OCP_RBC3819_n_44061 ( .a(FE_OCP_RBN3821_n_44061), .o(FE_OCP_RBN3819_n_44061) );
na02f80 g741909 ( .a(n_38171), .b(n_38090), .o(n_38242) );
in01f80 newInst_264 ( .a(newNet_180), .o(newNet_264) );
no02f80 g756419 ( .a(n_24156), .b(n_24155), .o(n_24259) );
no02f80 g764911 ( .a(FE_OCPN994_n_15552), .b(n_14588), .o(n_15553) );
oa22f80 FE_RC_524_0 ( .a(n_22992), .b(n_22985), .c(n_22993), .d(n_23040), .o(n_23136) );
no02f80 g778903 ( .a(n_2190), .b(n_2179), .o(n_3039) );
in01f80 newInst_3050 ( .a(newNet_3049), .o(newNet_3050) );
in01f80 g760705 ( .a(n_19701), .o(n_19702) );
na02f80 g768532 ( .a(n_12268), .b(n_12164), .o(n_12302) );
in01f80 FE_OCPC877_n_44734 ( .a(FE_OCP_RBN3366_n_44722), .o(FE_OCPN877_n_44734) );
in01f80 newInst_2139 ( .a(newNet_2138), .o(newNet_2139) );
na02f80 g739585 ( .a(FE_OCP_RBN3336_n_44610), .b(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .o(n_40610) );
no02f80 g748576 ( .a(FE_OCP_RBN1211_n_31515), .b(n_31360), .o(n_31588) );
no02f80 g778973 ( .a(n_2101), .b(n_1787), .o(n_2143) );
na02f80 g756749 ( .a(n_23429), .b(n_23428), .o(n_23430) );
oa12f80 g781008 ( .a(n_271), .b(n_273), .c(n_270), .o(n_479) );
in01f80 g761245 ( .a(n_19101), .o(n_19131) );
in01f80 g753594 ( .a(n_26774), .o(n_26775) );
na02f80 g775009 ( .a(n_6113), .b(n_5898), .o(n_6143) );
in01f80 newInst_2714 ( .a(newNet_2713), .o(newNet_2714) );
ao22s80 g775030 ( .a(n_6068), .b(n_5904), .c(n_6067), .d(n_5921), .o(n_6165) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_8_ ( .ck(newNet_3185), .d(n_35874), .o(delay_add_ln22_unr23_stage9_stallmux_q_8_) );
in01f80 g744830 ( .a(n_35219), .o(n_35220) );
oa22f80 FE_RC_4128_0 ( .a(n_22303), .b(n_22544), .c(n_22341), .d(n_22566), .o(n_22684) );
ao12f80 g763318 ( .a(n_16762), .b(n_16793), .c(n_16706), .o(n_16884) );
in01f80 FE_OCP_RBC3113_n_32254 ( .a(n_32254), .o(FE_OCP_RBN3113_n_32254) );
in01f80 g743487 ( .a(n_36626), .o(n_36627) );
na02f80 g774940 ( .a(n_6166), .b(n_6156), .o(n_6267) );
in01f80 FE_OCP_RBC2868_n_16088 ( .a(n_16088), .o(FE_OCP_RBN2868_n_16088) );
ao12f80 g772337 ( .a(n_8607), .b(n_8606), .c(n_8605), .o(n_8688) );
na02f80 FE_RC_2454_0 ( .a(FE_RN_982_0), .b(n_42639), .o(n_42654) );
ao12f80 g752017 ( .a(n_28122), .b(n_28121), .c(n_28120), .o(n_29317) );
na02f80 g741779 ( .a(n_38425), .b(n_38402), .o(n_38403) );
in01f80 newInst_3518 ( .a(newNet_872), .o(newNet_3518) );
in01f80 g776638 ( .a(n_4374), .o(n_4375) );
no02f80 g748878 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n_32441) );
in01f80 g760281 ( .a(n_20340), .o(n_20372) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_17_ ( .ck(newNet_3238), .d(n_36440), .o(delay_add_ln22_unr23_stage9_stallmux_q_17_) );
in01f80 g772211 ( .a(n_8637), .o(n_8669) );
na02f80 g755101 ( .a(n_25178), .b(n_24093), .o(n_25206) );
no02f80 g768123 ( .a(n_12605), .b(delay_add_ln22_unr8_stage4_stallmux_q_18_), .o(n_13412) );
na02f80 g776968 ( .a(n_3886), .b(n_3885), .o(n_3891) );
no02f80 g745853 ( .a(n_34097), .b(n_34096), .o(n_34114) );
na02f80 g753678 ( .a(n_26588), .b(FE_OCPN1526_n_26587), .o(n_26589) );
oa12f80 g738239 ( .a(n_41900), .b(n_41899), .c(n_41898), .o(n_41953) );
in01f80 g739929 ( .a(n_40050), .o(n_40092) );
no02f80 g744894 ( .a(FE_OCP_RBN2644_n_34980), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35032) );
no02f80 FE_RC_4217_0 ( .a(n_15053), .b(FE_RN_1846_0), .o(n_15108) );
na02f80 g759054 ( .a(n_21390), .b(n_45072), .o(n_21497) );
in01f80 g739022 ( .a(n_41218), .o(n_41629) );
in01f80 newInst_312 ( .a(newNet_311), .o(newNet_312) );
na02f80 g741169 ( .a(n_38847), .b(n_38859), .o(n_39061) );
ao12f80 g740715 ( .a(n_39417), .b(n_39416), .c(n_39415), .o(n_39495) );
in01f80 g751543 ( .a(n_28505), .o(n_28493) );
in01f80 g743045 ( .a(n_37176), .o(n_37177) );
in01f80 FE_OCP_RBC2905_n_16197 ( .a(n_16197), .o(FE_OCP_RBN2905_n_16197) );
in01f80 FE_OCPC1391_n_7925 ( .a(n_7925), .o(FE_OCPN1391_n_7925) );
na02f80 g771855 ( .a(n_44516), .b(n_10079), .o(n_10159) );
no02f80 FE_RC_1994_0 ( .a(n_19420), .b(FE_RN_651_0), .o(FE_RN_652_0) );
in01f80 g753093 ( .a(n_27467), .o(n_27468) );
na02f80 g756500 ( .a(n_23873), .b(n_23966), .o(n_23995) );
in01f80 g740349 ( .a(n_40388), .o(n_40389) );
in01f80 g776716 ( .a(n_4080), .o(n_4160) );
na02f80 g771977 ( .a(n_44516), .b(n_9994), .o(n_10154) );
oa12f80 g750961 ( .a(n_28681), .b(n_28934), .c(n_28568), .o(n_28965) );
oa22f80 g752694 ( .a(n_27358), .b(n_27101), .c(n_27359), .d(n_27102), .o(n_27472) );
na02f80 g774831 ( .a(n_45475), .b(n_5648), .o(n_6412) );
in01f80 FE_OCP_RBC2340_n_29470 ( .a(n_29470), .o(FE_OCP_RBN2340_n_29470) );
oa12f80 g759151 ( .a(n_21185), .b(n_21184), .c(n_21183), .o(n_21276) );
in01f80 FE_OCP_RBC2606_FE_OCPN899_n_44593 ( .a(FE_OCPN899_n_44593), .o(FE_OCP_RBN2606_FE_OCPN899_n_44593) );
in01f80 FE_RC_3750_0 ( .a(n_12026), .o(FE_RN_1646_0) );
in01f80 FE_OCP_RBC3719_n_39913 ( .a(FE_OCP_RBN3718_n_39913), .o(FE_OCP_RBN3719_n_39913) );
in01f80 g762686 ( .a(n_17895), .o(n_17923) );
in01f80 g780424 ( .a(n_902), .o(n_934) );
ao12f80 g743757 ( .a(n_36135), .b(n_36074), .c(n_36242), .o(n_36273) );
na02f80 g737511 ( .a(n_42595), .b(n_42520), .o(n_42648) );
in01f80 newInst_143 ( .a(newNet_142), .o(newNet_143) );
no02f80 g779567 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .o(n_1599) );
no02f80 g751694 ( .a(n_28384), .b(n_28361), .o(n_28450) );
no02f80 g776584 ( .a(n_4557), .b(n_4427), .o(n_4451) );
in01f80 g773378 ( .a(n_7612), .o(n_7598) );
na02f80 g739770 ( .a(n_40456), .b(n_40121), .o(n_40462) );
na02f80 g773768 ( .a(n_7159), .b(n_7030), .o(n_7194) );
na02f80 g771593 ( .a(n_8915), .b(FE_OCP_RBN3472_n_7886), .o(n_8946) );
in01f80 g779266 ( .a(n_1822), .o(n_1823) );
na02f80 FE_RC_1832_0 ( .a(n_14201), .b(FE_RN_550_0), .o(FE_RN_551_0) );
na02f80 g741708 ( .a(n_38477), .b(n_38504), .o(n_38573) );
na02f80 g756933 ( .a(n_23803), .b(n_23863), .o(n_23906) );
ao12f80 g759437 ( .a(n_20936), .b(n_20883), .c(n_20849), .o(n_21041) );
na02f80 g742820 ( .a(n_37297), .b(n_37279), .o(n_37310) );
na02f80 g745404 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35840), .o(n_35932) );
na02f80 g756613 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .o(n_23708) );
na02f80 g736944 ( .a(n_43242), .b(n_42883), .o(n_43458) );
in01f80 g765584 ( .a(n_15136), .o(n_15175) );
na02f80 g774953 ( .a(n_6059), .b(n_6055), .o(n_6110) );
no02f80 g780736 ( .a(n_608), .b(n_602), .o(n_603) );
in01f80 g778313 ( .a(n_2847), .o(n_2848) );
oa12f80 g761809 ( .a(n_18700), .b(n_19126), .c(n_18610), .o(n_19229) );
in01f80 FE_OCPC1388_n_11041 ( .a(FE_OCPN1387_n_11041), .o(FE_OCPN1388_n_11041) );
no02f80 g774187 ( .a(n_6872), .b(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .o(n_7141) );
oa12f80 g776528 ( .a(n_4519), .b(n_4518), .c(n_4553), .o(n_4590) );
in01f80 FE_OCP_RBC1155_n_18375 ( .a(FE_OCP_RBN1154_n_18375), .o(FE_OCP_RBN1155_n_18375) );
in01f80 newInst_3309 ( .a(newNet_1562), .o(newNet_3309) );
in01f80 g767401 ( .a(n_13365), .o(n_13385) );
na02f80 g748649 ( .a(n_31400), .b(n_31130), .o(n_31443) );
na02f80 g742401 ( .a(n_37761), .b(n_37724), .o(n_37791) );
no02f80 FE_RC_2647_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_5_), .b(n_32827), .o(FE_RN_1104_0) );
ao12f80 g756948 ( .a(n_23646), .b(n_23802), .c(n_23804), .o(n_23811) );
na02f80 FE_RC_1650_0 ( .a(FE_RN_461_0), .b(n_20854), .o(n_46969) );
no02f80 g761077 ( .a(FE_OCP_RBN1689_n_18986), .b(n_19140), .o(n_19180) );
in01f80 newInst_892 ( .a(newNet_891), .o(newNet_892) );
no02f80 g765158 ( .a(n_15932), .b(n_15832), .o(n_16024) );
in01f80 g736574 ( .a(n_43569), .o(n_43570) );
no02f80 g737372 ( .a(n_42811), .b(n_42340), .o(n_42830) );
no02f80 g773552 ( .a(n_7442), .b(n_7254), .o(n_7477) );
no02f80 g740393 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39538), .o(n_40242) );
in01f80 g778130 ( .a(n_2832), .o(n_2833) );
ao22s80 FE_RC_736_0 ( .a(n_8207), .b(n_7495), .c(n_7494), .d(n_8206), .o(n_8288) );
na02f80 g772884 ( .a(n_7974), .b(n_7973), .o(n_8054) );
no02f80 g750309 ( .a(n_29703), .b(n_29695), .o(n_29732) );
ao12f80 g765998 ( .a(n_14997), .b(n_14996), .c(n_14995), .o(n_15086) );
in01f80 g743794 ( .a(n_36015), .o(n_36047) );
in01f80 g766200 ( .a(n_14556), .o(n_14507) );
in01f80 FE_OCP_RBC1324_n_29056 ( .a(FE_OCP_RBN1323_n_29056), .o(FE_OCP_RBN1324_n_29056) );
in01f80 newInst_2158 ( .a(newNet_2157), .o(newNet_2158) );
na02f80 g761920 ( .a(n_18301), .b(n_18434), .o(n_18319) );
oa12f80 g761841 ( .a(n_18284), .b(n_18595), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n_18641) );
na02f80 g746819 ( .a(n_32919), .b(n_32918), .o(n_33166) );
oa12f80 g757376 ( .a(n_23383), .b(n_23400), .c(n_23382), .o(n_23903) );
in01f80 g761577 ( .a(n_20231), .o(n_22793) );
in01f80 FE_OCP_RBC2721_n_9494 ( .a(n_9494), .o(FE_OCP_RBN2721_n_9494) );
in01f80 g780259 ( .a(n_1010), .o(n_993) );
no02f80 g764457 ( .a(n_16422), .b(n_16266), .o(n_16416) );
no02f80 g774291 ( .a(n_6742), .b(n_6741), .o(n_6743) );
in01f80 FE_OCP_RBC1334_n_20249 ( .a(FE_OCP_RBN1332_n_20249), .o(FE_OCP_RBN1334_n_20249) );
ao12f80 g766902 ( .a(n_13793), .b(n_13848), .c(FE_OCP_RBN1925_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_13943) );
no02f80 g756498 ( .a(n_23922), .b(n_23921), .o(n_23943) );
no02f80 g749622 ( .a(FE_OCP_RBN1357_n_30298), .b(n_30444), .o(n_30446) );
no02f80 g739168 ( .a(n_40938), .b(n_40923), .o(n_40924) );
no02f80 g764425 ( .a(n_16169), .b(n_14650), .o(n_16166) );
no02f80 g750680 ( .a(n_29275), .b(n_28799), .o(n_29326) );
ao22s80 FE_RC_3742_0 ( .a(n_32101), .b(n_32296), .c(n_32102), .d(n_32300), .o(n_32380) );
in01f80 g781313 ( .a(n_53), .o(n_54) );
na02f80 g777129 ( .a(n_3557), .b(n_3444), .o(n_3569) );
na02f80 g755897 ( .a(n_24419), .b(n_25386), .o(n_24420) );
oa22f80 FE_RC_1470_0 ( .a(n_24350), .b(FE_OCP_RBN3132_n_27736), .c(n_27796), .d(n_27736), .o(n_27797) );
in01f80 newInst_3662 ( .a(newNet_3661), .o(newNet_3662) );
na02f80 g779278 ( .a(n_1785), .b(n_1784), .o(n_1919) );
in01f80 FE_OCP_DRV_C1566_n_28654 ( .a(FE_OCP_DRV_N1565_n_28654), .o(FE_OCP_DRV_N1566_n_28654) );
ao12f80 g759086 ( .a(n_21774), .b(n_21909), .c(n_21826), .o(n_22009) );
ao12f80 g752833 ( .a(n_28051), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n_28616) );
na02f80 g745628 ( .a(n_34286), .b(n_34590), .o(n_34648) );
ao12f80 g746336 ( .a(n_33608), .b(n_33607), .c(n_33606), .o(n_33673) );
oa12f80 g757763 ( .a(n_22466), .b(FE_OCP_RBN3106_n_22590), .c(n_22406), .o(n_22661) );
ao22s80 FE_RC_1230_0 ( .a(n_17389), .b(n_17694), .c(n_17324), .d(n_17659), .o(n_17729) );
oa22f80 FE_RC_334_0 ( .a(n_22337), .b(n_22685), .c(n_22336), .d(n_22719), .o(n_22874) );
no02f80 g750778 ( .a(n_30306), .b(n_30290), .o(n_30340) );
no02f80 g745948 ( .a(n_33967), .b(n_34013), .o(n_34053) );
oa12f80 g784647 ( .a(n_16628), .b(n_16607), .c(n_16585), .o(n_46977) );
na02f80 g764307 ( .a(n_16328), .b(n_14524), .o(n_16329) );
na02f80 g742499 ( .a(n_37595), .b(n_37625), .o(n_37662) );
no02f80 g757961 ( .a(n_22850), .b(n_22849), .o(n_22851) );
in01f80 newInst_3443 ( .a(newNet_969), .o(newNet_3443) );
in01f80 FE_RC_272_0 ( .a(FE_RN_83_0), .o(n_22171) );
no02f80 g739956 ( .a(n_40398), .b(n_40176), .o(n_40409) );
in01f80 g741953 ( .a(n_38060), .o(n_38061) );
na02f80 g779625 ( .a(n_1674), .b(n_1681), .o(n_2053) );
no02f80 g770363 ( .a(n_44053), .b(n_10624), .o(n_10626) );
in01f80 g763283 ( .a(n_17272), .o(n_17273) );
na02f80 g752525 ( .a(n_27646), .b(n_27531), .o(n_27701) );
in01f80 FE_OCP_RBC2222_n_13010 ( .a(n_13010), .o(FE_OCP_RBN2222_n_13010) );
in01f80 g738017 ( .a(n_42172), .o(n_42441) );
ao22s80 g736429 ( .a(n_43752), .b(n_43631), .c(FE_OCP_RBN3127_n_43752), .d(n_43630), .o(n_43794) );
na02f80 g758119 ( .a(n_44268), .b(n_22134), .o(n_22225) );
in01f80 newInst_1700 ( .a(newNet_569), .o(newNet_1700) );
oa12f80 g751430 ( .a(n_28458), .b(n_28577), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n_28579) );
in01f80 newInst_3690 ( .a(newNet_3328), .o(newNet_3690) );
na02f80 g770224 ( .a(n_10694), .b(n_10737), .o(n_10786) );
no02f80 g756401 ( .a(n_23640), .b(n_23443), .o(n_23691) );
ao12f80 g755858 ( .a(n_24106), .b(n_24906), .c(n_24154), .o(n_24958) );
oa12f80 g761772 ( .a(n_19161), .b(n_19160), .c(n_19159), .o(n_19760) );
no02f80 g736693 ( .a(n_43366), .b(n_43292), .o(n_43367) );
no02f80 g745939 ( .a(n_34077), .b(n_34111), .o(n_34140) );
oa12f80 g746715 ( .a(n_33007), .b(n_33145), .c(n_32968), .o(n_33204) );
na02f80 g765823 ( .a(n_14917), .b(n_14808), .o(n_14954) );
na02f80 g765965 ( .a(n_14750), .b(n_14679), .o(n_14751) );
no02f80 g764286 ( .a(n_16230), .b(n_14524), .o(n_16446) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_20_ ( .ck(newNet_1405), .d(n_36661), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_) );
in01f80 g740819 ( .a(n_39853), .o(n_39465) );
in01f80 newInst_2434 ( .a(newNet_1156), .o(newNet_2434) );
na02f80 g776641 ( .a(n_4401), .b(n_4400), .o(n_4402) );
oa12f80 g767573 ( .a(n_13056), .b(n_13055), .c(n_13054), .o(n_13222) );
na02f80 g753240 ( .a(n_27377), .b(n_27217), .o(n_27380) );
no02f80 g747255 ( .a(n_32773), .b(delay_add_ln22_unr20_stage8_stallmux_q_2_), .o(n_32817) );
in01f80 FE_OCP_RBC3482_n_13667 ( .a(n_13667), .o(FE_OCP_RBN3482_n_13667) );
in01f80 FE_OCP_DRV_C1576_n_28829 ( .a(FE_OCP_DRV_N1575_n_28829), .o(FE_OCP_DRV_N1576_n_28829) );
in01f80 FE_OFC839_n_4597 ( .a(n_4597), .o(FE_OFN839_n_4597) );
na02f80 g776722 ( .a(n_4213), .b(n_4087), .o(n_4214) );
in01f80 g762237 ( .a(n_18238), .o(n_18239) );
na02f80 g764158 ( .a(n_16852), .b(n_16102), .o(n_16889) );
no02f80 g767441 ( .a(n_13474), .b(n_13473), .o(n_13475) );
in01f80 g740115 ( .a(n_40223), .o(n_40224) );
na02f80 g740849 ( .a(n_39346), .b(n_39345), .o(n_39470) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_18_ ( .ck(newNet_3154), .d(n_40489), .o(delay_add_ln22_unr27_stage10_stallmux_q_18_) );
no02f80 g744847 ( .a(n_35113), .b(FE_OCPN1434_n_30614), .o(n_35138) );
no02f80 g740652 ( .a(FE_OCP_RBN2835_n_39586), .b(n_45840), .o(n_39611) );
no02f80 g774049 ( .a(n_6823), .b(n_6531), .o(n_6889) );
in01f80 g738506 ( .a(n_41635), .o(n_41586) );
in01f80 fopt783923 ( .a(n_45630), .o(n_45629) );
in01f80 newInst_2582 ( .a(newNet_2054), .o(newNet_2582) );
no02f80 g759995 ( .a(n_20532), .b(n_20534), .o(n_20632) );
in01f80 FE_RC_3293_0 ( .a(n_22890), .o(FE_RN_1448_0) );
in01f80 newInst_2835 ( .a(newNet_2834), .o(newNet_2835) );
in01f80 g777242 ( .a(n_5447), .o(n_3620) );
in01f80 g761544 ( .a(n_18864), .o(n_18897) );
na02f80 g744258 ( .a(FE_OCPN1510_n_44174), .b(n_34869), .o(n_36182) );
na02f80 g755889 ( .a(n_25522), .b(n_25548), .o(n_25637) );
in01f80 FE_OCPC1437_FE_OCP_RBN1330_n_18866 ( .a(FE_OCP_RBN1330_n_18866), .o(FE_OCPN1437_FE_OCP_RBN1330_n_18866) );
in01f80 g753237 ( .a(n_27175), .o(n_27219) );
na02f80 g738409 ( .a(n_41475), .b(n_41427), .o(n_41552) );
na02f80 g742554 ( .a(n_37559), .b(FE_OCP_RBN3392_n_37557), .o(n_37576) );
no02f80 g750095 ( .a(n_29841), .b(n_28888), .o(n_29893) );
in01f80 g747307 ( .a(n_32716), .o(n_32717) );
no02f80 g742600 ( .a(n_37554), .b(n_38279), .o(n_37555) );
no02f80 g750861 ( .a(n_29113), .b(n_30364), .o(n_29112) );
in01f80 FE_OCP_RBC1343_n_19077 ( .a(FE_OCP_RBN1342_n_19077), .o(FE_OCP_RBN1343_n_19077) );
no02f80 g748174 ( .a(n_31931), .b(n_32056), .o(n_32132) );
in01f80 g780474 ( .a(n_1159), .o(n_780) );
in01f80 g741650 ( .a(n_38583), .o(n_38587) );
no02f80 g759033 ( .a(n_21959), .b(n_21480), .o(n_21980) );
in01f80 g738753 ( .a(n_41729), .o(n_41600) );
in01f80 g743431 ( .a(n_36614), .o(n_36657) );
oa22f80 g779048 ( .a(FE_OCP_RBN3412_n_2100), .b(n_1876), .c(n_2100), .d(n_1877), .o(n_2173) );
no02f80 g755329 ( .a(n_24934), .b(n_23668), .o(n_24969) );
no02f80 FE_RC_4061_0 ( .a(FE_RN_1767_0), .b(n_36208), .o(n_36280) );
na02f80 g767639 ( .a(n_12745), .b(n_12521), .o(n_12772) );
na02f80 g739297 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_41053) );
in01f80 FE_OCP_RBC1373_n_35275 ( .a(n_35275), .o(FE_OCP_RBN1373_n_35275) );
oa22f80 FE_RC_3740_0 ( .a(n_15610), .b(n_15613), .c(n_15609), .d(n_15615), .o(n_15889) );
in01f80 g756521 ( .a(n_23941), .o(n_23942) );
oa22f80 g784340 ( .a(FE_OFN775_n_46137), .b(n_5538), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5569), .o(n_46146) );
no02f80 g763926 ( .a(n_17018), .b(FE_OCP_RBN3360_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17156) );
in01f80 g761951 ( .a(n_18269), .o(n_18289) );
no02f80 g748024 ( .a(n_31813), .b(n_31523), .o(n_31814) );
na02f80 g752051 ( .a(n_28044), .b(n_28043), .o(n_28332) );
oa12f80 g739845 ( .a(n_40091), .b(n_40265), .c(n_39983), .o(n_40301) );
no02f80 g742896 ( .a(n_37001), .b(n_37016), .o(n_37288) );
na02f80 g752229 ( .a(FE_OCPN877_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .o(n_27972) );
na02f80 g747438 ( .a(n_33746), .b(n_33360), .o(n_33533) );
no02f80 g760348 ( .a(n_18918), .b(n_20184), .o(n_20264) );
no02f80 g751928 ( .a(n_28150), .b(n_28126), .o(n_28228) );
no02f80 g762223 ( .a(n_18116), .b(n_18097), .o(n_18164) );
oa12f80 g778933 ( .a(n_2121), .b(n_2148), .c(n_2120), .o(n_2738) );
in01f80 g772224 ( .a(n_8711), .o(n_8762) );
na02f80 g784769 ( .a(n_34286), .b(FE_OCP_RBN1354_n_33584), .o(n_47255) );
no02f80 g755039 ( .a(n_25233), .b(n_25268), .o(n_25234) );
ao12f80 g738998 ( .a(n_41184), .b(n_41192), .c(n_41183), .o(n_41576) );
in01f80 g746171 ( .a(n_33827), .o(n_33847) );
na02f80 g763681 ( .a(n_16649), .b(n_16397), .o(n_16671) );
in01f80 g768068 ( .a(n_12700), .o(n_12701) );
na02f80 g758613 ( .a(n_21902), .b(FE_OCPN3178_n_21901), .o(n_21922) );
in01f80 g753035 ( .a(n_28336), .o(n_32566) );
no02f80 g755331 ( .a(n_24887), .b(n_24923), .o(n_24939) );
no02f80 FE_RC_3843_0 ( .a(FE_OCP_RBN1150_n_17239), .b(FE_RN_1675_0), .o(n_17341) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_14_ ( .ck(newNet_2115), .d(n_5971), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_14_) );
in01f80 newInst_71 ( .a(newNet_70), .o(newNet_71) );
na02f80 g779164 ( .a(n_1868), .b(n_1745), .o(n_1950) );
in01f80 g761145 ( .a(n_19172), .o(n_19201) );
in01f80 g784709 ( .a(FE_OCP_RBN2821_n_10023), .o(n_47184) );
no02f80 g765534 ( .a(n_15664), .b(n_15663), .o(n_15709) );
na02f80 g744741 ( .a(n_35220), .b(n_30633), .o(n_35285) );
no02f80 g779820 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_27_), .o(n_2109) );
na02f80 g736629 ( .a(n_43442), .b(n_43284), .o(n_43443) );
in01f80 g746842 ( .a(n_33366), .o(n_33367) );
in01f80 g776281 ( .a(n_47008), .o(n_4700) );
in01f80 g741836 ( .a(n_38388), .o(n_38441) );
na02f80 g747479 ( .a(n_32543), .b(n_44962), .o(n_32687) );
in01f80 g750034 ( .a(n_30139), .o(n_30140) );
ao22s80 g750995 ( .a(n_29880), .b(n_179), .c(n_29879), .d(n_186), .o(n_31043) );
na02f80 FE_RC_3849_0 ( .a(FE_RN_1679_0), .b(n_19139), .o(n_19166) );
in01f80 g741770 ( .a(n_38572), .o(n_38473) );
in01f80 g771318 ( .a(n_9148), .o(n_9162) );
in01f80 g769830 ( .a(n_11113), .o(n_11139) );
na02f80 g742942 ( .a(n_37204), .b(n_36944), .o(n_37228) );
ao12f80 g774202 ( .a(n_7121), .b(n_6872), .c(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .o(n_7161) );
in01f80 g742509 ( .a(n_37653), .o(n_37654) );
na02f80 g752011 ( .a(n_28919), .b(n_28691), .o(n_29332) );
in01f80 FE_RC_477_0 ( .a(n_23461), .o(FE_RN_141_0) );
na02f80 g759073 ( .a(n_21527), .b(n_21526), .o(n_21528) );
in01f80 g757208 ( .a(n_23079), .o(n_23080) );
oa22f80 g780532 ( .a(n_890), .b(n_809), .c(n_923), .d(n_620), .o(n_1062) );
no02f80 g771851 ( .a(n_44516), .b(n_10078), .o(n_10120) );
na02f80 FE_RC_4221_0 ( .a(FE_RN_1848_0), .b(FE_RN_1849_0), .o(FE_RN_1850_0) );
na02f80 g742866 ( .a(n_37237), .b(n_37236), .o(n_37238) );
in01f80 FE_OCP_RBC2119_n_45224 ( .a(FE_OCP_RBN2118_n_45224), .o(FE_OCP_RBN2119_n_45224) );
in01f80 g740077 ( .a(n_39919), .o(n_39920) );
no02f80 g775767 ( .a(n_5198), .b(n_5087), .o(n_5344) );
in01f80 FE_OCPC3760_n_2466 ( .a(n_2466), .o(FE_OCPN3760_n_2466) );
in01f80 g744868 ( .a(n_35097), .o(n_35098) );
no02f80 FE_RC_2249_0 ( .a(FE_RN_826_0), .b(FE_RN_827_0), .o(FE_RN_828_0) );
no02f80 g739925 ( .a(n_40436), .b(n_40332), .o(n_40437) );
na02f80 g740441 ( .a(n_39787), .b(n_39539), .o(n_39967) );
na02f80 g737939 ( .a(n_42277), .b(n_42106), .o(n_42296) );
oa12f80 g757893 ( .a(n_22041), .b(n_22172), .c(n_22087), .o(n_22173) );
in01f80 g768709 ( .a(n_12145), .o(n_12102) );
in01f80 FE_OCP_RBC2384_n_8342 ( .a(FE_OCP_RBN2383_n_8342), .o(FE_OCP_RBN2384_n_8342) );
in01f80 g762423 ( .a(n_18414), .o(n_18415) );
in01f80 FE_RC_2436_0 ( .a(n_32711), .o(FE_RN_971_0) );
in01f80 g741179 ( .a(n_38921), .o(n_39056) );
oa22f80 g774265 ( .a(n_6514), .b(n_6408), .c(n_6513), .d(n_6409), .o(n_6670) );
in01f80 newInst_383 ( .a(newNet_156), .o(newNet_383) );
no02f80 g776164 ( .a(n_4860), .b(n_4477), .o(n_4914) );
oa22f80 FE_RC_21_0 ( .a(n_6471), .b(n_6502), .c(n_6488), .d(n_6472), .o(n_6648) );
no02f80 g740892 ( .a(n_39306), .b(n_39270), .o(n_39343) );
in01f80 g778768 ( .a(n_2328), .o(n_2329) );
no02f80 g753867 ( .a(n_26179), .b(n_26302), .o(n_26303) );
in01f80 g740689 ( .a(n_39524), .o(n_39525) );
in01f80 fopt783177 ( .a(n_44718), .o(n_44717) );
na02f80 g744047 ( .a(n_44223), .b(n_34678), .o(n_35831) );
in01f80 g777323 ( .a(n_4598), .o(n_4599) );
na02f80 g743963 ( .a(n_35747), .b(n_34726), .o(n_35748) );
in01f80 g756342 ( .a(n_24000), .o(n_24018) );
na02f80 g760617 ( .a(n_19834), .b(n_19882), .o(n_19939) );
na02f80 g760887 ( .a(n_19505), .b(n_19425), .o(n_19556) );
in01f80 g776353 ( .a(n_4703), .o(n_4704) );
no02f80 g769812 ( .a(n_11192), .b(n_44498), .o(n_11230) );
no02f80 g761790 ( .a(n_19194), .b(n_19193), .o(n_19195) );
na02f80 g736984 ( .a(n_43120), .b(n_42982), .o(n_43389) );
no02f80 g770417 ( .a(FE_OCP_RBN2873_n_10477), .b(FE_OCP_RBN3637_n_44490), .o(n_10510) );
na02f80 g739994 ( .a(n_39955), .b(n_39857), .o(n_40022) );
no02f80 g761184 ( .a(n_19769), .b(n_19713), .o(n_19797) );
in01f80 newInst_35 ( .a(newNet_34), .o(newNet_35) );
ao22s80 g752409 ( .a(n_44723), .b(n_44696), .c(FE_OCP_RBN3306_n_44722), .d(n_44695), .o(n_27888) );
in01f80 g760081 ( .a(n_20294), .o(n_20317) );
ao12f80 FE_RC_3598_0 ( .a(FE_RN_1570_0), .b(FE_RN_1571_0), .c(n_13310), .o(n_13435) );
no02f80 g749856 ( .a(FE_OCP_RBN3018_n_31117), .b(n_31251), .o(n_31322) );
na02f80 g758924 ( .a(n_21604), .b(n_21496), .o(n_21647) );
na02f80 g756543 ( .a(n_23572), .b(n_23611), .o(n_23659) );
no02f80 FE_RC_3718_0 ( .a(FE_RN_1634_0), .b(FE_RN_1635_0), .o(FE_RN_1636_0) );
na02f80 g753837 ( .a(n_26368), .b(n_26303), .o(n_26401) );
na02f80 g748007 ( .a(n_33003), .b(n_32605), .o(n_33043) );
na02f80 g771958 ( .a(FE_OCPN906_n_44561), .b(n_9172), .o(n_9323) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_2_ ( .ck(newNet_1483), .d(n_31293), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_) );
na02f80 g756040 ( .a(n_25026), .b(n_25109), .o(n_25548) );
na02f80 g780599 ( .a(n_745), .b(n_773), .o(n_841) );
no02f80 g753726 ( .a(n_26496), .b(n_26559), .o(n_26624) );
no02f80 g759753 ( .a(n_21172), .b(n_21108), .o(n_21255) );
in01f80 FE_RC_3503_0 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .o(FE_RN_1512_0) );
no02f80 g759346 ( .a(n_20826), .b(FE_OCP_RBN1728_FE_RN_1583_0), .o(n_20944) );
in01f80 newInst_3608 ( .a(newNet_1581), .o(newNet_3608) );
ao12f80 g749741 ( .a(FE_OCP_RBN3012_n_31117), .b(n_31289), .c(n_31288), .o(n_31290) );
oa12f80 g777864 ( .a(n_3196), .b(n_3215), .c(n_2759), .o(n_3271) );
na02f80 g764592 ( .a(n_16504), .b(n_15877), .o(n_16541) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_7_ ( .ck(newNet_1679), .d(n_21933), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_) );
in01f80 g743792 ( .a(n_36047), .o(n_36074) );
na02f80 g768046 ( .a(n_12721), .b(n_12720), .o(n_12774) );
no02f80 g737733 ( .a(n_42392), .b(n_42114), .o(n_42526) );
na02f80 g759682 ( .a(n_21877), .b(n_21106), .o(n_21300) );
in01f80 FE_OCPC954_n_44460 ( .a(FE_OCPN996_n_44460), .o(FE_OCPN954_n_44460) );
in01f80 fopt782742 ( .a(n_17686), .o(n_44153) );
na02f80 FE_RC_2679_0 ( .a(FE_RN_1119_0), .b(FE_RN_1121_0), .o(n_4517) );
in01f80 g754808 ( .a(n_25457), .o(n_25490) );
na02f80 g780710 ( .a(n_628), .b(n_581), .o(n_634) );
oa12f80 g749043 ( .a(n_30855), .b(n_30883), .c(n_29896), .o(n_31001) );
in01f80 g753162 ( .a(n_27482), .o(n_27483) );
in01f80 FE_RC_3728_0 ( .a(n_19064), .o(FE_RN_1640_0) );
in01f80 g775316 ( .a(n_5674), .o(n_5675) );
na02f80 g754494 ( .a(n_26687), .b(n_26741), .o(n_26772) );
in01f80 g754339 ( .a(n_27142), .o(n_25851) );
ao12f80 g741797 ( .a(n_38395), .b(n_38394), .c(n_38393), .o(n_38873) );
ao12f80 g754812 ( .a(n_25116), .b(n_25282), .c(n_25069), .o(n_25366) );
in01f80 g773151 ( .a(n_7824), .o(n_7995) );
no02f80 FE_RC_1785_0 ( .a(FE_RN_520_0), .b(FE_RN_522_0), .o(FE_RN_523_0) );
no02f80 FE_RC_767_0 ( .a(FE_RN_237_0), .b(FE_RN_238_0), .o(FE_RN_239_0) );
no02f80 g778199 ( .a(n_45505), .b(n_2383), .o(n_2742) );
oa12f80 g757915 ( .a(n_21936), .b(n_22086), .c(n_21937), .o(n_22140) );
no02f80 g748684 ( .a(n_31142), .b(n_30996), .o(n_31209) );
ao12f80 g765371 ( .a(n_15667), .b(n_15874), .c(n_15786), .o(n_16508) );
no02f80 g773240 ( .a(n_45616), .b(n_8531), .o(n_7639) );
in01f80 newInst_304 ( .a(newNet_303), .o(newNet_304) );
in01f80 newInst_2859 ( .a(newNet_2858), .o(newNet_2859) );
oa22f80 g779891 ( .a(FE_OCPN875_n_44672), .b(n_1005), .c(n_44623), .d(n_949), .o(n_1297) );
no02f80 g760711 ( .a(n_19736), .b(n_19698), .o(n_19737) );
no02f80 g757899 ( .a(n_22887), .b(n_22730), .o(n_22888) );
no02f80 g754520 ( .a(n_26233), .b(n_26164), .o(n_26313) );
in01f80 g775244 ( .a(n_5959), .o(n_5957) );
in01f80 g738253 ( .a(n_42358), .o(n_41936) );
oa12f80 g757856 ( .a(n_23085), .b(n_23007), .c(FE_OFN735_n_22641), .o(n_23121) );
no02f80 g780914 ( .a(n_420), .b(n_443), .o(n_467) );
na02f80 g761325 ( .a(n_19905), .b(n_19823), .o(n_20512) );
oa22f80 FE_RC_3287_0 ( .a(n_30658), .b(n_30706), .c(n_30657), .d(n_30707), .o(n_30860) );
no02f80 g747748 ( .a(n_33440), .b(n_33462), .o(n_33797) );
in01f80 g738957 ( .a(n_41223), .o(n_41224) );
in01f80 g781239 ( .a(n_138), .o(n_139) );
no02f80 g779104 ( .a(n_2042), .b(n_1770), .o(n_2076) );
oa22f80 g737876 ( .a(n_42270), .b(n_42046), .c(FE_OCPN1231_n_42201), .d(n_42026), .o(n_42612) );
in01f80 g770490 ( .a(n_10320), .o(n_10321) );
in01f80 g758974 ( .a(n_22119), .o(n_22056) );
na02f80 g751746 ( .a(n_29050), .b(n_28990), .o(n_29078) );
na02f80 g759225 ( .a(n_21073), .b(n_45024), .o(n_21222) );
no02f80 g738986 ( .a(n_41204), .b(n_40867), .o(n_41235) );
in01f80 newInst_1058 ( .a(newNet_747), .o(newNet_1058) );
na02f80 g777808 ( .a(FE_OCP_RBN2464_n_4336), .b(n_2913), .o(n_3285) );
in01f80 g746069 ( .a(n_33956), .o(n_33975) );
oa12f80 g737855 ( .a(n_42248), .b(n_42547), .c(n_42232), .o(n_42602) );
in01f80 newInst_3372 ( .a(newNet_3371), .o(newNet_3372) );
in01f80 FE_RC_2410_0 ( .a(n_2005), .o(FE_RN_950_0) );
no02f80 g738411 ( .a(n_41511), .b(n_41548), .o(n_41872) );
in01f80 g770260 ( .a(n_10779), .o(n_10813) );
ao22s80 g773626 ( .a(FE_OCP_RBN2190_n_7346), .b(n_7109), .c(n_7346), .d(n_7108), .o(n_7702) );
in01f80 g744025 ( .a(n_35625), .o(n_36305) );
no02f80 g742745 ( .a(n_37340), .b(n_37339), .o(n_37341) );
no02f80 g752287 ( .a(FE_OCP_RBN2126_n_44734), .b(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .o(n_28219) );
na02f80 g768836 ( .a(n_11978), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_), .o(n_12019) );
oa22f80 FE_RC_3368_0 ( .a(n_30595), .b(FE_OCPN1410_n_27014), .c(FE_OCP_DRV_N3158_n_27062), .d(n_30575), .o(n_30692) );
no02f80 g740262 ( .a(n_40059), .b(n_39989), .o(n_40031) );
no02f80 g774286 ( .a(n_6756), .b(n_6755), .o(n_6813) );
no02f80 g760531 ( .a(n_19924), .b(n_19784), .o(n_19976) );
in01f80 FE_OCP_RBC3622_n_15135 ( .a(FE_OCP_RBN3620_n_15135), .o(FE_OCP_RBN3622_n_15135) );
na02f80 g777935 ( .a(n_47022), .b(FE_OCP_RBN2344_FE_OCPN870_n_2737), .o(n_3132) );
in01f80 newInst_723 ( .a(newNet_722), .o(newNet_723) );
in01f80 g771152 ( .a(n_9362), .o(n_9363) );
in01f80 g761446 ( .a(n_20218), .o(n_20219) );
ao22s80 FE_RC_3_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .b(n_1528), .c(n_1549), .d(n_1590), .o(n_1591) );
no02f80 g760781 ( .a(n_19530), .b(n_19442), .o(n_19570) );
no02f80 g745100 ( .a(n_35749), .b(n_34712), .o(n_34713) );
no02f80 g767021 ( .a(FE_OCP_RBN2457_n_13765), .b(n_13135), .o(n_13902) );
na02f80 g749527 ( .a(n_30389), .b(n_30143), .o(n_30429) );
in01f80 FE_OCP_RBC2626_n_3848 ( .a(n_3848), .o(FE_OCP_RBN2626_n_3848) );
in01f80 FE_OCP_RBC3403_n_28597 ( .a(FE_OCP_RBN2192_n_28597), .o(FE_OCP_RBN3403_n_28597) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_10_ ( .ck(newNet_2794), .d(n_16212), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_10_) );
no02f80 g745456 ( .a(n_34406), .b(n_34382), .o(n_34459) );
in01f80 g758162 ( .a(n_22221), .o(n_22220) );
in01f80 g779487 ( .a(n_2090), .o(n_2091) );
in01f80 g766116 ( .a(n_14706), .o(n_14738) );
in01f80 newInst_2982 ( .a(newNet_1986), .o(newNet_2982) );
in01f80 FE_OCP_RBC2004_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN2004_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
no02f80 g774298 ( .a(n_6688), .b(n_6687), .o(n_7170) );
no02f80 g743376 ( .a(n_36583), .b(n_36750), .o(n_36660) );
in01f80 newInst_1622 ( .a(newNet_1128), .o(newNet_1622) );
no02f80 g746454 ( .a(n_35017), .b(n_34645), .o(n_34646) );
oa12f80 g773624 ( .a(n_7102), .b(FE_OCP_RBN2189_n_7346), .c(n_7068), .o(n_7417) );
no02f80 g762320 ( .a(n_18090), .b(n_17920), .o(n_18135) );
oa12f80 g748206 ( .a(n_32767), .b(n_32766), .c(n_32765), .o(n_33294) );
no02f80 g744717 ( .a(n_35205), .b(n_35230), .o(n_35345) );
in01f80 g739859 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_7_), .o(n_40695) );
in01f80 newInst_2318 ( .a(newNet_866), .o(newNet_2318) );
in01f80 g758873 ( .a(n_22117), .o(n_22209) );
no02f80 g748138 ( .a(n_31903), .b(n_31872), .o(n_31932) );
oa22f80 FE_RC_2767_0 ( .a(n_12899), .b(n_13694), .c(n_13663), .d(n_12898), .o(n_13756) );
in01f80 g774990 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_18_), .o(n_7353) );
in01f80 newInst_3423 ( .a(newNet_3422), .o(newNet_3423) );
in01f80 g759785 ( .a(n_21861), .o(n_21862) );
in01f80 g749917 ( .a(n_30200), .o(n_30201) );
in01f80 newInst_3490 ( .a(newNet_3489), .o(newNet_3490) );
na02f80 g739123 ( .a(n_40979), .b(n_40905), .o(n_41060) );
na02f80 g741156 ( .a(FE_OCP_RBN2635_n_38806), .b(n_38820), .o(n_38834) );
na02f80 FE_RC_2798_0 ( .a(FE_RN_1196_0), .b(n_34574), .o(n_34632) );
na02f80 g766123 ( .a(n_14546), .b(n_44849), .o(n_14602) );
in01f80 FE_RC_2283_0 ( .a(n_33738), .o(FE_RN_854_0) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_17_ ( .ck(newNet_3064), .d(n_1025), .o(delay_add_ln22_unr2_stage2_stallmux_q_17_) );
na02f80 g761374 ( .a(n_18923), .b(n_18947), .o(n_19055) );
no02f80 g741295 ( .a(n_44944), .b(n_38890), .o(n_38927) );
in01f80 g742068 ( .a(n_38005), .o(n_38006) );
in01f80 g774063 ( .a(n_6860), .o(n_6861) );
na02f80 g753213 ( .a(n_27087), .b(n_26011), .o(n_27144) );
in01f80 g750155 ( .a(n_29952), .o(n_29953) );
na02f80 g776346 ( .a(n_4494), .b(n_4398), .o(n_4565) );
in01f80 newInst_1010 ( .a(newNet_1009), .o(newNet_1010) );
na02f80 g781343 ( .a(n_29), .b(beta_4), .o(n_146) );
na02f80 g768015 ( .a(n_12729), .b(n_11528), .o(n_12847) );
in01f80 g772908 ( .a(n_7978), .o(n_7979) );
in01f80 g757805 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_), .o(n_23603) );
ao12f80 g765858 ( .a(n_14662), .b(n_14771), .c(n_14719), .o(n_14862) );
na02f80 FE_RC_1804_0 ( .a(n_23445), .b(n_23330), .o(n_23545) );
na02f80 g741999 ( .a(n_38283), .b(n_38237), .o(n_38337) );
in01f80 newInst_2292 ( .a(newNet_2291), .o(newNet_2292) );
na02f80 g771198 ( .a(n_9111), .b(n_8232), .o(n_9196) );
no02f80 FE_RC_2750_0 ( .a(n_43349), .b(n_43646), .o(FE_RN_1168_0) );
na02f80 g770245 ( .a(n_46989), .b(FE_OCP_RBN2613_n_9075), .o(n_10914) );
in01f80 g780063 ( .a(n_1230), .o(n_1231) );
oa12f80 g743806 ( .a(n_36243), .b(n_35877), .c(n_36185), .o(n_36322) );
in01f80 newInst_1937 ( .a(newNet_1892), .o(newNet_1937) );
no02f80 g776368 ( .a(n_4720), .b(n_4719), .o(n_4774) );
na02f80 g739090 ( .a(n_41051), .b(n_41032), .o(n_41033) );
no02f80 FE_RC_54_0 ( .a(FE_RN_12_0), .b(FE_RN_13_0), .o(FE_RN_14_0) );
in01f80 g762196 ( .a(n_18216), .o(n_18377) );
na02f80 g781294 ( .a(beta_31), .b(beta_9), .o(n_101) );
in01f80 FE_OCP_RBC1850_n_22639 ( .a(n_22639), .o(FE_OCP_RBN1850_n_22639) );
in01f80 newInst_124 ( .a(newNet_123), .o(newNet_124) );
in01f80 FE_OCP_DRV_C3738_n_29439 ( .a(n_29439), .o(FE_OCP_DRV_N3738_n_29439) );
in01f80 g760817 ( .a(n_19617), .o(n_19618) );
na02f80 g765903 ( .a(n_14772), .b(n_14411), .o(n_14804) );
in01f80 g750487 ( .a(n_29564), .o(n_29565) );
in01f80 FE_OCP_RBC3507_n_13860 ( .a(FE_OCP_RBN3505_n_13860), .o(FE_OCP_RBN3507_n_13860) );
no02f80 g746976 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .o(n_32957) );
na02f80 FE_RC_2462_0 ( .a(FE_RN_987_0), .b(n_13906), .o(FE_RN_988_0) );
ao12f80 g775601 ( .a(n_5266), .b(n_5571), .c(n_5358), .o(n_5663) );
in01f80 g745978 ( .a(n_33983), .o(n_33984) );
oa22f80 g769310 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .c(n_10387), .d(FE_OCPN1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12201) );
in01f80 g780056 ( .a(n_1232), .o(n_1233) );
oa12f80 g766909 ( .a(n_13826), .b(n_13825), .c(n_13824), .o(n_13907) );
in01f80 FE_OCP_RBC2926_n_16446 ( .a(n_16446), .o(FE_OCP_RBN2926_n_16446) );
in01f80 g736363 ( .a(n_43809), .o(n_43810) );
na02f80 g777066 ( .a(n_3882), .b(n_3912), .o(n_4063) );
in01f80 g775745 ( .a(n_5418), .o(n_5483) );
in01f80 FE_OCP_RBC2798_n_10106 ( .a(FE_OCP_RBN2796_n_10106), .o(FE_OCP_RBN2798_n_10106) );
na02f80 g744322 ( .a(n_35512), .b(n_34151), .o(n_35545) );
in01f80 FE_OCPC951_n_41540 ( .a(n_41540), .o(FE_OCPN951_n_41540) );
no02f80 g754033 ( .a(n_26085), .b(n_24432), .o(n_26186) );
oa12f80 g738549 ( .a(n_41420), .b(n_41631), .c(n_41576), .o(n_41749) );
ao12f80 g752114 ( .a(n_28262), .b(n_28709), .c(n_28173), .o(n_28754) );
no02f80 g749008 ( .a(n_31094), .b(n_31095), .o(n_31177) );
na02f80 g744785 ( .a(n_35100), .b(n_47233), .o(n_35177) );
in01f80 g768448 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_21_), .o(n_12404) );
no02f80 g748803 ( .a(n_32417), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n_32492) );
oa22f80 g753159 ( .a(n_26993), .b(n_26954), .c(n_26922), .d(n_26955), .o(n_27029) );
na02f80 FE_RC_3092_0 ( .a(n_21497), .b(n_21703), .o(FE_RN_1366_0) );
in01f80 FE_OCP_RBC2979_n_5656 ( .a(n_5656), .o(FE_OCP_RBN2979_n_5656) );
na02f80 g773814 ( .a(n_7129), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_), .o(n_7166) );
na02f80 g745442 ( .a(FE_OCP_RBN2993_n_35539), .b(n_35189), .o(n_35795) );
oa22f80 g748671 ( .a(n_31357), .b(n_31375), .c(n_31399), .d(n_31376), .o(n_31435) );
in01f80 newInst_3702 ( .a(newNet_3701), .o(newNet_3702) );
in01f80 g762438 ( .a(n_18127), .o(n_18146) );
na02f80 g742469 ( .a(n_37623), .b(n_37646), .o(n_37647) );
no02f80 g753774 ( .a(FE_OCP_RBN2884_n_26292), .b(n_26366), .o(n_26447) );
in01f80 g751669 ( .a(FE_OCP_RBN2218_FE_OCPN950_n_28595), .o(n_28817) );
in01f80 g764764 ( .a(n_15704), .o(n_15703) );
in01f80 newInst_1039 ( .a(newNet_432), .o(newNet_1039) );
no02f80 g741064 ( .a(n_39042), .b(FE_OCP_RBN2546_n_44944), .o(n_39157) );
na02f80 g766924 ( .a(n_13973), .b(n_14006), .o(n_14007) );
na02f80 g757599 ( .a(n_23276), .b(n_22812), .o(n_23320) );
oa22f80 g767741 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_29_), .c(n_12823), .d(n_13086), .o(n_13130) );
in01f80 g775502 ( .a(n_5812), .o(n_5879) );
no02f80 g756054 ( .a(n_25188), .b(n_24901), .o(n_25771) );
in01f80 newInst_781 ( .a(newNet_780), .o(newNet_781) );
in01f80 FE_OCPC957_n_39096 ( .a(FE_OCPN956_n_39096), .o(FE_OCPN957_n_39096) );
in01f80 g764937 ( .a(n_15656), .o(n_15549) );
in01f80 g755001 ( .a(n_25270), .o(n_25481) );
na02f80 g759273 ( .a(n_20948), .b(n_20922), .o(n_21046) );
na02f80 g784469 ( .a(n_11364), .b(n_10385), .o(n_46285) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_12_ ( .ck(newNet_1256), .d(n_5399), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_) );
in01f80 g746315 ( .a(n_33655), .o(n_33656) );
oa22f80 g744927 ( .a(n_34906), .b(n_34447), .c(n_34907), .d(n_34448), .o(n_35003) );
in01f80 newInst_1073 ( .a(newNet_1072), .o(newNet_1073) );
ao22s80 FE_RC_1059_0 ( .a(n_11767), .b(n_11994), .c(n_11768), .d(n_11995), .o(n_12195) );
in01f80 newInst_1952 ( .a(newNet_1951), .o(newNet_1952) );
na02f80 g776708 ( .a(n_4041), .b(n_3938), .o(n_4042) );
na02f80 g736567 ( .a(n_43528), .b(n_43530), .o(n_43531) );
in01f80 g756881 ( .a(n_23958), .o(n_23865) );
in01f80 g752564 ( .a(n_27681), .o(n_27682) );
no02f80 g763165 ( .a(n_17787), .b(n_17369), .o(n_17816) );
in01f80 FE_RC_3134_0 ( .a(FE_OCP_RBN2777_n_15595), .o(FE_RN_1389_0) );
in01f80 newInst_1729 ( .a(newNet_1728), .o(newNet_1729) );
na02f80 g743359 ( .a(n_36618), .b(n_36595), .o(n_36675) );
na02f80 g738371 ( .a(n_41636), .b(FE_OCP_RBN2313_n_41420), .o(n_41711) );
na02f80 g775627 ( .a(n_5628), .b(n_47012), .o(n_5783) );
na02f80 g742198 ( .a(n_44872), .b(n_38209), .o(n_37903) );
in01f80 newInst_1035 ( .a(newNet_1034), .o(newNet_1035) );
no02f80 g777938 ( .a(n_2987), .b(n_3138), .o(n_3167) );
oa22f80 FE_RC_1321_0 ( .a(FE_OCP_RBN2580_n_3734), .b(n_3819), .c(n_3817), .d(n_3690), .o(n_3881) );
na02f80 g767972 ( .a(n_12886), .b(n_13196), .o(n_13674) );
no02f80 g759933 ( .a(FE_OCP_RBN3679_n_21051), .b(n_21371), .o(n_21482) );
in01f80 g755081 ( .a(n_25583), .o(n_25584) );
in01f80 g737417 ( .a(n_42796), .o(n_42775) );
na02f80 g748383 ( .a(n_31449), .b(n_31448), .o(n_31475) );
no02f80 g741661 ( .a(n_38573), .b(n_38572), .o(n_38574) );
in01f80 g748299 ( .a(n_31919), .o(n_31920) );
in01f80 newInst_610 ( .a(newNet_609), .o(newNet_610) );
no02f80 g736976 ( .a(FE_OCPN913_n_43022), .b(n_43299), .o(n_43357) );
na02f80 g776562 ( .a(n_4375), .b(n_4387), .o(n_4515) );
in01f80 g778417 ( .a(n_2790), .o(n_3592) );
in01f80 g759406 ( .a(n_20855), .o(n_20856) );
in01f80 newInst_2808 ( .a(newNet_2807), .o(newNet_2808) );
in01f80 newInst_2691 ( .a(newNet_2690), .o(newNet_2691) );
in01f80 g761720 ( .a(n_18653), .o(n_18654) );
no02f80 g776811 ( .a(n_3888), .b(n_3871), .o(n_4015) );
in01f80 g766478 ( .a(FE_OCPN1054_n_14098), .o(n_14514) );
no02f80 g756794 ( .a(n_47245), .b(n_23098), .o(n_23421) );
ao12f80 g742757 ( .a(n_37009), .b(n_37298), .c(n_37131), .o(n_37355) );
oa12f80 g780471 ( .a(n_893), .b(n_816), .c(n_779), .o(n_888) );
in01f80 g777975 ( .a(n_3096), .o(n_3075) );
oa22f80 g749053 ( .a(n_32227), .b(n_31430), .c(n_32245), .d(n_31429), .o(n_32291) );
oa22f80 g780395 ( .a(n_836), .b(n_420), .c(n_846), .d(n_580), .o(n_941) );
ao12f80 g749565 ( .a(n_30378), .b(n_30377), .c(n_30376), .o(n_31770) );
in01f80 g780362 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .o(n_959) );
in01f80 g767936 ( .a(n_12722), .o(n_12723) );
ao22s80 FE_RC_1509_0 ( .a(n_45070), .b(FE_OCP_RBN1711_n_21087), .c(n_45023), .d(n_21087), .o(n_21233) );
na02f80 g769920 ( .a(n_10878), .b(n_44464), .o(n_10912) );
in01f80 g768111 ( .a(n_12755), .o(n_12756) );
no02f80 g736458 ( .a(n_43705), .b(n_43412), .o(n_43744) );
in01f80 g736673 ( .a(n_43369), .o(n_43409) );
no02f80 g770620 ( .a(n_10355), .b(n_10310), .o(n_10356) );
oa12f80 g772911 ( .a(n_7912), .b(n_7865), .c(n_7810), .o(n_7966) );
in01f80 g761448 ( .a(n_19901), .o(n_20112) );
na02f80 g763481 ( .a(FE_OCP_RBN1209_n_16814), .b(FE_OCP_RBN2867_n_16088), .o(n_16948) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_6_ ( .ck(newNet_946), .d(n_22794), .o(delay_xor_ln21_unr15_stage6_stallmux_q_6_) );
in01f80 g775921 ( .a(n_5315), .o(n_5316) );
no02f80 g761862 ( .a(n_18549), .b(n_18548), .o(n_18550) );
na02f80 g764996 ( .a(n_15429), .b(n_14419), .o(n_15504) );
in01f80 g736622 ( .a(n_43240), .o(n_43241) );
oa22f80 g771345 ( .a(FE_OCP_RBN2655_n_9198), .b(FE_OCP_RBN2556_n_44576), .c(n_9198), .d(FE_OCP_RBN3573_n_44563), .o(n_9410) );
no02f80 g764438 ( .a(n_16084), .b(n_14524), .o(n_16125) );
in01f80 FE_OCP_RBC3102_n_27571 ( .a(n_27571), .o(FE_OCP_RBN3102_n_27571) );
in01f80 FE_OCP_RBC1701_n_19353 ( .a(FE_OCP_RBN1700_n_19353), .o(FE_OCP_RBN1701_n_19353) );
na02f80 g774092 ( .a(n_6762), .b(n_6564), .o(n_6957) );
na02f80 g767030 ( .a(n_14758), .b(n_13714), .o(n_14258) );
no02f80 g763193 ( .a(n_17340), .b(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n_17399) );
in01f80 g760309 ( .a(n_20279), .o(n_20280) );
in01f80 FE_OCP_RBC2645_n_34980 ( .a(n_34980), .o(FE_OCP_RBN2645_n_34980) );
no02f80 g757948 ( .a(n_22135), .b(n_44277), .o(n_22233) );
in01f80 g775131 ( .a(n_5997), .o(n_5998) );
oa12f80 g780434 ( .a(n_709), .b(n_708), .c(n_707), .o(n_729) );
in01f80 g745986 ( .a(n_34048), .o(n_34087) );
ao12f80 g784437 ( .a(n_37631), .b(n_36746), .c(n_46197), .o(n_46249) );
na02f80 g738140 ( .a(n_42012), .b(n_41853), .o(n_42040) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_16_ ( .ck(newNet_3067), .d(n_973), .o(delay_add_ln22_unr2_stage2_stallmux_q_16_) );
in01f80 g751126 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30504) );
na02f80 g745840 ( .a(n_44104), .b(FE_OCP_RBN3458_n_33872), .o(n_34338) );
no02f80 g756591 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .o(n_23921) );
in01f80 g766782 ( .a(n_13751), .o(n_13785) );
in01f80 g754893 ( .a(n_25331), .o(n_25398) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_13_ ( .ck(newNet_846), .d(n_1288), .o(delay_xor_ln21_unr3_stage2_stallmux_q_13_) );
in01f80 g767862 ( .a(n_12793), .o(n_12794) );
na02f80 g755137 ( .a(n_25373), .b(n_45633), .o(n_25613) );
no02f80 g754219 ( .a(n_26037), .b(n_23398), .o(n_26136) );
in01f80 g749400 ( .a(n_32006), .o(n_32007) );
ao12f80 g747354 ( .a(n_32662), .b(n_32661), .c(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n_33544) );
in01f80 newInst_3462 ( .a(newNet_1487), .o(newNet_3462) );
na02f80 g745384 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35931), .o(n_35927) );
in01f80 g777334 ( .a(n_5241), .o(n_5298) );
in01f80 newInst_2299 ( .a(newNet_2298), .o(newNet_2299) );
no02f80 g763845 ( .a(n_16645), .b(FE_OCP_RBN3608_n_14905), .o(n_16667) );
in01f80 FE_OCP_RBC3593_n_8902 ( .a(n_8902), .o(FE_OCP_RBN3593_n_8902) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_31_ ( .ck(newNet_2063), .d(n_6774), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_) );
in01f80 newInst_1164 ( .a(newNet_1163), .o(newNet_1164) );
in01f80 g764753 ( .a(n_15845), .o(n_15893) );
na04m80 g742669 ( .a(n_37357), .b(n_37366), .c(n_37353), .d(n_37049), .o(n_37400) );
na02f80 FE_RC_1946_0 ( .a(FE_RN_621_0), .b(n_13866), .o(FE_RN_622_0) );
no02f80 g741746 ( .a(n_38427), .b(n_38426), .o(n_38428) );
no02f80 g778726 ( .a(FE_OCPN871_n_2737), .b(n_2644), .o(n_2803) );
no02f80 g774729 ( .a(n_6294), .b(n_6228), .o(n_6371) );
in01f80 g743054 ( .a(n_37008), .o(n_36952) );
in01f80 g756271 ( .a(n_24670), .o(n_24671) );
in01f80 newInst_3307 ( .a(newNet_3306), .o(newNet_3307) );
na02f80 g755368 ( .a(n_24703), .b(n_24702), .o(n_24787) );
na02f80 g746123 ( .a(n_33852), .b(n_33851), .o(n_33853) );
no02f80 g779781 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .o(n_1415) );
na02f80 g743378 ( .a(n_36566), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36618) );
in01f80 g780145 ( .a(n_1175), .o(n_1176) );
no02f80 g777030 ( .a(n_3777), .b(n_3839), .o(n_4008) );
na02f80 g738185 ( .a(n_41995), .b(n_41986), .o(n_41987) );
na02f80 g745537 ( .a(n_34486), .b(n_34506), .o(n_34507) );
in01f80 newInst_8 ( .a(newNet_7), .o(newNet_8) );
na02f80 g762245 ( .a(n_18578), .b(n_18580), .o(n_18587) );
in01f80 FE_OCP_RBC3799_delay_xor_ln22_unr12_stage5_stallmux_q_0_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_0_), .o(FE_OCP_RBN3799_delay_xor_ln22_unr12_stage5_stallmux_q_0_) );
in01f80 g747572 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .o(n_32912) );
no02f80 g772983 ( .a(n_7753), .b(n_7774), .o(n_7884) );
no02f80 g745076 ( .a(FE_OCP_RBN2575_n_34822), .b(n_34626), .o(n_34927) );
no02f80 g765648 ( .a(n_14988), .b(FE_OCP_RBN2503_n_13896), .o(n_15053) );
no02f80 g771817 ( .a(n_9309), .b(n_9308), .o(n_9310) );
oa22f80 g739776 ( .a(n_40450), .b(n_40394), .c(n_40451), .d(n_40395), .o(n_40490) );
no02f80 g742785 ( .a(n_37287), .b(n_37282), .o(n_37875) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_19_ ( .ck(newNet_2566), .d(n_27643), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_) );
ao22s80 g743575 ( .a(n_36501), .b(n_36196), .c(n_36532), .d(n_36197), .o(n_36559) );
no02f80 g745306 ( .a(n_35582), .b(n_35188), .o(n_35635) );
na02f80 g749934 ( .a(n_30973), .b(n_30972), .o(n_30974) );
ao22s80 g756950 ( .a(n_24188), .b(n_23979), .c(n_24059), .d(n_23954), .o(n_24454) );
na02f80 g740562 ( .a(n_39704), .b(n_38794), .o(n_39722) );
in01f80 FE_RC_1330_0 ( .a(n_39840), .o(FE_RN_393_0) );
in01f80 g779184 ( .a(n_2487), .o(n_1911) );
in01f80 newInst_3016 ( .a(newNet_3015), .o(newNet_3016) );
ao12f80 g742805 ( .a(n_37244), .b(n_37243), .c(n_37242), .o(n_37869) );
in01f80 newInst_448 ( .a(newNet_447), .o(newNet_448) );
no02f80 g759975 ( .a(n_20367), .b(n_45060), .o(n_20416) );
in01f80 g768959 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_22_), .o(n_11868) );
na02f80 g749289 ( .a(n_30656), .b(n_30629), .o(n_30771) );
na02f80 g745758 ( .a(n_35407), .b(n_34806), .o(n_35431) );
na02f80 g770074 ( .a(n_10849), .b(n_10897), .o(n_10930) );
no02f80 g766942 ( .a(n_13974), .b(FE_RN_995_0), .o(n_14530) );
in01f80 g753116 ( .a(n_27348), .o(n_27349) );
na02f80 g738580 ( .a(n_41721), .b(n_41608), .o(n_42014) );
ao12f80 g761290 ( .a(n_20012), .b(n_19952), .c(n_19980), .o(n_20781) );
in01f80 g750046 ( .a(n_29899), .o(n_29870) );
in01f80 g765850 ( .a(n_14923), .o(n_14951) );
no02f80 g775062 ( .a(n_6014), .b(n_6037), .o(n_6132) );
na02f80 g739654 ( .a(n_40546), .b(n_40555), .o(n_40579) );
no02f80 g746693 ( .a(n_33163), .b(n_32996), .o(n_33164) );
oa12f80 g778562 ( .a(n_2304), .b(n_2303), .c(n_2302), .o(n_3058) );
na02f80 g778096 ( .a(n_2940), .b(n_2851), .o(n_3055) );
na02f80 g753912 ( .a(n_27003), .b(n_26645), .o(n_27067) );
na02f80 g751036 ( .a(n_29824), .b(n_29823), .o(n_29825) );
oa22f80 FE_RC_3167_0 ( .a(n_22961), .b(n_22903), .c(n_22833), .d(n_22860), .o(n_22963) );
no02f80 g746491 ( .a(n_34814), .b(n_34810), .o(n_34890) );
no02f80 g774360 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_14_), .o(n_6985) );
in01f80 g744354 ( .a(n_46225), .o(n_36826) );
in01f80 g740804 ( .a(n_39466), .o(n_39467) );
in01f80 newInst_2625 ( .a(newNet_2624), .o(newNet_2625) );
in01f80 FE_OCP_RBC2533_n_47018 ( .a(FE_OCP_RBN2532_n_47018), .o(FE_OCP_RBN2533_n_47018) );
in01f80 g768775 ( .a(n_12037), .o(n_12114) );
in01f80 newInst_2531 ( .a(newNet_2530), .o(newNet_2531) );
in01f80 g768597 ( .a(n_12309), .o(n_12310) );
in01f80 FE_OCP_RBC2632_n_30170 ( .a(n_30170), .o(FE_OCP_RBN2632_n_30170) );
no02f80 g781250 ( .a(n_140), .b(n_73), .o(n_249) );
in01f80 FE_OCP_RBC2353_n_13858 ( .a(FE_OCP_RBN1171_n_13858), .o(FE_OCP_RBN2353_n_13858) );
oa12f80 g739838 ( .a(n_40136), .b(n_40432), .c(n_40066), .o(n_40444) );
na02f80 g740350 ( .a(n_40266), .b(n_39859), .o(n_40388) );
ao12f80 g745147 ( .a(n_34577), .b(n_34576), .c(n_34575), .o(n_35749) );
oa12f80 g775558 ( .a(n_5134), .b(n_5138), .c(n_5041), .o(n_5272) );
na02f80 g778439 ( .a(n_2419), .b(n_2394), .o(n_2395) );
in01f80 g778221 ( .a(n_2753), .o(n_2727) );
in01f80 FE_OCP_RBC2532_n_47018 ( .a(n_47018), .o(FE_OCP_RBN2532_n_47018) );
in01f80 newInst_3198 ( .a(newNet_1975), .o(newNet_3198) );
oa12f80 g767563 ( .a(n_12512), .b(n_12805), .c(n_12483), .o(n_12904) );
in01f80 g774544 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_29_), .o(n_6473) );
oa22f80 g753144 ( .a(n_26991), .b(n_26840), .c(n_26992), .d(n_26839), .o(n_27046) );
in01f80 g780628 ( .a(n_900), .o(n_945) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_22_ ( .ck(newNet_716), .d(n_46186), .o(delay_xor_ln21_unr6_stage3_stallmux_q_22_) );
in01f80 g736865 ( .a(n_43611), .o(n_43612) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_29_ ( .ck(newNet_1970), .d(n_12196), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_) );
na02f80 g776855 ( .a(n_3744), .b(n_3613), .o(n_3775) );
na02f80 g774765 ( .a(n_6364), .b(n_6338), .o(n_6465) );
na02f80 g774931 ( .a(n_6235), .b(n_6218), .o(n_6268) );
in01f80 g743331 ( .a(n_37855), .o(n_37899) );
na02f80 g767748 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n_13126) );
in01f80 FE_RC_1217_0 ( .a(n_33402), .o(FE_RN_366_0) );
no02f80 g745158 ( .a(n_34820), .b(n_34819), .o(n_34821) );
na02f80 g778030 ( .a(n_3018), .b(FE_OCP_RBN2297_n_2438), .o(n_3047) );
no02f80 g773108 ( .a(n_7922), .b(n_7829), .o(n_8494) );
in01f80 FE_OCP_RBC2121_n_45224 ( .a(FE_OCP_RBN2119_n_45224), .o(FE_OCP_RBN2121_n_45224) );
in01f80 g779653 ( .a(n_1798), .o(n_1799) );
na02f80 g761705 ( .a(n_19338), .b(n_18933), .o(n_19403) );
oa22f80 g739274 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_9_), .c(n_45153), .d(n_40499), .o(n_41074) );
no02f80 g737953 ( .a(n_42201), .b(n_42045), .o(n_42368) );
no02f80 g777740 ( .a(n_3405), .b(n_3349), .o(n_3447) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_28_ ( .ck(newNet_1820), .d(n_17014), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_) );
na02f80 g765907 ( .a(n_14880), .b(n_14848), .o(n_14917) );
ao12f80 g749967 ( .a(n_29928), .b(n_29869), .c(n_29898), .o(n_30457) );
in01f80 g775225 ( .a(n_5970), .o(n_5996) );
na02f80 g762293 ( .a(n_18616), .b(n_18728), .o(n_19196) );
in01f80 newInst_2193 ( .a(newNet_2192), .o(newNet_2193) );
oa12f80 g736373 ( .a(n_300), .b(n_43770), .c(FE_OFN3_n_43918), .o(n_43804) );
in01f80 g765353 ( .a(n_15404), .o(n_15405) );
na02f80 g745513 ( .a(n_34383), .b(n_34339), .o(n_34406) );
na02f80 g756819 ( .a(n_23865), .b(n_23909), .o(n_23937) );
no02f80 g762345 ( .a(n_45002), .b(n_18526), .o(n_18726) );
oa22f80 g775946 ( .a(n_4684), .b(n_4533), .c(n_4683), .d(n_4532), .o(n_4858) );
na02f80 g758906 ( .a(n_21677), .b(n_21727), .o(n_21759) );
in01f80 g756425 ( .a(n_24299), .o(n_25001) );
no03m80 FE_RC_2617_0 ( .a(n_12402), .b(n_12136), .c(n_12401), .o(n_12445) );
no02f80 g749358 ( .a(n_30643), .b(FE_OCPN1410_n_27014), .o(n_30674) );
ao22s80 FE_RC_523_0 ( .a(n_23881), .b(n_24209), .c(n_23882), .d(n_24208), .o(n_24293) );
in01f80 FE_OCP_RBC2369_n_38545 ( .a(FE_OCP_RBN2368_n_38545), .o(FE_OCP_RBN2369_n_38545) );
in01f80 newInst_1399 ( .a(newNet_1398), .o(newNet_1399) );
oa12f80 g767421 ( .a(n_13171), .b(n_13472), .c(n_13200), .o(n_13585) );
na02f80 g753482 ( .a(n_26842), .b(n_26497), .o(n_26878) );
in01f80 g742841 ( .a(n_37230), .o(n_37222) );
no02f80 g765190 ( .a(n_15840), .b(n_15839), .o(n_15841) );
oa12f80 g752165 ( .a(n_28590), .b(n_28589), .c(n_28588), .o(n_28664) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_9_ ( .ck(newNet_2431), .d(n_31806), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_9_) );
in01f80 g777251 ( .a(n_3666), .o(n_3667) );
na02f80 g760091 ( .a(n_20537), .b(FE_OCP_RBN3840_n_19513), .o(n_20606) );
oa22f80 g771174 ( .a(n_9297), .b(n_9438), .c(n_9357), .d(n_9368), .o(n_9629) );
in01f80 newInst_2183 ( .a(newNet_2182), .o(newNet_2183) );
na02f80 g761262 ( .a(n_19681), .b(n_19680), .o(n_19682) );
oa12f80 g761220 ( .a(n_19956), .b(n_19931), .c(n_20086), .o(n_20987) );
na02f80 g755614 ( .a(n_24565), .b(n_24527), .o(n_24638) );
no02f80 g747710 ( .a(n_33242), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_33243) );
no02f80 g758898 ( .a(n_21435), .b(n_21434), .o(n_21473) );
no02f80 g779586 ( .a(FE_OCP_RBN3249_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_3_), .o(n_1542) );
no02f80 g751943 ( .a(n_28125), .b(n_28124), .o(n_28147) );
no02f80 g748653 ( .a(n_31209), .b(n_30995), .o(n_31246) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_0_ ( .ck(newNet_936), .d(n_27708), .o(n_44695) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_22_ ( .ck(newNet_1111), .d(n_11068), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_7_ ( .ck(newNet_878), .d(n_32350), .o(delay_xor_ln21_unr21_stage8_stallmux_q_7_) );
na02f80 g762364 ( .a(n_45002), .b(n_18102), .o(n_18617) );
no02f80 g751909 ( .a(n_28919), .b(n_29026), .o(n_29129) );
in01f80 FE_OCP_RBC2792_n_9910 ( .a(n_9910), .o(FE_OCP_RBN2792_n_9910) );
no02f80 g756433 ( .a(n_24109), .b(n_23743), .o(n_24156) );
in01f80 FE_OCP_RBC2897_n_45484 ( .a(n_45484), .o(FE_OCP_RBN2897_n_45484) );
ao22s80 FE_RC_3450_0 ( .a(n_24868), .b(n_25071), .c(n_24869), .d(n_25072), .o(n_25149) );
in01f80 g755512 ( .a(n_24799), .o(n_24798) );
in01f80 g767439 ( .a(n_13358), .o(n_13359) );
no02f80 g765780 ( .a(n_14958), .b(n_14903), .o(n_15019) );
in01f80 FE_OCP_RBC2251_n_13017 ( .a(FE_OCP_RBN2250_n_13017), .o(FE_OCP_RBN2251_n_13017) );
na02f80 g760497 ( .a(n_20001), .b(n_20023), .o(n_20094) );
oa22f80 g769397 ( .a(n_11384), .b(n_10383), .c(n_11385), .d(n_10384), .o(n_11433) );
in01f80 g744627 ( .a(n_36621), .o(n_36622) );
na02f80 g770043 ( .a(n_11106), .b(n_10985), .o(n_11063) );
na02f80 g765520 ( .a(FE_OFN765_n_15670), .b(n_15666), .o(n_15714) );
oa12f80 g748708 ( .a(n_32586), .b(n_32493), .c(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32796) );
in01f80 g757883 ( .a(n_22205), .o(n_22238) );
in01f80 g760394 ( .a(n_20212), .o(n_20203) );
no02f80 g745368 ( .a(FE_OCP_RBN3698_n_35543), .b(n_35763), .o(n_35850) );
in01f80 FE_RC_2024_0 ( .a(FE_RN_673_0), .o(n_14369) );
na02f80 g770585 ( .a(FE_OCP_RBN2794_n_10106), .b(n_8992), .o(n_10280) );
no02f80 g771388 ( .a(n_9093), .b(n_9099), .o(n_9152) );
oa22f80 FE_RC_2111_0 ( .a(n_26456), .b(n_27008), .c(FE_OCP_RBN2938_n_26456), .d(n_27017), .o(n_27083) );
oa12f80 g745348 ( .a(n_35719), .b(FE_OCP_RBN2995_n_35539), .c(n_35678), .o(n_36159) );
in01f80 newInst_2286 ( .a(newNet_2096), .o(newNet_2286) );
in01f80 g779467 ( .a(n_1476), .o(n_1477) );
in01f80 newInst_3577 ( .a(newNet_2344), .o(newNet_3577) );
oa12f80 g757709 ( .a(FE_OCP_RBN3065_n_22170), .b(n_22543), .c(n_22138), .o(n_22564) );
na02f80 FE_RC_2747_0 ( .a(FE_RN_1166_0), .b(n_38906), .o(FE_RN_1167_0) );
no02f80 g767279 ( .a(n_13697), .b(n_13379), .o(n_13698) );
in01f80 g757430 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .o(n_23773) );
in01f80 FE_OCP_RBC2140_FE_OCPN861_n_45450 ( .a(FE_OCPN861_n_45450), .o(FE_OCP_RBN2140_FE_OCPN861_n_45450) );
na02f80 g747717 ( .a(n_32088), .b(n_31808), .o(n_32089) );
no02f80 g749902 ( .a(n_29928), .b(n_29897), .o(n_29929) );
in01f80 newInst_3719 ( .a(newNet_2124), .o(newNet_3719) );
oa12f80 g744632 ( .a(n_35311), .b(n_35345), .c(n_35310), .o(n_35380) );
in01f80 FE_OCP_RBC2622_n_3601 ( .a(n_3601), .o(FE_OCP_RBN2622_n_3601) );
na02f80 g748944 ( .a(n_31198), .b(n_31197), .o(n_31296) );
in01f80 g770021 ( .a(n_10878), .o(n_10879) );
in01f80 FE_OCP_RBC2344_FE_OCPN870_n_2737 ( .a(FE_OCP_RBN2343_FE_OCPN870_n_2737), .o(FE_OCP_RBN2344_FE_OCPN870_n_2737) );
ao12f80 g762009 ( .a(n_18781), .b(n_18780), .c(n_18779), .o(n_19913) );
in01f80 g777539 ( .a(n_4759), .o(n_4675) );
in01f80 g777603 ( .a(n_3545), .o(n_3546) );
oa22f80 FE_RC_3306_0 ( .a(n_36790), .b(n_36758), .c(n_36757), .d(n_36791), .o(n_36845) );
oa22f80 g742040 ( .a(FE_OCP_RBN3441_n_37945), .b(n_37520), .c(FE_OCP_RBN3445_n_37945), .d(n_37499), .o(n_38480) );
no02f80 g778103 ( .a(n_2957), .b(FE_OCP_RBN3488_n_3390), .o(n_2981) );
in01f80 newInst_1355 ( .a(newNet_1354), .o(newNet_1355) );
oa12f80 g772310 ( .a(n_8484), .b(n_8553), .c(n_8423), .o(n_8632) );
no02f80 g740074 ( .a(n_40111), .b(n_40005), .o(n_40006) );
na02f80 g737715 ( .a(n_42394), .b(n_42390), .o(n_42463) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_5_ ( .ck(newNet_2516), .d(n_26761), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_) );
na02f80 g774775 ( .a(n_6344), .b(n_6360), .o(n_6476) );
in01f80 newInst_959 ( .a(newNet_958), .o(newNet_959) );
in01f80 g752965 ( .a(n_28198), .o(n_28173) );
in01f80 FE_OCP_RBC1215_n_20595 ( .a(n_20595), .o(FE_OCP_RBN1215_n_20595) );
na02f80 g776425 ( .a(n_4343), .b(n_4093), .o(n_4397) );
in01f80 g764657 ( .a(n_15908), .o(n_15909) );
in01f80 g743147 ( .a(n_36921), .o(n_36995) );
na02f80 g769801 ( .a(n_11118), .b(n_44464), .o(n_11144) );
oa22f80 FE_RC_201_0 ( .a(n_17313), .b(n_17557), .c(n_17314), .d(n_17558), .o(n_17725) );
in01f80 FE_OCP_RBC2046_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2046_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
na02f80 g740364 ( .a(FE_OCP_RBN3031_n_39942), .b(n_40202), .o(n_40309) );
na02f80 g774756 ( .a(n_6368), .b(n_6268), .o(n_6375) );
in01f80 g759874 ( .a(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_22111) );
na02f80 g769574 ( .a(n_11376), .b(n_47185), .o(n_11476) );
no02f80 g767962 ( .a(n_13079), .b(n_13080), .o(n_13036) );
na02f80 g762216 ( .a(n_18615), .b(n_19400), .o(n_18776) );
in01f80 g751458 ( .a(n_28603), .o(n_28604) );
no02f80 g748069 ( .a(n_32025), .b(n_32059), .o(n_32105) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_3_ ( .ck(newNet_158), .d(n_46383), .o(delay_xor_ln22_unr9_stage4_stallmux_q_3_) );
no02f80 g772333 ( .a(n_8659), .b(n_8628), .o(n_8755) );
in01f80 FE_OCP_RBC2958_n_26231 ( .a(FE_OCP_RBN2955_n_26231), .o(FE_OCP_RBN2958_n_26231) );
in01f80 FE_RC_1233_0 ( .a(n_6389), .o(FE_RN_370_0) );
ao12f80 g780326 ( .a(n_964), .b(n_907), .c(n_1203), .o(n_984) );
in01f80 g737724 ( .a(n_42387), .o(n_42388) );
in01f80 fopt783334 ( .a(n_44869), .o(n_44920) );
in01f80 g775110 ( .a(n_6063), .o(n_6043) );
oa22f80 FE_RC_1691_0 ( .a(FE_OCP_RBN2507_n_13896), .b(n_14768), .c(FE_OCPN1005_n_13962), .d(FE_OCP_RBN2680_n_14768), .o(n_14873) );
no02f80 g772005 ( .a(n_44464), .b(n_9478), .o(n_9695) );
no02f80 FE_RC_3731_0 ( .a(FE_RN_1642_0), .b(n_19566), .o(n_19606) );
in01f80 g737397 ( .a(n_42808), .o(n_42838) );
in01f80 g737405 ( .a(n_42811), .o(n_42806) );
in01f80 g751079 ( .a(n_28894), .o(n_28933) );
in01f80 g766971 ( .a(n_13683), .o(n_13739) );
in01f80 g743033 ( .a(n_37151), .o(n_37152) );
oa12f80 g752691 ( .a(n_28202), .b(n_28129), .c(n_27923), .o(n_28216) );
na02f80 g742130 ( .a(n_38227), .b(n_38230), .o(n_38355) );
in01f80 g756095 ( .a(n_24981), .o(n_24953) );
oa12f80 g780262 ( .a(n_909), .b(n_908), .c(n_1148), .o(n_1018) );
in01f80 g775994 ( .a(n_4815), .o(n_4816) );
in01f80 FE_OCP_RBC2214_FE_OCPN950_n_28595 ( .a(FE_OCP_RBN3406_n_28597), .o(FE_OCP_RBN2214_FE_OCPN950_n_28595) );
na02f80 g760647 ( .a(n_19730), .b(n_18117), .o(n_19812) );
no02f80 g749783 ( .a(n_31407), .b(n_31411), .o(n_31429) );
in01f80 g764182 ( .a(n_16887), .o(n_16888) );
in01f80 newInst_2437 ( .a(newNet_2436), .o(newNet_2437) );
no02f80 g761254 ( .a(n_18951), .b(n_18324), .o(n_18990) );
ao22s80 g764533 ( .a(n_15907), .b(n_15635), .c(n_15857), .d(n_15636), .o(n_16086) );
in01f80 g770101 ( .a(n_10797), .o(n_10778) );
in01f80 newInst_2794 ( .a(newNet_2793), .o(newNet_2794) );
no02f80 g760653 ( .a(n_19802), .b(FE_OCPUNCON1806_n_19801), .o(n_19833) );
oa22f80 g749803 ( .a(n_29835), .b(n_29848), .c(n_29811), .d(n_29796), .o(n_31403) );
in01f80 g770086 ( .a(n_10765), .o(n_10766) );
na02f80 g764615 ( .a(n_15999), .b(n_15903), .o(n_16000) );
in01f80 g749654 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_31778) );
in01f80 g749238 ( .a(n_32174), .o(n_32175) );
na02f80 g762096 ( .a(n_18266), .b(delay_add_ln22_unr11_stage5_stallmux_q_19_), .o(n_18313) );
in01f80 FE_OCP_RBC1920_n_22476 ( .a(FE_OCP_RBN1919_n_22476), .o(FE_OCP_RBN1920_n_22476) );
ao12f80 g737496 ( .a(n_42539), .b(n_42538), .c(n_42537), .o(n_42597) );
in01f80 g747779 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_32276) );
in01f80 g744050 ( .a(n_35696), .o(n_35697) );
ao12f80 g748087 ( .a(n_32628), .b(n_32809), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .o(n_32826) );
no02f80 FE_RC_4230_0 ( .a(n_15225), .b(n_15137), .o(FE_RN_1857_0) );
na03f80 FE_RC_4267_0 ( .a(n_13780), .b(n_13727), .c(n_13731), .o(n_13883) );
in01f80 g744777 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_36497) );
na02f80 g773201 ( .a(n_7817), .b(n_7877), .o(n_7916) );
no02f80 g743829 ( .a(n_36071), .b(n_36039), .o(n_36203) );
no02f80 g760192 ( .a(n_20929), .b(n_20901), .o(n_20902) );
na02f80 g740866 ( .a(n_39288), .b(n_39275), .o(n_39345) );
oa12f80 g767993 ( .a(n_12474), .b(n_12629), .c(n_12432), .o(n_12668) );
oa12f80 g779190 ( .a(n_1792), .b(n_44812), .c(n_1569), .o(n_1894) );
na02f80 g769321 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .o(n_11794) );
oa12f80 g775877 ( .a(n_4802), .b(n_5217), .c(n_4842), .o(n_5346) );
in01f80 FE_RC_2757_0 ( .a(n_18300), .o(FE_RN_1173_0) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_8_ ( .ck(newNet_2334), .d(n_35757), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_) );
na02f80 g769220 ( .a(n_11575), .b(n_11465), .o(n_11629) );
na02f80 g751987 ( .a(n_28793), .b(n_28862), .o(n_28905) );
na02f80 g745803 ( .a(n_44102), .b(n_33499), .o(n_34479) );
na02f80 g778997 ( .a(n_2195), .b(n_2194), .o(n_2196) );
in01f80 newInst_2225 ( .a(newNet_2224), .o(newNet_2225) );
na02f80 g783817 ( .a(n_15392), .b(n_15353), .o(n_45502) );
na02f80 FE_RC_3763_0 ( .a(FE_RN_1653_0), .b(FE_OCPN932_n_40736), .o(n_44026) );
in01f80 FE_RC_3395_0 ( .a(n_16567), .o(FE_RN_1470_0) );
in01f80 FE_OCP_RBC3414_n_12739 ( .a(n_12739), .o(FE_OCP_RBN3414_n_12739) );
no02f80 g742485 ( .a(n_37627), .b(n_37643), .o(n_37702) );
in01f80 FE_RC_2056_0 ( .a(FE_RN_696_0), .o(n_26220) );
na02f80 g739092 ( .a(n_40997), .b(n_40751), .o(n_41031) );
no02f80 g739386 ( .a(n_45181), .b(n_40500), .o(n_40749) );
in01f80 FE_OCP_RBC1185_n_14823 ( .a(n_14823), .o(FE_OCP_RBN1185_n_14823) );
in01f80 g743079 ( .a(n_46254), .o(n_37082) );
ao12f80 g768713 ( .a(n_12031), .b(n_12030), .c(n_12029), .o(n_12134) );
na02f80 g768462 ( .a(n_12378), .b(n_12253), .o(n_12375) );
no02f80 g747377 ( .a(n_32525), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n_32692) );
no02f80 g744688 ( .a(n_35213), .b(n_35183), .o(n_35234) );
in01f80 g752309 ( .a(FE_OFN811_n_29140), .o(n_27961) );
na02f80 g759050 ( .a(n_21466), .b(FE_OCPN1524_n_45072), .o(n_21496) );
ao12f80 g745862 ( .a(n_44100), .b(n_34123), .c(n_34122), .o(n_34135) );
ao12f80 g746325 ( .a(n_33507), .b(n_33506), .c(n_33505), .o(n_34350) );
ao12f80 g779425 ( .a(n_2082), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .o(n_2439) );
no02f80 g779564 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_10_), .o(n_1554) );
in01f80 g781263 ( .a(n_125), .o(n_126) );
oa22f80 g755939 ( .a(n_25160), .b(n_25085), .c(n_25188), .d(n_24382), .o(n_25576) );
in01f80 g758769 ( .a(n_22284), .o(n_22285) );
in01f80 FE_OCP_RBC3623_n_39097 ( .a(n_39097), .o(FE_OCP_RBN3623_n_39097) );
no02f80 g749510 ( .a(n_30529), .b(n_30509), .o(n_30598) );
in01f80 g781392 ( .a(beta_14), .o(n_40) );
oa12f80 g766767 ( .a(n_13099), .b(n_13664), .c(n_13083), .o(n_13709) );
ao12f80 g768242 ( .a(n_12611), .b(n_12623), .c(n_12610), .o(n_12887) );
in01f80 g740961 ( .a(n_39110), .o(n_39111) );
na02f80 FE_RC_2786_0 ( .a(FE_RN_1188_0), .b(FE_RN_1189_0), .o(n_19747) );
oa12f80 g736657 ( .a(n_334), .b(n_43074), .c(FE_OFN5_n_43918), .o(n_43155) );
in01f80 g776270 ( .a(n_4554), .o(n_4555) );
in01f80 FE_OCP_RBC2232_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2232_n_13141) );
oa22f80 g743719 ( .a(n_36276), .b(n_36367), .c(n_36275), .d(n_36368), .o(n_36423) );
no02f80 g769680 ( .a(FE_OCP_RBN3705_n_11146), .b(n_44516), .o(n_11205) );
no02f80 g764324 ( .a(n_16319), .b(FE_OCP_RBN2629_n_14590), .o(n_16438) );
in01f80 g767790 ( .a(n_13120), .o(n_13121) );
in01f80 g753212 ( .a(n_27144), .o(n_27178) );
no02f80 g742187 ( .a(n_44869), .b(n_37875), .o(n_37876) );
in01f80 newInst_2347 ( .a(newNet_2346), .o(newNet_2347) );
no02f80 g751370 ( .a(n_28745), .b(n_28607), .o(n_29036) );
in01f80 newInst_1351 ( .a(newNet_933), .o(newNet_1351) );
in01f80 g748179 ( .a(n_32126), .o(n_32127) );
no02f80 g775660 ( .a(n_5215), .b(n_4759), .o(n_5266) );
na02f80 g765398 ( .a(n_15403), .b(n_15328), .o(n_15449) );
in01f80 newInst_3522 ( .a(newNet_3521), .o(newNet_3522) );
na02f80 FE_RC_2472_0 ( .a(FE_RN_996_0), .b(n_14457), .o(FE_RN_997_0) );
in01f80 g770904 ( .a(n_9942), .o(n_10008) );
no02f80 g736648 ( .a(n_43413), .b(n_43370), .o(n_43441) );
no02f80 g757383 ( .a(n_22828), .b(FE_OCP_RBN3819_n_44061), .o(n_22912) );
no02f80 g738572 ( .a(n_41532), .b(n_41531), .o(n_41569) );
no02f80 g777774 ( .a(n_3347), .b(n_2913), .o(n_3349) );
na02f80 g749840 ( .a(FE_OCP_RBN3013_n_31117), .b(n_31189), .o(n_31185) );
na02f80 g773642 ( .a(n_7342), .b(n_7371), .o(n_7378) );
na02f80 g738011 ( .a(n_42167), .b(n_42165), .o(n_42175) );
in01f80 g762899 ( .a(n_17597), .o(n_17598) );
no02f80 g770049 ( .a(n_10889), .b(n_10835), .o(n_10934) );
in01f80 g750539 ( .a(n_29555), .o(n_29556) );
na02f80 g769943 ( .a(n_10962), .b(FE_OCP_RBN3693_n_10852), .o(n_10977) );
no02f80 g747276 ( .a(n_45753), .b(n_33444), .o(n_33724) );
ms00f80 delay_sub_ln23_0_unr26_stage9_stallmux_q_reg_1_ ( .ck(newNet_1450), .d(n_33337), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_) );
ao12f80 g750663 ( .a(n_30304), .b(n_30337), .c(n_29887), .o(n_30394) );
in01f80 newInst_3451 ( .a(newNet_3450), .o(newNet_3451) );
na02f80 g759309 ( .a(n_21042), .b(n_21041), .o(n_21043) );
in01f80 newInst_3549 ( .a(newNet_3548), .o(newNet_3549) );
no02f80 g749379 ( .a(n_30544), .b(n_30278), .o(n_30609) );
in01f80 g747149 ( .a(n_32708), .o(n_32743) );
no02f80 g777987 ( .a(n_3048), .b(n_2850), .o(n_3100) );
in01f80 g767732 ( .a(n_12846), .o(n_12868) );
ao22s80 FE_RC_1087_0 ( .a(n_29662), .b(n_29808), .c(n_29772), .d(n_29646), .o(n_29839) );
in01f80 g759062 ( .a(n_21280), .o(n_21322) );
in01f80 g773480 ( .a(n_7544), .o(n_7584) );
in01f80 g753643 ( .a(n_26654), .o(n_26655) );
in01f80 newInst_1600 ( .a(newNet_98), .o(newNet_1600) );
na02f80 FE_RC_3524_0 ( .a(FE_RN_1521_0), .b(FE_RN_1523_0), .o(n_34873) );
na02f80 g768592 ( .a(n_12294), .b(n_12293), .o(n_12314) );
no02f80 g780603 ( .a(n_666), .b(n_665), .o(n_682) );
no02f80 g741573 ( .a(n_38627), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38646) );
na02f80 g766425 ( .a(n_14564), .b(n_14108), .o(n_14653) );
in01f80 g780370 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .o(n_892) );
oa12f80 g756955 ( .a(n_23593), .b(n_23592), .c(n_23591), .o(n_24150) );
na02f80 g750576 ( .a(n_29382), .b(n_29403), .o(n_29505) );
in01f80 FE_OCPC3792_n_31804 ( .a(n_31804), .o(FE_OCPN3792_n_31804) );
in01f80 newInst_307 ( .a(newNet_306), .o(newNet_307) );
in01f80 g779681 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .o(n_1366) );
in01f80 g754969 ( .a(n_25212), .o(n_25213) );
no02f80 g743872 ( .a(n_35712), .b(n_35622), .o(n_35832) );
na02f80 g743493 ( .a(n_36519), .b(n_36510), .o(n_36588) );
na02f80 g744579 ( .a(n_35380), .b(n_35379), .o(n_35381) );
in01f80 newInst_363 ( .a(newNet_207), .o(newNet_363) );
in01f80 FE_OCP_RBC2658_n_4101 ( .a(n_4101), .o(FE_OCP_RBN2658_n_4101) );
na02f80 g741629 ( .a(n_38568), .b(n_38778), .o(n_38589) );
no02f80 FE_RC_2642_0 ( .a(n_2913), .b(FE_OCP_RBN2526_n_3421), .o(FE_RN_1102_0) );
na02f80 FE_RC_3926_0 ( .a(n_45622), .b(FE_OCP_RBN3272_n_45224), .o(FE_RN_1698_0) );
in01f80 FE_OFC811_n_29140 ( .a(FE_OFN828_n_29140), .o(FE_OFN811_n_29140) );
no02f80 g765165 ( .a(n_15637), .b(n_15515), .o(n_16347) );
no02f80 g755593 ( .a(n_45633), .b(n_24555), .o(n_24642) );
in01f80 g746783 ( .a(n_33378), .o(n_33379) );
no02f80 g755236 ( .a(n_25607), .b(n_25606), .o(n_25608) );
no02f80 g772655 ( .a(n_8229), .b(FE_OCPN891_n_7802), .o(n_8230) );
in01f80 newInst_3374 ( .a(newNet_1364), .o(newNet_3374) );
oa12f80 g784659 ( .a(n_10719), .b(FE_OCP_RBN2936_n_10626), .c(n_10682), .o(n_46989) );
in01f80 FE_OCP_RBC1199_n_25763 ( .a(n_25763), .o(FE_OCP_RBN1199_n_25763) );
in01f80 g781241 ( .a(n_141), .o(n_142) );
na02f80 g778213 ( .a(n_2792), .b(n_2649), .o(n_2843) );
no02f80 g752822 ( .a(n_27276), .b(n_27234), .o(n_27312) );
na02f80 g764579 ( .a(n_16547), .b(n_16546), .o(n_16548) );
in01f80 FE_RC_2297_0 ( .a(n_25189), .o(FE_RN_865_0) );
in01f80 g741728 ( .a(n_38499), .o(n_38500) );
no02f80 g739200 ( .a(n_40680), .b(n_45180), .o(n_40747) );
na02f80 g777094 ( .a(n_3929), .b(FE_OCP_RBN2582_n_3734), .o(n_4098) );
no02f80 g775041 ( .a(n_5976), .b(n_4759), .o(n_6013) );
ao22s80 FE_RC_2673_0 ( .a(FE_OCP_RBN1137_n_11779), .b(FE_RN_594_0), .c(n_11779), .d(n_11813), .o(n_12036) );
na02f80 g761969 ( .a(n_18911), .b(n_18622), .o(n_18969) );
in01f80 newInst_1810 ( .a(newNet_1809), .o(newNet_1810) );
in01f80 newInst_1644 ( .a(newNet_996), .o(newNet_1644) );
oa22f80 g775363 ( .a(n_5721), .b(n_5463), .c(n_5673), .d(n_5464), .o(n_5840) );
in01f80 g758181 ( .a(n_22020), .o(n_22021) );
ao22s80 g737181 ( .a(n_42984), .b(n_42692), .c(n_42983), .d(n_42691), .o(n_43006) );
in01f80 g778084 ( .a(n_2980), .o(n_3020) );
in01f80 g747454 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_7_), .o(n_32399) );
in01f80 g757135 ( .a(n_24059), .o(n_24188) );
no02f80 g757085 ( .a(n_23301), .b(n_23300), .o(n_23302) );
no02f80 g738455 ( .a(n_41784), .b(n_41763), .o(n_41810) );
no02f80 g747840 ( .a(n_33392), .b(n_33511), .o(n_33701) );
in01f80 newInst_3483 ( .a(newNet_2789), .o(newNet_3483) );
no02f80 g767950 ( .a(n_12918), .b(n_12882), .o(n_12919) );
na02f80 g751179 ( .a(n_29944), .b(n_29992), .o(n_30065) );
na02f80 g760464 ( .a(n_20072), .b(n_18803), .o(n_20144) );
in01f80 g746863 ( .a(n_33066), .o(n_33016) );
oa12f80 g759335 ( .a(n_21208), .b(n_21207), .c(n_21206), .o(n_21302) );
na02f80 g759776 ( .a(n_21297), .b(n_21335), .o(n_21336) );
na02f80 g771948 ( .a(FE_OCP_RBN3644_n_44490), .b(n_9598), .o(n_9811) );
in01f80 FE_RC_2721_0 ( .a(n_8306), .o(FE_RN_1149_0) );
in01f80 newInst_840 ( .a(newNet_839), .o(newNet_840) );
in01f80 FE_RC_1545_0 ( .a(n_28001), .o(FE_RN_436_0) );
no02f80 g739589 ( .a(n_40638), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n_40636) );
na02f80 g770424 ( .a(n_10653), .b(n_10579), .o(n_10684) );
na02f80 g759186 ( .a(n_21095), .b(n_19408), .o(n_21186) );
in01f80 g736345 ( .a(n_43827), .o(n_43828) );
in01f80 newInst_3415 ( .a(newNet_3414), .o(newNet_3415) );
no02f80 g772746 ( .a(n_8169), .b(n_8160), .o(n_8161) );
in01f80 newInst_2641 ( .a(newNet_1232), .o(newNet_2641) );
in01f80 g755921 ( .a(n_24310), .o(n_24386) );
in01f80 g773220 ( .a(n_45887), .o(n_7696) );
no02f80 g778512 ( .a(n_2310), .b(n_2323), .o(n_2475) );
na02f80 g742646 ( .a(n_37400), .b(n_37312), .o(n_37461) );
oa22f80 FE_RC_1598_0 ( .a(n_27481), .b(n_27692), .c(n_27480), .d(n_27717), .o(n_27805) );
in01f80 g738021 ( .a(n_42169), .o(n_42170) );
in01f80 newInst_561 ( .a(newNet_560), .o(newNet_561) );
in01f80 FE_OFC819_n_4298 ( .a(FE_OFN837_n_4298), .o(FE_OFN819_n_4298) );
no02f80 g740019 ( .a(n_40012), .b(FE_OCP_RBN3056_n_39913), .o(n_40083) );
no03m80 g784114 ( .a(n_45858), .b(n_7413), .c(n_6862), .o(n_45864) );
ms00f80 delay_sub_ln23_0_unr29_stage10_stallmux_q_reg ( .ck(newNet_1351), .d(n_45891), .o(delay_sub_ln23_0_unr29_stage10_stallmux_q) );
na02f80 g747477 ( .a(FE_OCP_RBN3333_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .o(n_32368) );
oa22f80 g740993 ( .a(n_38992), .b(n_39051), .c(n_38991), .d(n_39107), .o(n_39785) );
oa12f80 g752491 ( .a(FE_OCPN1448_n_27463), .b(n_44265), .c(n_27415), .o(n_27670) );
in01f80 FE_OCP_RBC3695_n_5284 ( .a(n_5284), .o(FE_OCP_RBN3695_n_5284) );
in01f80 newInst_236 ( .a(newNet_196), .o(newNet_236) );
no02f80 g773730 ( .a(n_7194), .b(n_7190), .o(n_7191) );
ao12f80 g752838 ( .a(n_27881), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n_28276) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_19_ ( .ck(newNet_643), .d(n_46358), .o(delay_xor_ln21_unr9_stage4_stallmux_q_19_) );
na02f80 g763496 ( .a(FE_OCP_RBN1209_n_16814), .b(n_15948), .o(n_16986) );
na02f80 g741405 ( .a(n_38812), .b(n_38068), .o(n_38868) );
in01f80 g742686 ( .a(n_37412), .o(n_37413) );
in01f80 g757339 ( .a(n_23127), .o(n_23128) );
in01f80 newInst_897 ( .a(newNet_896), .o(newNet_897) );
in01f80 g761519 ( .a(FE_OCP_RBN2259_n_18899), .o(n_18944) );
no02f80 FE_RC_3501_0 ( .a(n_27308), .b(n_45766), .o(FE_RN_1511_0) );
no02f80 g770473 ( .a(n_10328), .b(n_10368), .o(n_10478) );
na02f80 g737217 ( .a(n_42908), .b(n_42798), .o(n_42935) );
no02f80 g740528 ( .a(n_39731), .b(n_39723), .o(n_39766) );
na02f80 g751383 ( .a(n_28682), .b(n_28522), .o(n_28683) );
no02f80 g771967 ( .a(FE_OCP_RBN3647_n_44490), .b(n_8689), .o(n_9828) );
in01f80 g755756 ( .a(n_24520), .o(n_24488) );
no02f80 g777297 ( .a(FE_OCP_RBN2727_n_4219), .b(n_4777), .o(n_4864) );
in01f80 FE_OCP_DRV_C1535_n_12633 ( .a(n_12633), .o(FE_OCP_DRV_N1535_n_12633) );
no02f80 g758243 ( .a(n_22455), .b(FE_OFN735_n_22641), .o(n_22734) );
in01f80 newInst_542 ( .a(newNet_541), .o(newNet_542) );
in01f80 g765985 ( .a(n_14696), .o(n_14722) );
in01f80 g773538 ( .a(n_7493), .o(n_7525) );
in01f80 fopt783561 ( .a(n_45180), .o(n_45149) );
na02f80 g743165 ( .a(n_36946), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_6_), .o(n_37084) );
na02f80 g769656 ( .a(n_11333), .b(n_10285), .o(n_11364) );
in01f80 g775851 ( .a(n_5508), .o(n_5509) );
in01f80 FE_RC_2422_0 ( .a(n_6676), .o(FE_RN_959_0) );
in01f80 g741073 ( .a(n_39301), .o(n_39302) );
in01f80 g746881 ( .a(n_33338), .o(n_33339) );
in01f80 g746355 ( .a(n_33616), .o(n_33542) );
oa12f80 g778188 ( .a(n_3209), .b(n_3208), .c(n_3207), .o(n_4018) );
na02f80 g738687 ( .a(n_41716), .b(n_41562), .o(n_41877) );
in01f80 g746621 ( .a(n_34606), .o(n_34607) );
in01f80 g771200 ( .a(n_9570), .o(n_9571) );
in01f80 g762795 ( .a(n_17778), .o(n_17779) );
in01f80 g774132 ( .a(n_6759), .o(n_6833) );
in01f80 g774365 ( .a(n_6656), .o(n_6579) );
no02f80 FE_RC_2564_0 ( .a(FE_RN_1052_0), .b(n_6708), .o(n_6612) );
na02f80 g764732 ( .a(n_15800), .b(n_15701), .o(n_15801) );
ao22s80 g736395 ( .a(n_43782), .b(n_43348), .c(n_43781), .d(n_43347), .o(n_43839) );
in01f80 g748822 ( .a(n_32479), .o(n_32480) );
in01f80 FE_OCPC1032_n_28448 ( .a(FE_OCPN1031_n_28448), .o(FE_OCPN1032_n_28448) );
in01f80 g772298 ( .a(n_8776), .o(n_8777) );
in01f80 g742047 ( .a(n_37984), .o(n_37949) );
in01f80 FE_OCP_RBC3645_n_44490 ( .a(FE_OCP_RBN3641_n_44490), .o(FE_OCP_RBN3645_n_44490) );
oa12f80 g773510 ( .a(n_7506), .b(n_7507), .c(n_7505), .o(n_7676) );
in01f80 g758770 ( .a(n_22246), .o(n_22284) );
in01f80 newInst_1908 ( .a(newNet_1907), .o(newNet_1908) );
in01f80 g767816 ( .a(n_12849), .o(n_12770) );
in01f80 g767607 ( .a(n_13190), .o(n_13262) );
ao12f80 g740692 ( .a(n_39099), .b(n_39450), .c(FE_OCP_RBN3623_n_39097), .o(n_39481) );
in01f80 newInst_1158 ( .a(newNet_368), .o(newNet_1158) );
ao12f80 g756253 ( .a(n_24666), .b(n_24665), .c(n_24664), .o(n_25250) );
in01f80 g756461 ( .a(n_23769), .o(n_23770) );
in01f80 newInst_3363 ( .a(newNet_3362), .o(newNet_3363) );
ao12f80 g772033 ( .a(n_8651), .b(n_8710), .c(n_8652), .o(n_8815) );
no02f80 g741214 ( .a(n_38857), .b(n_38856), .o(n_38858) );
no02f80 g756051 ( .a(n_25026), .b(n_25130), .o(n_25216) );
no02f80 g744605 ( .a(n_35293), .b(n_35292), .o(n_35351) );
in01f80 FE_OCPC966_n_47020 ( .a(FE_OCPN965_n_47020), .o(FE_OCPN966_n_47020) );
na02f80 g755992 ( .a(n_24178), .b(n_21852), .o(n_24229) );
in01f80 newInst_3655 ( .a(newNet_3654), .o(newNet_3655) );
na02f80 g752782 ( .a(n_28196), .b(n_27790), .o(n_28238) );
oa12f80 g738441 ( .a(n_41589), .b(FE_OCPN953_n_41540), .c(n_41637), .o(n_41902) );
no02f80 g779501 ( .a(n_1440), .b(n_1406), .o(n_1529) );
in01f80 g762756 ( .a(n_17997), .o(n_17943) );
ao12f80 g772031 ( .a(n_8151), .b(n_8900), .c(n_8172), .o(n_8962) );
in01f80 g746821 ( .a(n_33196), .o(n_33197) );
no02f80 g777281 ( .a(n_4219), .b(n_4686), .o(n_4731) );
in01f80 newInst_91 ( .a(newNet_90), .o(newNet_91) );
in01f80 FE_RC_2908_0 ( .a(n_13054), .o(FE_RN_1263_0) );
no02f80 g758648 ( .a(n_21744), .b(n_21617), .o(n_21849) );
ao22s80 g774627 ( .a(n_6356), .b(n_6334), .c(n_6357), .d(n_6335), .o(n_6477) );
oa22f80 FE_RC_4122_0 ( .a(n_12681), .b(n_13410), .c(n_12682), .d(n_13411), .o(n_13497) );
na02f80 g774226 ( .a(n_6525), .b(n_6607), .o(n_6649) );
na02f80 g758206 ( .a(n_22410), .b(n_22374), .o(n_22492) );
no02f80 g771990 ( .a(FE_OCP_RBN3548_n_44575), .b(n_9172), .o(n_9225) );
in01f80 FE_RC_4228_0 ( .a(FE_RN_1856_0), .o(FE_OCP_RBN1222_n_45522) );
na02f80 g761760 ( .a(n_18710), .b(n_18472), .o(n_18870) );
ao12f80 g748623 ( .a(n_33028), .b(n_32453), .c(n_46107), .o(n_32723) );
na02f80 g736703 ( .a(n_43112), .b(FE_OCPN912_n_43022), .o(n_43190) );
oa22f80 g750973 ( .a(n_30166), .b(n_30303), .c(n_29883), .d(n_30156), .o(n_31119) );
in01f80 g766150 ( .a(n_14577), .o(n_14598) );
na02f80 g738512 ( .a(FE_OCP_RBN2312_n_41420), .b(n_41626), .o(n_41696) );
oa22f80 g746870 ( .a(FE_OCP_RBN2169_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .c(FE_OCP_RBN2172_n_32892), .d(n_33155), .o(n_33178) );
in01f80 g767689 ( .a(n_12961), .o(n_12962) );
na02f80 g740555 ( .a(n_39629), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39672) );
no02f80 g747119 ( .a(n_32871), .b(n_32716), .o(n_32907) );
oa12f80 g766565 ( .a(n_13981), .b(n_14019), .c(n_14051), .o(n_14052) );
in01f80 FE_OCPC1476_n_23708 ( .a(FE_OCPN1475_n_23708), .o(FE_OCPN1476_n_23708) );
na02f80 g739215 ( .a(n_40814), .b(n_40829), .o(n_40830) );
in01f80 g775158 ( .a(n_6047), .o(n_6005) );
na02f80 g763105 ( .a(n_17507), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .o(n_17619) );
na02f80 g750927 ( .a(n_30229), .b(n_30208), .o(n_30253) );
ao12f80 g744760 ( .a(FE_OCPN1794_n_30612), .b(n_35249), .c(n_35143), .o(n_35283) );
in01f80 FE_OCP_RBC3388_n_33108 ( .a(FE_OCP_RBN3387_n_33108), .o(FE_OCP_RBN3388_n_33108) );
in01f80 g757622 ( .a(n_22684), .o(n_22637) );
no02f80 g742879 ( .a(n_37194), .b(n_37203), .o(n_37249) );
in01f80 FE_OCP_RBC2217_FE_OCPN950_n_28595 ( .a(FE_OCP_RBN2216_FE_OCPN950_n_28595), .o(FE_OCP_RBN2217_FE_OCPN950_n_28595) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_17_ ( .ck(newNet_834), .d(n_1343), .o(delay_xor_ln21_unr3_stage2_stallmux_q_17_) );
no02f80 g758752 ( .a(n_21618), .b(n_21617), .o(n_21709) );
no02f80 g746253 ( .a(n_33570), .b(n_33550), .o(n_33664) );
in01f80 g737586 ( .a(n_42767), .o(n_42768) );
in01f80 newInst_1586 ( .a(newNet_1585), .o(newNet_1586) );
in01f80 g777837 ( .a(n_3232), .o(n_3202) );
in01f80 g771873 ( .a(n_9036), .o(n_9051) );
oa12f80 g748733 ( .a(n_31140), .b(n_31139), .c(n_31138), .o(n_31182) );
na02f80 g776435 ( .a(n_4379), .b(FE_OCP_RBN2691_FE_OCPN843_n_3912), .o(n_4546) );
in01f80 g763233 ( .a(n_17561), .o(n_17410) );
in01f80 FE_RC_2066_0 ( .a(n_34955), .o(FE_RN_702_0) );
na02f80 g741025 ( .a(n_38880), .b(n_38886), .o(n_38932) );
no02f80 g757985 ( .a(n_22308), .b(n_22130), .o(n_22309) );
in01f80 FE_OCP_RBC1693_n_19052 ( .a(FE_OCPN1738_n_19052), .o(FE_OCP_RBN1693_n_19052) );
no02f80 g746955 ( .a(n_33014), .b(delay_add_ln22_unr20_stage8_stallmux_q_10_), .o(n_33032) );
na02f80 g773720 ( .a(n_8174), .b(n_7364), .o(n_7357) );
no02f80 g758300 ( .a(FE_OCPN991_n_22249), .b(n_21283), .o(n_22435) );
no02f80 FE_RC_2852_0 ( .a(n_13887), .b(n_14104), .o(FE_RN_1228_0) );
in01f80 newInst_3479 ( .a(newNet_3478), .o(newNet_3479) );
in01f80 g754366 ( .a(n_25845), .o(n_25846) );
no02f80 g778176 ( .a(n_2853), .b(n_2852), .o(n_2854) );
no02f80 g770154 ( .a(n_10770), .b(n_10390), .o(n_10771) );
na02f80 g746607 ( .a(n_34473), .b(n_34585), .o(n_34609) );
no02f80 g747959 ( .a(n_32081), .b(n_31860), .o(n_32142) );
in01f80 newInst_1258 ( .a(newNet_1257), .o(newNet_1258) );
ao12f80 g760048 ( .a(n_20037), .b(n_21050), .c(n_21019), .o(n_21141) );
oa12f80 g770111 ( .a(n_10347), .b(n_10770), .c(n_10768), .o(n_10798) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_2_ ( .ck(newNet_3018), .d(n_835), .o(delay_add_ln22_unr2_stage2_stallmux_q_2_) );
in01f80 g772459 ( .a(n_8515), .o(n_8516) );
no02f80 FE_RC_3629_0 ( .a(FE_RN_1589_0), .b(n_20951), .o(FE_RN_1590_0) );
na02f80 g757443 ( .a(n_22822), .b(n_22930), .o(n_22964) );
no02f80 g755692 ( .a(n_25343), .b(n_25220), .o(n_25344) );
ao12f80 g752626 ( .a(n_28243), .b(n_28242), .c(n_28241), .o(n_28862) );
in01f80 g758866 ( .a(n_21503), .o(n_21504) );
in01f80 FE_OCP_RBC3822_n_44061 ( .a(FE_OCP_RBN3823_n_44061), .o(FE_OCP_RBN3822_n_44061) );
in01f80 g759604 ( .a(n_20767), .o(n_20764) );
na02f80 g751511 ( .a(n_28469), .b(n_28504), .o(n_28779) );
na02f80 g751659 ( .a(n_28383), .b(n_28360), .o(n_28419) );
in01f80 g745327 ( .a(n_36217), .o(n_36218) );
na02f80 g764633 ( .a(n_16071), .b(FE_OCP_RBN2483_n_14326), .o(n_16107) );
in01f80 newInst_2543 ( .a(newNet_2542), .o(newNet_2543) );
in01f80 g767921 ( .a(n_12799), .o(n_12798) );
no02f80 g750327 ( .a(n_29672), .b(n_45758), .o(n_29688) );
no02f80 g772728 ( .a(n_8227), .b(n_8226), .o(n_8313) );
oa22f80 FE_RC_1583_0 ( .a(n_17584), .b(n_17687), .c(n_16339), .d(n_17649), .o(n_17752) );
oa12f80 g743561 ( .a(n_36199), .b(n_36532), .c(n_36531), .o(n_36546) );
no02f80 g756763 ( .a(n_23424), .b(delay_add_ln22_unr14_stage6_stallmux_q_12_), .o(n_23443) );
na02f80 g767389 ( .a(n_13406), .b(n_13405), .o(n_13433) );
in01f80 g773494 ( .a(n_7465), .o(n_7466) );
no02f80 g762262 ( .a(n_18499), .b(n_18498), .o(n_18500) );
na02f80 g755685 ( .a(n_24500), .b(n_24498), .o(n_24499) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_0_ ( .ck(newNet_280), .d(n_46172), .o(delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
in01f80 newInst_1122 ( .a(newNet_1043), .o(newNet_1122) );
in01f80 g737521 ( .a(n_42594), .o(n_42595) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_9_ ( .ck(newNet_1937), .d(n_10680), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_) );
in01f80 newInst_3135 ( .a(newNet_3134), .o(newNet_3135) );
in01f80 newInst_3161 ( .a(newNet_3160), .o(newNet_3161) );
no02f80 g736689 ( .a(n_43471), .b(n_43470), .o(n_43472) );
no02f80 g758911 ( .a(n_21610), .b(n_21638), .o(n_21764) );
in01f80 fopt783150 ( .a(n_1282), .o(n_44672) );
in01f80 g755470 ( .a(n_24656), .o(n_24657) );
no02f80 FE_RC_4181_0 ( .a(FE_RN_1821_0), .b(n_33827), .o(FE_RN_1828_0) );
na02f80 g746603 ( .a(n_34473), .b(n_34696), .o(n_34694) );
in01f80 newInst_451 ( .a(newNet_450), .o(newNet_451) );
oa12f80 g773653 ( .a(n_7315), .b(n_7314), .c(n_7313), .o(n_7794) );
na02f80 g757499 ( .a(n_22827), .b(delay_add_ln22_unr14_stage6_stallmux_q_1_), .o(n_22867) );
no02f80 FE_RC_3107_0 ( .a(n_26799), .b(n_26692), .o(FE_RN_1374_0) );
oa22f80 g778017 ( .a(n_3076), .b(n_3058), .c(FE_OCP_RBN2462_n_3076), .d(n_3125), .o(n_3152) );
no02f80 g771051 ( .a(n_9419), .b(n_8362), .o(n_9420) );
in01f80 g757184 ( .a(n_23215), .o(n_23232) );
no02f80 g761788 ( .a(n_18894), .b(n_18559), .o(n_18560) );
no02f80 FE_RC_3624_0 ( .a(FE_RN_1586_0), .b(n_20771), .o(FE_RN_1587_0) );
na02f80 g741654 ( .a(n_38580), .b(n_38778), .o(n_38597) );
in01f80 g774970 ( .a(n_6237), .o(n_6257) );
no02f80 FE_RC_2973_0 ( .a(FE_RN_1300_0), .b(n_44222), .o(n_35693) );
ao12f80 g778754 ( .a(n_2185), .b(n_2184), .c(n_2183), .o(n_2719) );
no02f80 g768754 ( .a(n_12030), .b(n_12029), .o(n_12031) );
na02f80 FE_RC_1823_0 ( .a(FE_RN_544_0), .b(n_35275), .o(n_35290) );
no02f80 g781078 ( .a(n_262), .b(n_46), .o(n_263) );
no02f80 g763731 ( .a(n_17211), .b(n_17260), .o(n_17470) );
in01f80 g739755 ( .a(n_40473), .o(n_40474) );
no02f80 g745259 ( .a(n_35807), .b(n_35715), .o(n_35808) );
in01f80 g768688 ( .a(n_47211), .o(n_12185) );
in01f80 g775014 ( .a(n_6179), .o(n_6180) );
no02f80 g767286 ( .a(n_13499), .b(FE_OCP_RBN2271_n_13489), .o(n_13552) );
no02f80 g772254 ( .a(n_8733), .b(n_8173), .o(n_8759) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_28_ ( .ck(newNet_1489), .d(n_32341), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_) );
in01f80 newInst_2574 ( .a(newNet_2573), .o(newNet_2574) );
in01f80 g772484 ( .a(n_8474), .o(n_8513) );
oa22f80 FE_RC_1302_0 ( .a(n_3615), .b(n_3616), .c(n_3610), .d(n_3029), .o(n_3776) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_3_ ( .ck(newNet_495), .d(n_22671), .o(delay_xor_ln22_unr15_stage6_stallmux_q_3_) );
na02f80 FE_RC_2819_0 ( .a(n_34297), .b(FE_RN_1207_0), .o(FE_RN_1208_0) );
na02f80 g736933 ( .a(n_43038), .b(n_46942), .o(n_43092) );
in01f80 FE_OCP_RBC1370_n_20763 ( .a(FE_OCP_RBN1369_n_20763), .o(FE_OCP_RBN1370_n_20763) );
in01f80 newInst_1613 ( .a(newNet_729), .o(newNet_1613) );
oa22f80 g750028 ( .a(n_29869), .b(n_29485), .c(n_29896), .d(n_29507), .o(n_30367) );
in01f80 FE_OCP_RBC3713_n_31466 ( .a(FE_OCP_RBN3712_n_31466), .o(FE_OCP_RBN3713_n_31466) );
ms00f80 mux_while_ln12_psv_q_reg_5_ ( .ck(newNet_108), .d(n_213), .o(mux_while_ln12_psv_q_5_) );
na02f80 g751608 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n_28815) );
na02f80 g746317 ( .a(n_33545), .b(n_34296), .o(n_33546) );
in01f80 g767763 ( .a(n_13356), .o(n_13277) );
no02f80 FE_RC_3453_0 ( .a(n_26394), .b(FE_RN_1484_0), .o(FE_RN_1485_0) );
ao12f80 g746564 ( .a(n_34758), .b(n_34810), .c(n_34229), .o(n_35434) );
na02f80 g773166 ( .a(n_7802), .b(n_7853), .o(n_7880) );
in01f80 newInst_3532 ( .a(newNet_3531), .o(newNet_3532) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_5_ ( .ck(newNet_1071), .d(n_9957), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_) );
oa22f80 FE_RC_3117_0 ( .a(n_45091), .b(FE_OCP_RBN1721_n_21004), .c(n_45024), .d(n_21004), .o(n_21157) );
no02f80 g759356 ( .a(n_21006), .b(n_45091), .o(n_21039) );
na02f80 FE_RC_2777_0 ( .a(FE_RN_1184_0), .b(n_38342), .o(FE_RN_1185_0) );
in01f80 newInst_3616 ( .a(newNet_3545), .o(newNet_3616) );
in01f80 g758735 ( .a(n_21833), .o(n_21834) );
in01f80 g780980 ( .a(n_403), .o(n_420) );
na02f80 g764967 ( .a(n_15316), .b(FE_RN_1314_0), .o(n_15353) );
in01f80 g775181 ( .a(n_5839), .o(n_5868) );
na02f80 g746983 ( .a(n_32892), .b(n_32363), .o(n_32911) );
oa22f80 g757941 ( .a(n_22021), .b(n_21938), .c(n_22020), .d(n_21939), .o(n_22112) );
na02f80 g752046 ( .a(n_28142), .b(n_28094), .o(n_28161) );
oa12f80 g739048 ( .a(n_41152), .b(n_41151), .c(n_41150), .o(n_41542) );
na02f80 g759344 ( .a(n_21061), .b(n_21062), .o(n_21148) );
no02f80 g763122 ( .a(n_17343), .b(n_17444), .o(n_17445) );
na02f80 g762876 ( .a(n_17842), .b(n_17744), .o(n_17889) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_23_ ( .ck(newNet_2550), .d(n_27720), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_) );
na02f80 g778907 ( .a(n_2177), .b(n_2176), .o(n_2178) );
no02f80 g741687 ( .a(n_38534), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38552) );
no02f80 g773429 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n_7555) );
oa12f80 g768406 ( .a(n_12115), .b(n_12418), .c(n_12007), .o(n_12443) );
ao12f80 g761529 ( .a(n_19543), .b(n_19542), .c(n_19541), .o(n_19648) );
in01f80 FE_OCP_RBC2776_n_15110 ( .a(n_15110), .o(FE_OCP_RBN2776_n_15110) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_2_ ( .ck(newNet_1373), .d(n_36281), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_) );
no02f80 g779595 ( .a(FE_OCP_RBN3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n_1494) );
na02f80 g744263 ( .a(n_44180), .b(n_35611), .o(n_35547) );
in01f80 newInst_3420 ( .a(newNet_3419), .o(newNet_3420) );
in01f80 g737460 ( .a(n_42654), .o(n_42655) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_9_ ( .ck(newNet_1060), .d(n_10295), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_) );
ao22s80 g736291 ( .a(FE_OCP_RBN3111_n_43871), .b(n_43559), .c(n_43871), .d(n_43558), .o(n_43900) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_7_ ( .ck(newNet_2234), .d(n_40416), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_) );
in01f80 g746363 ( .a(n_33545), .o(n_34347) );
ao12f80 g768612 ( .a(n_12200), .b(n_12199), .c(n_12198), .o(n_12738) );
no02f80 g755346 ( .a(n_24891), .b(FE_OCPN1512_n_22280), .o(n_24917) );
in01f80 g751618 ( .a(n_28484), .o(n_28485) );
ms00f80 sin_out_reg_22_ ( .ck(newNet_53), .d(n_43898), .o(sin_out_22) );
na02f80 g769863 ( .a(n_44454), .b(n_11078), .o(n_11150) );
no02f80 g739229 ( .a(n_40765), .b(n_40862), .o(n_41248) );
na02f80 g780080 ( .a(n_1213), .b(n_1212), .o(n_1214) );
na02f80 g738337 ( .a(n_41476), .b(n_41523), .o(n_41524) );
na02f80 g768290 ( .a(n_12538), .b(n_12537), .o(n_12576) );
in01f80 FE_OCP_RBC3123_n_6557 ( .a(n_6557), .o(FE_OCP_RBN3123_n_6557) );
in01f80 g769703 ( .a(n_11359), .o(n_11360) );
oa12f80 g766619 ( .a(n_14262), .b(n_14261), .c(n_14260), .o(n_15631) );
no02f80 g744127 ( .a(n_35531), .b(n_35554), .o(n_35555) );
in01f80 g740637 ( .a(n_40028), .o(n_39612) );
na02f80 g744450 ( .a(n_35472), .b(n_35486), .o(n_35512) );
na02f80 g774797 ( .a(n_45475), .b(n_5732), .o(n_6353) );
in01f80 g751707 ( .a(n_28417), .o(n_28418) );
na02f80 g753983 ( .a(n_26201), .b(n_26110), .o(n_26247) );
ao22s80 g739139 ( .a(n_40990), .b(n_41036), .c(n_40975), .d(n_41037), .o(n_41406) );
na02f80 g770565 ( .a(FE_OCP_RBN3666_n_10106), .b(n_9041), .o(n_10282) );
in01f80 newInst_2682 ( .a(newNet_2120), .o(newNet_2682) );
oa12f80 g739689 ( .a(n_40375), .b(n_40524), .c(n_40138), .o(n_40534) );
in01f80 newInst_3399 ( .a(newNet_3398), .o(newNet_3399) );
no02f80 g762375 ( .a(FE_OFN750_n_45003), .b(n_18574), .o(n_18737) );
na02f80 g761832 ( .a(n_18481), .b(n_18479), .o(n_18480) );
oa22f80 g752845 ( .a(n_27047), .b(n_27005), .c(n_27013), .d(n_27004), .o(n_27059) );
oa22f80 g758560 ( .a(n_22488), .b(n_21827), .c(n_22487), .d(n_21828), .o(n_22568) );
in01f80 g754556 ( .a(n_26574), .o(n_26575) );
no02f80 g765036 ( .a(n_15206), .b(FE_OCP_RBN2507_n_13896), .o(n_15241) );
oa12f80 g764670 ( .a(n_16032), .b(n_16031), .c(n_16030), .o(n_16106) );
no02f80 g738352 ( .a(n_41773), .b(n_41752), .o(n_41791) );
in01f80 newInst_697 ( .a(newNet_198), .o(newNet_697) );
in01f80 g738151 ( .a(n_42115), .o(n_42049) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_8_ ( .ck(newNet_1063), .d(n_10168), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_) );
no02f80 g743341 ( .a(n_36716), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36752) );
no02f80 g777266 ( .a(n_3543), .b(n_3601), .o(n_3640) );
in01f80 g764668 ( .a(n_15989), .o(n_15990) );
in01f80 g759606 ( .a(n_21724), .o(n_21725) );
no02f80 g748871 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_24_), .o(n_32489) );
in01f80 g749514 ( .a(n_31939), .o(n_31940) );
no02f80 g749872 ( .a(n_31311), .b(n_30971), .o(n_31407) );
na02f80 g779522 ( .a(n_1404), .b(n_1382), .o(n_1478) );
in01f80 g772816 ( .a(n_8251), .o(n_8137) );
na02f80 g756771 ( .a(n_23476), .b(n_23475), .o(n_23541) );
no02f80 g762090 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n_18590) );
na02f80 g779304 ( .a(n_1699), .b(n_1656), .o(n_1696) );
in01f80 FE_OCP_RBC3543_n_44575 ( .a(n_44575), .o(FE_OCP_RBN3543_n_44575) );
na02f80 g762278 ( .a(n_18620), .b(n_18580), .o(n_18993) );
in01f80 g755262 ( .a(n_25038), .o(n_25039) );
no02f80 g751758 ( .a(n_28306), .b(n_28305), .o(n_28320) );
in01f80 newInst_3056 ( .a(newNet_3055), .o(newNet_3056) );
na02f80 g751861 ( .a(n_28191), .b(n_28189), .o(n_28190) );
na02f80 g765796 ( .a(n_15093), .b(n_15092), .o(n_15094) );
in01f80 g758231 ( .a(n_22808), .o(n_22917) );
in01f80 g753451 ( .a(n_26918), .o(n_26958) );
in01f80 FE_OCP_RBC3485_n_13667 ( .a(FE_OCP_RBN3483_n_13667), .o(FE_OCP_RBN3485_n_13667) );
in01f80 g760809 ( .a(n_20180), .o(n_21169) );
no02f80 g749860 ( .a(FE_OCP_RBN3019_n_31117), .b(n_31184), .o(n_31279) );
na02f80 g777652 ( .a(n_3474), .b(n_3473), .o(n_3505) );
ao12f80 g761827 ( .a(n_18583), .b(n_19097), .c(n_18657), .o(n_19160) );
na02f80 g771371 ( .a(n_9485), .b(n_9378), .o(n_9588) );
no02f80 g760795 ( .a(n_19516), .b(n_19224), .o(n_19603) );
in01f80 newInst_3070 ( .a(newNet_2275), .o(newNet_3070) );
oa12f80 g755771 ( .a(n_24343), .b(n_24342), .c(n_24341), .o(n_24432) );
no02f80 g746992 ( .a(n_34075), .b(n_34074), .o(n_34107) );
in01f80 g757038 ( .a(n_23834), .o(n_23779) );
in01f80 g740870 ( .a(n_39440), .o(n_39376) );
in01f80 g738524 ( .a(n_41546), .o(n_41510) );
na02f80 g778948 ( .a(n_2264), .b(n_2263), .o(n_2280) );
na02f80 g765569 ( .a(n_15103), .b(n_15250), .o(n_15252) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_14_ ( .ck(newNet_586), .d(n_17754), .o(delay_xor_ln22_unr12_stage5_stallmux_q_14_) );
na02f80 g770836 ( .a(n_10182), .b(n_10139), .o(n_10140) );
in01f80 g775567 ( .a(n_5676), .o(n_5748) );
no02f80 g750822 ( .a(n_29154), .b(FE_OCP_RBN2235_n_29055), .o(n_29186) );
in01f80 FE_RC_1532_0 ( .a(n_28092), .o(FE_RN_432_0) );
oa12f80 g742697 ( .a(n_37327), .b(n_37326), .c(n_37325), .o(n_37852) );
in01f80 g775943 ( .a(n_4903), .o(n_4904) );
in01f80 newInst_2832 ( .a(newNet_2468), .o(newNet_2832) );
in01f80 g747081 ( .a(n_33015), .o(n_33034) );
in01f80 FE_OCP_RBC2584_n_3858 ( .a(n_3858), .o(FE_OCP_RBN2584_n_3858) );
na02f80 g762117 ( .a(n_19402), .b(n_18767), .o(n_18883) );
in01f80 newInst_521 ( .a(newNet_520), .o(newNet_521) );
in01f80 FE_RC_2618_0 ( .a(n_40572), .o(FE_RN_1090_0) );
no02f80 g775269 ( .a(n_5600), .b(n_5574), .o(n_5750) );
in01f80 g763409 ( .a(n_17072), .o(n_17073) );
no02f80 g742986 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n_37001) );
in01f80 g767336 ( .a(n_13547), .o(n_13568) );
in01f80 FE_OCP_RBC3587_n_47016 ( .a(n_47016), .o(FE_OCP_RBN3587_n_47016) );
ao22s80 g784424 ( .a(n_36354), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_46236) );
no02f80 g776774 ( .a(n_3913), .b(n_3680), .o(n_3961) );
in01f80 g779264 ( .a(n_1865), .o(n_1866) );
no02f80 g756725 ( .a(n_24036), .b(n_23984), .o(n_24107) );
no02f80 g760157 ( .a(n_20537), .b(n_19503), .o(n_20556) );
na02f80 g766188 ( .a(n_14998), .b(n_14733), .o(n_14734) );
oa12f80 g739179 ( .a(n_40800), .b(n_40801), .c(n_40799), .o(n_41383) );
oa12f80 g745197 ( .a(n_35770), .b(n_35810), .c(FE_OCP_RBN2988_n_35539), .o(n_36230) );
no02f80 g776937 ( .a(n_4023), .b(n_4022), .o(n_4065) );
in01f80 FE_OCPC1054_n_14098 ( .a(FE_OCPN1053_n_14098), .o(FE_OCPN1054_n_14098) );
na02f80 g738601 ( .a(n_41443), .b(n_41398), .o(n_41508) );
no02f80 g745746 ( .a(n_34161), .b(n_34179), .o(n_34603) );
ao12f80 g772828 ( .a(n_7721), .b(n_7959), .c(n_8021), .o(n_8073) );
ao12f80 g739246 ( .a(n_40861), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n_41272) );
in01f80 FE_OCPC1009_n_28439 ( .a(FE_OCPN1008_n_28439), .o(FE_OCPN1009_n_28439) );
in01f80 FE_RC_2899_0 ( .a(n_20124), .o(FE_RN_1256_0) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_10_ ( .ck(newNet_526), .d(n_22872), .o(delay_xor_ln22_unr15_stage6_stallmux_q_10_) );
na02f80 g738426 ( .a(n_41740), .b(n_41605), .o(n_41768) );
in01f80 g739461 ( .a(n_40837), .o(n_40838) );
no02f80 g747836 ( .a(n_33372), .b(n_33573), .o(n_33680) );
na02f80 g779110 ( .a(n_1943), .b(n_1815), .o(n_2009) );
no02f80 FE_RC_2304_0 ( .a(FE_RN_870_0), .b(FE_RN_871_0), .o(FE_RN_872_0) );
in01f80 newInst_327 ( .a(newNet_326), .o(newNet_327) );
no02f80 g752577 ( .a(n_28298), .b(n_28280), .o(n_28281) );
ao12f80 g774219 ( .a(n_6770), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .o(n_6855) );
in01f80 g779313 ( .a(n_1753), .o(n_1754) );
na02f80 g776785 ( .a(n_3867), .b(FE_OCP_RBN2583_n_3734), .o(n_3868) );
in01f80 newInst_1793 ( .a(newNet_1792), .o(newNet_1793) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_7_ ( .ck(newNet_944), .d(n_22766), .o(delay_xor_ln21_unr15_stage6_stallmux_q_7_) );
in01f80 g761354 ( .a(n_19072), .o(n_19073) );
in01f80 g779802 ( .a(n_1433), .o(n_1403) );
no02f80 g743384 ( .a(n_36615), .b(n_36750), .o(n_36616) );
ao12f80 g784620 ( .a(n_39494), .b(n_39408), .c(n_39455), .o(n_46949) );
na02f80 g774811 ( .a(n_6290), .b(n_5852), .o(n_6364) );
in01f80 g763976 ( .a(n_17783), .o(n_17815) );
no02f80 g737606 ( .a(n_42334), .b(n_42374), .o(n_42375) );
no02f80 g779038 ( .a(n_2153), .b(n_2112), .o(n_2587) );
oa12f80 g745035 ( .a(n_34238), .b(n_34753), .c(n_47254), .o(n_34793) );
na02f80 g756486 ( .a(FE_OCP_RBN2275_n_24077), .b(n_24111), .o(n_24112) );
in01f80 FE_OCP_RBC1678_n_44847 ( .a(n_44847), .o(FE_OCP_RBN1678_n_44847) );
na02f80 g764683 ( .a(n_15765), .b(n_14419), .o(n_15999) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_12_ ( .ck(newNet_590), .d(n_17677), .o(delay_xor_ln22_unr12_stage5_stallmux_q_12_) );
in01f80 newInst_2556 ( .a(newNet_2555), .o(newNet_2556) );
ao12f80 g746409 ( .a(n_33083), .b(n_33331), .c(n_33067), .o(n_33427) );
na02f80 g768306 ( .a(n_12607), .b(n_12411), .o(n_12644) );
in01f80 g767111 ( .a(FE_OCP_RBN2506_n_13896), .o(n_14758) );
ao12f80 g773570 ( .a(n_7429), .b(n_45865), .c(n_7428), .o(n_7908) );
na02f80 g744934 ( .a(n_34932), .b(FE_OCPN1796_n_30546), .o(n_34959) );
in01f80 newInst_1590 ( .a(newNet_1589), .o(newNet_1590) );
no02f80 g757021 ( .a(n_23700), .b(n_23800), .o(n_23747) );
no02f80 g738078 ( .a(FE_OCP_RBN2444_n_42051), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42098) );
in01f80 g748888 ( .a(n_32413), .o(n_32487) );
oa22f80 g779867 ( .a(n_44652), .b(n_1188), .c(n_44637), .d(n_1186), .o(n_1329) );
in01f80 g762139 ( .a(n_18843), .o(n_18844) );
in01f80 FE_RC_900_0 ( .a(n_30292), .o(FE_RN_264_0) );
in01f80 FE_OCP_RBC2164_n_28249 ( .a(n_28249), .o(FE_OCP_RBN2164_n_28249) );
no02f80 g760867 ( .a(n_20057), .b(n_20069), .o(n_20121) );
in01f80 FE_OCP_RBC2820_n_4872 ( .a(n_4872), .o(FE_OCP_RBN2820_n_4872) );
no02f80 FE_RC_2290_0 ( .a(FE_RN_859_0), .b(n_17663), .o(FE_RN_860_0) );
in01f80 g741234 ( .a(n_39173), .o(n_39174) );
oa12f80 g776512 ( .a(n_4090), .b(n_4432), .c(n_3990), .o(n_4608) );
na02f80 g762996 ( .a(n_17646), .b(n_17671), .o(n_17762) );
no02f80 g759193 ( .a(n_20982), .b(n_20981), .o(n_21164) );
in01f80 FE_OFC788_n_25834 ( .a(FE_OFN786_n_25834), .o(FE_OFN788_n_25834) );
no02f80 g784125 ( .a(n_7212), .b(n_7211), .o(n_45872) );
na02f80 g763740 ( .a(n_17532), .b(n_17466), .o(n_18255) );
in01f80 FE_OFC50_n_1045 ( .a(FE_OFN49_n_1045), .o(FE_OFN50_n_1045) );
ao22s80 g739694 ( .a(n_40550), .b(n_40213), .c(n_40543), .d(n_40212), .o(n_40574) );
na02f80 g754146 ( .a(n_25920), .b(n_23259), .o(n_25947) );
no02f80 g748713 ( .a(n_31202), .b(n_31201), .o(n_31244) );
no02f80 g781214 ( .a(n_120), .b(n_119), .o(n_121) );
in01f80 g770024 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_12_), .o(n_12462) );
in01f80 g748833 ( .a(n_31297), .o(n_31298) );
na02f80 g777823 ( .a(n_3227), .b(n_2804), .o(n_3291) );
in01f80 newInst_2120 ( .a(newNet_441), .o(newNet_2120) );
in01f80 g755499 ( .a(n_24800), .o(n_24820) );
ao22s80 g751519 ( .a(n_28460), .b(n_27834), .c(n_28467), .d(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_28822) );
in01f80 FE_OCP_RBC2796_n_10106 ( .a(FE_OCP_RBN2794_n_10106), .o(FE_OCP_RBN2796_n_10106) );
in01f80 FE_RC_4246_0 ( .a(FE_RN_1868_0), .o(n_26987) );
in01f80 g779675 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n_1371) );
oa12f80 g745219 ( .a(n_34521), .b(n_34520), .c(n_34519), .o(n_35648) );
na02f80 g778956 ( .a(n_2228), .b(n_1141), .o(n_2324) );
no02f80 g741059 ( .a(n_39097), .b(n_38608), .o(n_39132) );
no02f80 g753421 ( .a(n_27192), .b(n_26918), .o(n_27021) );
no02f80 g751191 ( .a(n_29837), .b(n_29359), .o(n_30256) );
oa12f80 g784799 ( .a(n_16372), .b(n_16322), .c(n_16274), .o(n_47340) );
oa22f80 g739780 ( .a(n_40442), .b(n_40356), .c(n_40443), .d(n_40355), .o(n_40486) );
in01f80 g761900 ( .a(n_18637), .o(n_18638) );
no02f80 g762925 ( .a(n_17797), .b(n_17745), .o(n_17842) );
ao22s80 g736591 ( .a(n_43376), .b(n_43633), .c(n_43377), .d(n_43632), .o(n_43656) );
ao22s80 g738842 ( .a(n_41300), .b(n_41309), .c(n_41310), .d(n_40657), .o(n_42204) );
na02f80 g766898 ( .a(n_13647), .b(FE_OCP_DRV_N1538_n_13646), .o(n_13705) );
na02f80 g747829 ( .a(n_33372), .b(n_33371), .o(n_33390) );
in01f80 FE_OCP_RBC3676_n_21039 ( .a(n_21039), .o(FE_OCP_RBN3676_n_21039) );
in01f80 FE_RC_2717_0 ( .a(FE_OCPN891_n_7802), .o(FE_RN_1146_0) );
in01f80 FE_RC_3056_0 ( .a(n_26804), .o(FE_RN_1339_0) );
ao12f80 g745108 ( .a(n_34655), .b(n_34767), .c(n_34539), .o(n_34788) );
no02f80 g748128 ( .a(n_31987), .b(FE_OCP_RBN3735_n_31819), .o(n_32059) );
in01f80 g773922 ( .a(n_7031), .o(n_7094) );
na02f80 g759126 ( .a(n_21909), .b(n_21957), .o(n_21958) );
in01f80 g743399 ( .a(n_36715), .o(n_36716) );
ao12f80 g741851 ( .a(n_38384), .b(n_38383), .c(n_38382), .o(n_38484) );
ao12f80 g760414 ( .a(n_19958), .b(n_20655), .c(n_19926), .o(n_20782) );
in01f80 FE_OCPC935_n_42192 ( .a(n_42192), .o(FE_OCPN935_n_42192) );
na02f80 g762256 ( .a(n_18535), .b(n_18534), .o(n_18536) );
no02f80 g756394 ( .a(n_24014), .b(n_23945), .o(n_24015) );
in01f80 g767884 ( .a(n_12766), .o(n_12791) );
na02f80 g762885 ( .a(n_17766), .b(n_17719), .o(n_17794) );
in01f80 FE_OFC767_n_15670 ( .a(FE_OFN763_n_15670), .o(FE_OFN767_n_15670) );
no02f80 g749264 ( .a(n_30677), .b(n_45489), .o(n_30741) );
in01f80 g736914 ( .a(n_43110), .o(n_43136) );
in01f80 g770676 ( .a(n_10264), .o(n_10265) );
in01f80 g753894 ( .a(n_26392), .o(n_26393) );
in01f80 FE_RC_3595_0 ( .a(n_13272), .o(FE_RN_1569_0) );
na02f80 g737015 ( .a(n_43230), .b(n_43494), .o(n_43495) );
no02f80 g773465 ( .a(n_7500), .b(delay_add_ln22_unr5_stage3_stallmux_q_24_), .o(n_7511) );
na02f80 g748582 ( .a(n_31404), .b(FE_OCPN1520_n_31403), .o(n_31467) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_7_ ( .ck(newNet_1360), .d(n_36384), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_) );
in01f80 g780168 ( .a(n_1124), .o(n_1100) );
no02f80 g750430 ( .a(n_29594), .b(n_29630), .o(n_29595) );
oa22f80 FE_RC_333_0 ( .a(n_22387), .b(n_22603), .c(n_22340), .d(n_22619), .o(n_22778) );
na02f80 g755784 ( .a(n_24313), .b(n_23971), .o(n_24398) );
in01f80 g769416 ( .a(n_11453), .o(n_11422) );
in01f80 newInst_425 ( .a(newNet_424), .o(newNet_425) );
in01f80 g748369 ( .a(n_32750), .o(n_32780) );
in01f80 g781172 ( .a(n_182), .o(n_178) );
in01f80 g756645 ( .a(n_23600), .o(n_23601) );
in01f80 newInst_3313 ( .a(newNet_3312), .o(newNet_3313) );
no02f80 g766959 ( .a(n_13637), .b(FE_RN_1222_0), .o(n_13685) );
in01f80 g747701 ( .a(n_33420), .o(n_33464) );
oa22f80 g784561 ( .a(FE_OFN800_n_46285), .b(n_10848), .c(FE_OCP_RBN3709_n_46337), .d(n_10814), .o(n_46382) );
ao12f80 g754309 ( .a(n_25723), .b(n_25870), .c(n_25751), .o(n_25954) );
na02f80 g747155 ( .a(n_32906), .b(delay_add_ln22_unr20_stage8_stallmux_q_6_), .o(n_32925) );
no02f80 g752340 ( .a(n_44723), .b(delay_xor_ln21_unr18_stage7_stallmux_q_5_), .o(n_28092) );
oa12f80 g738300 ( .a(n_41837), .b(n_41836), .c(n_41835), .o(n_42286) );
oa12f80 g762810 ( .a(n_17235), .b(n_17694), .c(n_17120), .o(n_17693) );
in01f80 newInst_1675 ( .a(newNet_1674), .o(newNet_1675) );
ao12f80 g784681 ( .a(n_3974), .b(n_3905), .c(n_3835), .o(n_47011) );
no02f80 g778914 ( .a(n_2284), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .o(n_2314) );
oa12f80 g736519 ( .a(n_287), .b(n_43662), .c(FE_OFN2_n_43918), .o(n_43702) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_21_ ( .ck(newNet_3619), .d(n_17460), .o(delay_add_ln22_unr11_stage5_stallmux_q_21_) );
in01f80 g766675 ( .a(n_15564), .o(n_14354) );
no02f80 g777612 ( .a(n_3419), .b(n_2681), .o(n_3480) );
na02f80 g767481 ( .a(n_13234), .b(n_13154), .o(n_13294) );
in01f80 g742238 ( .a(n_38078), .o(n_38134) );
no02f80 g737248 ( .a(n_42898), .b(n_42765), .o(n_42919) );
na02f80 g750090 ( .a(n_29841), .b(n_29866), .o(n_29868) );
no02f80 g736435 ( .a(n_43762), .b(n_43636), .o(n_43783) );
in01f80 g779693 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_3_), .o(n_1364) );
ao12f80 g746511 ( .a(n_34666), .b(n_34938), .c(n_34889), .o(n_34913) );
na02f80 g773704 ( .a(n_7273), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_16_), .o(n_7337) );
no02f80 g759764 ( .a(n_21378), .b(n_20485), .o(n_21337) );
no02f80 g750560 ( .a(n_29475), .b(n_29351), .o(n_29494) );
na02f80 g774926 ( .a(n_6150), .b(n_6197), .o(n_6215) );
no02f80 g751301 ( .a(n_29675), .b(n_29098), .o(n_29721) );
in01f80 fopt783920 ( .a(n_38671), .o(n_45623) );
in01f80 g775405 ( .a(n_5767), .o(n_5768) );
in01f80 g751870 ( .a(n_28293), .o(n_28264) );
in01f80 g737639 ( .a(n_42825), .o(n_42826) );
no02f80 g756458 ( .a(n_23580), .b(n_23613), .o(n_23614) );
in01f80 g738880 ( .a(n_41258), .o(n_41259) );
in01f80 g741872 ( .a(n_38483), .o(n_39230) );
in01f80 g766402 ( .a(n_15666), .o(n_14652) );
na02f80 FE_RC_1729_0 ( .a(n_23456), .b(FE_RN_479_0), .o(FE_RN_480_0) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_28_ ( .ck(newNet_2732), .d(n_17688), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_) );
in01f80 g776821 ( .a(n_47013), .o(n_4076) );
na02f80 g758514 ( .a(n_21940), .b(n_21922), .o(n_21941) );
in01f80 g754977 ( .a(n_25128), .o(n_25185) );
na02f80 g773838 ( .a(n_7054), .b(delay_add_ln22_unr5_stage3_stallmux_q_11_), .o(n_7117) );
in01f80 FE_OCP_RBC3572_n_44563 ( .a(n_44563), .o(FE_OCP_RBN3572_n_44563) );
na02f80 g766431 ( .a(n_14147), .b(n_14230), .o(n_14268) );
no02f80 g757495 ( .a(n_22990), .b(n_22932), .o(n_23040) );
na02f80 g757058 ( .a(n_24188), .b(n_24087), .o(n_24352) );
in01f80 newInst_382 ( .a(newNet_381), .o(newNet_382) );
na02f80 g753169 ( .a(n_27414), .b(n_27381), .o(n_27521) );
in01f80 g778788 ( .a(n_2365), .o(n_2414) );
oa12f80 g779330 ( .a(n_1452), .b(n_1635), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(n_1636) );
na02f80 g760912 ( .a(n_19381), .b(n_19430), .o(n_19431) );
na02f80 g771701 ( .a(n_8786), .b(n_8795), .o(n_8881) );
in01f80 g781339 ( .a(n_72), .o(n_73) );
na02f80 g739892 ( .a(n_40124), .b(n_39922), .o(n_40265) );
in01f80 g775984 ( .a(n_5288), .o(n_5289) );
in01f80 FE_OCP_RBC2625_n_3848 ( .a(n_3848), .o(FE_OCP_RBN2625_n_3848) );
na02f80 g740922 ( .a(n_39114), .b(n_39277), .o(n_39336) );
no02f80 g760120 ( .a(FE_OCP_RBN3850_n_20290), .b(n_20187), .o(n_20314) );
no02f80 g775868 ( .a(n_5248), .b(n_5184), .o(n_5249) );
na02f80 FE_RC_2996_0 ( .a(n_6412), .b(n_6535), .o(FE_RN_1310_0) );
in01f80 g774807 ( .a(n_6272), .o(n_6394) );
na02f80 g760927 ( .a(n_19499), .b(n_19498), .o(n_19500) );
no02f80 g755728 ( .a(n_25006), .b(n_24954), .o(n_25063) );
na02f80 g755696 ( .a(n_24484), .b(n_23282), .o(n_24553) );
oa12f80 g742859 ( .a(n_37135), .b(n_44039), .c(n_37082), .o(n_37188) );
in01f80 g770078 ( .a(n_10986), .o(n_10987) );
na02f80 g737567 ( .a(n_42428), .b(n_42371), .o(n_42429) );
in01f80 g753680 ( .a(n_26647), .o(n_26648) );
ao12f80 g778508 ( .a(n_2319), .b(n_2318), .c(n_2317), .o(n_3127) );
no02f80 g759544 ( .a(n_20843), .b(n_20791), .o(n_20881) );
na02f80 g780566 ( .a(n_679), .b(n_695), .o(n_882) );
na02f80 g776620 ( .a(n_4012), .b(n_3082), .o(n_4358) );
no02f80 g750654 ( .a(n_29373), .b(n_29372), .o(n_29374) );
in01f80 FE_RC_3862_0 ( .a(n_21736), .o(FE_RN_1687_0) );
in01f80 g743300 ( .a(n_36780), .o(n_36781) );
no02f80 g748000 ( .a(n_31814), .b(n_31667), .o(n_31908) );
na02f80 g773712 ( .a(n_7287), .b(n_7098), .o(n_7323) );
na02f80 g742079 ( .a(FE_OCP_RBN3445_n_37945), .b(n_38279), .o(n_38352) );
in01f80 g740108 ( .a(n_40279), .o(n_40280) );
ao12f80 g781273 ( .a(n_119), .b(n_7), .c(beta_26), .o(n_153) );
no02f80 g778987 ( .a(n_2093), .b(n_2092), .o(n_2094) );
no02f80 g739434 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .o(n_40723) );
na02f80 g746070 ( .a(n_33903), .b(n_33876), .o(n_33956) );
in01f80 g757405 ( .a(n_23097), .o(n_23098) );
in01f80 g754134 ( .a(n_26085), .o(n_26086) );
in01f80 g767595 ( .a(n_13052), .o(n_13053) );
in01f80 newInst_494 ( .a(newNet_313), .o(newNet_494) );
oa22f80 g784554 ( .a(FE_OFN800_n_46285), .b(n_11061), .c(FE_OCP_RBN3709_n_46337), .d(n_11036), .o(n_46375) );
in01f80 g774386 ( .a(n_6892), .o(n_6893) );
in01f80 newInst_1878 ( .a(newNet_1503), .o(newNet_1878) );
na02f80 g759041 ( .a(n_21318), .b(n_21317), .o(n_21356) );
oa12f80 g750308 ( .a(n_29657), .b(n_29648), .c(n_29702), .o(n_29719) );
oa12f80 g749640 ( .a(n_30266), .b(n_30283), .c(n_30265), .o(n_30322) );
in01f80 newInst_12 ( .a(newNet_9), .o(newNet_12) );
no02f80 g759007 ( .a(n_21495), .b(n_21533), .o(n_22038) );
na02f80 g781059 ( .a(sin_out_4), .b(FE_OFN4_n_43918), .o(n_318) );
in01f80 g744873 ( .a(n_35165), .o(n_36062) );
in01f80 newInst_2485 ( .a(newNet_2484), .o(newNet_2485) );
in01f80 g757543 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .o(n_22865) );
oa12f80 g768606 ( .a(n_12179), .b(n_12260), .c(n_12092), .o(n_12334) );
oa22f80 g752608 ( .a(n_28239), .b(n_28024), .c(n_28240), .d(n_28023), .o(n_28923) );
in01f80 newInst_3446 ( .a(newNet_3445), .o(newNet_3446) );
no02f80 g746387 ( .a(n_34778), .b(n_34815), .o(n_34868) );
in01f80 FE_OCP_RBC2452_n_38537 ( .a(n_38537), .o(FE_OCP_RBN2452_n_38537) );
in01f80 g767364 ( .a(n_13649), .o(n_13650) );
no02f80 g769607 ( .a(n_11367), .b(n_11269), .o(n_11413) );
na03f80 FE_RC_3989_0 ( .a(FE_RN_1729_0), .b(n_29815), .c(n_29903), .o(FE_RN_1730_0) );
in01f80 g741188 ( .a(n_39004), .o(n_38950) );
na02f80 g772365 ( .a(n_8677), .b(n_8676), .o(n_8771) );
no02f80 g751323 ( .a(n_28684), .b(n_28658), .o(n_28659) );
in01f80 g737599 ( .a(n_42465), .o(n_42466) );
in01f80 FE_OCPC1418_n_31504 ( .a(FE_OCPN1417_n_31504), .o(FE_OCPN1418_n_31504) );
na02f80 g745934 ( .a(n_34049), .b(FE_OCP_RBN2323_n_33942), .o(n_34079) );
in01f80 g755901 ( .a(n_24320), .o(n_24311) );
na02f80 g738192 ( .a(n_41993), .b(n_41992), .o(n_41994) );
in01f80 FE_OCP_RBC2667_n_4158 ( .a(n_4158), .o(FE_OCP_RBN2667_n_4158) );
in01f80 g768983 ( .a(n_12017), .o(n_12018) );
in01f80 g768850 ( .a(n_12221), .o(n_12222) );
in01f80 g739456 ( .a(n_40669), .o(n_40670) );
in01f80 newInst_2209 ( .a(newNet_571), .o(newNet_2209) );
na02f80 g764400 ( .a(n_16277), .b(n_16194), .o(n_16363) );
in01f80 g763916 ( .a(n_17098), .o(n_17263) );
in01f80 g755193 ( .a(n_25745), .o(n_26512) );
no02f80 g741400 ( .a(n_38785), .b(n_38771), .o(n_38806) );
no02f80 g759296 ( .a(n_21065), .b(n_45023), .o(n_21219) );
in01f80 g761642 ( .a(n_19794), .o(n_19571) );
no02f80 FE_RC_2450_0 ( .a(FE_RN_977_0), .b(FE_RN_979_0), .o(FE_RN_980_0) );
in01f80 g737932 ( .a(n_42556), .o(n_42557) );
na02f80 g772651 ( .a(n_8243), .b(FE_OCP_RBN2415_n_8219), .o(n_8284) );
na02f80 g766395 ( .a(n_14128), .b(n_14122), .o(n_14184) );
na02f80 g743218 ( .a(n_35473), .b(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .o(n_37032) );
na02f80 g763004 ( .a(n_17616), .b(n_17617), .o(n_17646) );
in01f80 g751521 ( .a(n_28820), .o(n_28821) );
in01f80 g740054 ( .a(n_40076), .o(n_40077) );
in01f80 g765357 ( .a(n_15256), .o(n_15257) );
na02f80 FE_RC_2891_0 ( .a(n_33880), .b(n_33925), .o(FE_RN_1252_0) );
na02f80 g739735 ( .a(n_40472), .b(n_40147), .o(n_40524) );
in01f80 newInst_69 ( .a(newNet_36), .o(newNet_69) );
no02f80 g736706 ( .a(n_43219), .b(n_43120), .o(n_43327) );
no02f80 g757810 ( .a(n_23027), .b(n_22655), .o(n_23089) );
na02f80 g757358 ( .a(n_23161), .b(n_23160), .o(n_23515) );
in01f80 FE_RC_3617_0 ( .a(n_45067), .o(FE_RN_1582_0) );
in01f80 newInst_3536 ( .a(newNet_3535), .o(newNet_3536) );
na02f80 g742907 ( .a(n_37133), .b(n_37010), .o(n_37464) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_1_ ( .ck(newNet_825), .d(n_1307), .o(delay_xor_ln21_unr3_stage2_stallmux_q_1_) );
no02f80 g776088 ( .a(n_4840), .b(n_4848), .o(n_4872) );
na02f80 g737883 ( .a(n_42270), .b(n_42570), .o(n_42657) );
in01f80 newInst_860 ( .a(newNet_859), .o(newNet_860) );
oa12f80 g765119 ( .a(n_15414), .b(n_15413), .c(n_15412), .o(n_15488) );
no02f80 g760513 ( .a(n_19892), .b(n_18553), .o(n_20004) );
oa22f80 FE_RC_3369_0 ( .a(FE_RN_795_0), .b(FE_RN_796_0), .c(FE_RN_797_0), .d(n_20820), .o(n_20849) );
oa12f80 g766141 ( .a(n_14510), .b(n_14467), .c(n_44850), .o(n_14600) );
in01f80 FE_OCP_RBC3126_n_27632 ( .a(n_27632), .o(FE_OCP_RBN3126_n_27632) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_16_ ( .ck(newNet_252), .d(n_46177), .o(delay_xor_ln22_unr6_stage3_stallmux_q_16_) );
in01f80 g752633 ( .a(n_27590), .o(n_27591) );
in01f80 newInst_3209 ( .a(newNet_3208), .o(newNet_3209) );
in01f80 FE_OCP_RBC3086_n_31819 ( .a(FE_OCP_RBN3084_n_31819), .o(FE_OCP_RBN3086_n_31819) );
no02f80 FE_RC_2960_0 ( .a(FE_RN_1292_0), .b(n_39816), .o(n_39872) );
in01f80 g778851 ( .a(n_2913), .o(n_3029) );
no02f80 g763817 ( .a(n_17153), .b(n_17308), .o(n_18083) );
in01f80 g745104 ( .a(n_34711), .o(n_34728) );
na02f80 g746291 ( .a(n_33657), .b(n_33636), .o(n_33706) );
na02f80 g759066 ( .a(n_21354), .b(n_21353), .o(n_21355) );
in01f80 FE_RC_3049_0 ( .a(FE_RN_1336_0), .o(n_26783) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_9_ ( .ck(newNet_895), .d(n_27894), .o(delay_xor_ln21_unr18_stage7_stallmux_q_9_) );
oa22f80 g743600 ( .a(n_36378), .b(n_36255), .c(n_36379), .d(n_36254), .o(n_36433) );
na02f80 g747822 ( .a(n_33226), .b(n_33279), .o(n_33293) );
in01f80 newInst_947 ( .a(newNet_349), .o(newNet_947) );
in01f80 newInst_3297 ( .a(newNet_1710), .o(newNet_3297) );
in01f80 FE_OCP_RBC3584_n_14681 ( .a(n_14681), .o(FE_OCP_RBN3584_n_14681) );
na02f80 g755580 ( .a(n_24534), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24535) );
oa12f80 g745953 ( .a(n_34699), .b(n_35299), .c(n_35070), .o(n_35338) );
ao12f80 g784607 ( .a(n_42996), .b(n_42985), .c(n_42708), .o(n_46935) );
na02f80 g736949 ( .a(n_43242), .b(n_43211), .o(n_43521) );
na02f80 g765925 ( .a(FE_OCP_RBN3595_n_14785), .b(n_14215), .o(n_14848) );
na02f80 g767781 ( .a(n_12823), .b(n_11886), .o(n_12824) );
ao12f80 g774902 ( .a(n_6198), .b(n_6235), .c(n_6234), .o(n_6261) );
in01f80 g738811 ( .a(n_41382), .o(n_41456) );
in01f80 g768540 ( .a(n_12352), .o(n_12330) );
in01f80 g753149 ( .a(n_27488), .o(n_27489) );
na02f80 g770324 ( .a(n_10570), .b(n_44463), .o(n_10591) );
no02f80 g746431 ( .a(n_33456), .b(n_33455), .o(n_33457) );
no02f80 g739234 ( .a(n_41010), .b(n_40785), .o(n_41165) );
in01f80 newInst_738 ( .a(newNet_737), .o(newNet_738) );
no02f80 g763468 ( .a(n_17129), .b(n_16973), .o(n_17247) );
in01f80 newInst_1842 ( .a(newNet_1841), .o(newNet_1842) );
no02f80 g759516 ( .a(n_20853), .b(n_20852), .o(n_20936) );
no02f80 g741204 ( .a(n_38870), .b(FE_OCP_RBN2370_n_38545), .o(n_39097) );
no02f80 g748290 ( .a(n_31591), .b(n_31610), .o(n_31611) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_22_ ( .ck(newNet_1990), .d(n_11731), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_) );
na02f80 g775633 ( .a(n_5192), .b(n_5152), .o(n_5232) );
na02f80 g749882 ( .a(n_29894), .b(n_29927), .o(n_29989) );
na02f80 FE_RC_2217_0 ( .a(n_32533), .b(FE_RN_800_0), .o(FE_RN_801_0) );
in01f80 newInst_3008 ( .a(newNet_3007), .o(newNet_3008) );
in01f80 newInst_1534 ( .a(newNet_977), .o(newNet_1534) );
in01f80 newInst_1463 ( .a(newNet_1200), .o(newNet_1463) );
no02f80 FE_RC_1953_0 ( .a(FE_RN_625_0), .b(FE_RN_628_0), .o(n_25940) );
in01f80 FE_RC_984_0 ( .a(FE_RN_284_0), .o(n_27675) );
na02f80 g745071 ( .a(n_34717), .b(n_34716), .o(n_34718) );
in01f80 g767767 ( .a(n_13369), .o(n_13370) );
oa22f80 FE_RC_3362_0 ( .a(n_31829), .b(n_32244), .c(n_31830), .d(n_32226), .o(n_32340) );
oa22f80 g777225 ( .a(n_3705), .b(n_3717), .c(n_3698), .d(n_3715), .o(n_3803) );
no02f80 g780385 ( .a(n_937), .b(n_860), .o(n_861) );
in01f80 g741316 ( .a(n_39131), .o(n_39129) );
oa12f80 g767317 ( .a(n_12809), .b(n_13336), .c(n_12731), .o(n_13409) );
no02f80 g742119 ( .a(n_38180), .b(n_38213), .o(n_38233) );
no02f80 g775136 ( .a(n_5787), .b(n_5769), .o(n_5907) );
na02f80 g749970 ( .a(n_30114), .b(n_30053), .o(n_30141) );
in01f80 g765049 ( .a(n_15496), .o(n_15608) );
in01f80 g752018 ( .a(n_29155), .o(n_29290) );
na02f80 g744286 ( .a(FE_OCP_RBN2902_n_44174), .b(FE_OCP_RBN2642_n_34921), .o(n_35776) );
no02f80 g755146 ( .a(n_25745), .b(n_26451), .o(n_25746) );
in01f80 g762110 ( .a(n_18462), .o(n_18424) );
in01f80 FE_RC_2262_0 ( .a(n_25081), .o(FE_RN_838_0) );
in01f80 newInst_552 ( .a(newNet_551), .o(newNet_552) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_7_ ( .ck(newNet_2704), .d(n_15842), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_) );
in01f80 g755148 ( .a(n_25071), .o(n_25072) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_18_ ( .ck(newNet_3062), .d(n_1001), .o(delay_add_ln22_unr2_stage2_stallmux_q_18_) );
in01f80 g739150 ( .a(n_40915), .o(n_40964) );
no02f80 g776554 ( .a(n_4307), .b(n_3297), .o(n_4308) );
na02f80 g775955 ( .a(n_4807), .b(n_4801), .o(n_4908) );
in01f80 FE_OCP_RBC3654_n_10100 ( .a(FE_OCP_RBN3652_n_10100), .o(FE_OCP_RBN3654_n_10100) );
in01f80 g767425 ( .a(n_13587), .o(n_13620) );
in01f80 g740796 ( .a(n_39384), .o(n_39385) );
in01f80 newInst_2606 ( .a(newNet_2605), .o(newNet_2606) );
oa12f80 g771698 ( .a(n_7554), .b(n_8863), .c(n_8840), .o(n_8864) );
in01f80 g769707 ( .a(n_11369), .o(n_11338) );
na02f80 g773092 ( .a(n_7811), .b(n_7921), .o(n_8468) );
no02f80 g755338 ( .a(n_24917), .b(n_24896), .o(n_24966) );
in01f80 g749032 ( .a(n_30947), .o(n_30948) );
no02f80 g774518 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .o(n_6765) );
no02f80 g769368 ( .a(FE_OCPN858_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n_12082) );
na02f80 g765274 ( .a(n_15116), .b(n_14340), .o(n_15117) );
na02f80 FE_RC_2962_0 ( .a(FE_OCP_RBN2523_n_8951), .b(n_9162), .o(FE_RN_1293_0) );
in01f80 g775861 ( .a(n_5230), .o(n_5231) );
na02f80 g774009 ( .a(n_6802), .b(n_6801), .o(n_6822) );
in01f80 g766993 ( .a(n_13582), .o(n_13583) );
na02f80 g769201 ( .a(n_12115), .b(n_12008), .o(n_12165) );
oa12f80 g751814 ( .a(n_28919), .b(n_29077), .c(n_29076), .o(n_29103) );
in01f80 g756098 ( .a(n_24981), .o(n_24994) );
in01f80 g773753 ( .a(n_7272), .o(n_7273) );
oa12f80 g749736 ( .a(n_31311), .b(n_31372), .c(n_31371), .o(n_31391) );
na02f80 g757188 ( .a(n_23214), .b(n_23213), .o(n_23300) );
no02f80 g744803 ( .a(n_35165), .b(FE_OCPN1794_n_30612), .o(n_35196) );
oa12f80 g772509 ( .a(n_8028), .b(n_8433), .c(n_7988), .o(n_8639) );
no02f80 g778295 ( .a(n_2517), .b(n_2443), .o(n_2709) );
oa12f80 g739083 ( .a(n_41033), .b(n_41051), .c(n_41032), .o(n_41438) );
in01f80 newInst_999 ( .a(newNet_998), .o(newNet_999) );
no02f80 g764726 ( .a(n_15741), .b(n_15767), .o(n_15951) );
in01f80 FE_OCP_RBC3041_n_46337 ( .a(n_46337), .o(FE_OCP_RBN3041_n_46337) );
in01f80 newInst_179 ( .a(newNet_153), .o(newNet_179) );
no02f80 g779347 ( .a(n_1623), .b(n_1622), .o(n_1653) );
na02f80 g774323 ( .a(n_6551), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6577) );
na02f80 g755296 ( .a(n_24968), .b(n_24745), .o(n_25010) );
na02f80 g760089 ( .a(FE_OCP_RBN1694_n_19052), .b(n_20300), .o(n_20342) );
in01f80 FE_OCP_RBC2383_n_8342 ( .a(n_8342), .o(FE_OCP_RBN2383_n_8342) );
oa12f80 g743631 ( .a(n_36205), .b(n_36410), .c(n_36270), .o(n_36482) );
in01f80 g771076 ( .a(n_10067), .o(n_10204) );
in01f80 g754918 ( .a(n_25389), .o(n_25422) );
na02f80 g738320 ( .a(n_41831), .b(n_41755), .o(n_41885) );
in01f80 newInst_1540 ( .a(newNet_622), .o(newNet_1540) );
ms00f80 sin_out_reg_23_ ( .ck(newNet_49), .d(n_43903), .o(sin_out_23) );
na02f80 g750149 ( .a(n_29869), .b(n_29211), .o(n_30071) );
na02f80 g769793 ( .a(n_11095), .b(n_11130), .o(n_11252) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_10_ ( .ck(newNet_1147), .d(n_10301), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_) );
in01f80 g748359 ( .a(n_33415), .o(n_33576) );
in01f80 newInst_749 ( .a(newNet_748), .o(newNet_749) );
no02f80 g766661 ( .a(n_13839), .b(n_13352), .o(n_13894) );
in01f80 newInst_2003 ( .a(newNet_2002), .o(newNet_2003) );
no02f80 g748319 ( .a(n_31594), .b(n_30871), .o(n_31606) );
in01f80 g738721 ( .a(n_41485), .o(n_41486) );
na02f80 g737918 ( .a(n_42270), .b(n_41952), .o(n_42558) );
ao12f80 g770194 ( .a(n_10556), .b(n_10745), .c(n_10603), .o(n_10821) );
no02f80 FE_RC_3947_0 ( .a(n_32835), .b(FE_RN_1707_0), .o(n_33168) );
in01f80 newInst_2468 ( .a(newNet_2467), .o(newNet_2468) );
na02f80 g745971 ( .a(n_33962), .b(n_33964), .o(n_33965) );
no02f80 g777693 ( .a(n_3447), .b(n_3369), .o(n_3468) );
na02f80 g769173 ( .a(n_11971), .b(n_11893), .o(n_12170) );
no02f80 g739514 ( .a(n_40685), .b(n_40684), .o(n_40808) );
in01f80 g753934 ( .a(n_26226), .o(n_26227) );
no02f80 FE_RC_2555_0 ( .a(FE_RN_1047_0), .b(n_37412), .o(n_37515) );
oa12f80 g744331 ( .a(n_35494), .b(n_35493), .c(n_35503), .o(n_35518) );
in01f80 g752386 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n_27778) );
no02f80 g759714 ( .a(FE_OCP_RBN3631_n_20504), .b(FE_OFN751_n_45003), .o(n_20589) );
in01f80 g738007 ( .a(n_42192), .o(n_42202) );
in01f80 g755438 ( .a(n_24756), .o(n_24757) );
in01f80 g770963 ( .a(n_9851), .o(n_9852) );
in01f80 newInst_3272 ( .a(newNet_3271), .o(newNet_3272) );
in01f80 g779300 ( .a(n_1733), .o(n_1734) );
no02f80 g742793 ( .a(n_37344), .b(n_37343), .o(n_37387) );
in01f80 newInst_1781 ( .a(newNet_1780), .o(newNet_1781) );
na02f80 g743135 ( .a(n_36986), .b(n_36985), .o(n_36987) );
na02f80 g774974 ( .a(n_6179), .b(n_6116), .o(n_6194) );
ao22s80 FE_RC_322_0 ( .a(FE_OCP_RBN1920_n_22476), .b(n_22502), .c(FE_OCP_RBN1921_n_22476), .d(FE_OCP_RBN3100_n_22502), .o(n_22622) );
in01f80 g743089 ( .a(n_37106), .o(n_37050) );
in01f80 FE_RC_3585_0 ( .a(FE_RN_1564_0), .o(FE_RN_1563_0) );
na02f80 g777070 ( .a(n_5329), .b(n_5328), .o(n_5333) );
ao12f80 g751435 ( .a(FE_OCP_RBN2216_FE_OCPN950_n_28595), .b(n_28773), .c(n_28795), .o(n_28804) );
na02f80 g777077 ( .a(n_3661), .b(n_3705), .o(n_3813) );
no02f80 g767008 ( .a(n_14419), .b(n_14207), .o(n_14486) );
na02f80 g740065 ( .a(n_40073), .b(n_40072), .o(n_40114) );
in01f80 fopt783262 ( .a(n_36410), .o(n_44831) );
no02f80 g768021 ( .a(n_12679), .b(n_12678), .o(n_12680) );
in01f80 g741801 ( .a(n_38562), .o(n_39393) );
no02f80 g750427 ( .a(n_29562), .b(FE_OCPN1406_n_25859), .o(n_29702) );
no02f80 g738576 ( .a(n_41614), .b(n_41613), .o(n_41615) );
no02f80 g756905 ( .a(n_23310), .b(n_23309), .o(n_23311) );
no02f80 g767016 ( .a(FE_OCP_RBN2503_n_13896), .b(n_14038), .o(n_14171) );
oa12f80 g741454 ( .a(n_38809), .b(n_38808), .c(n_38807), .o(n_39738) );
no02f80 g761764 ( .a(n_18517), .b(FE_OCP_RBN1166_n_18437), .o(n_18599) );
na02f80 g746733 ( .a(n_33144), .b(n_33099), .o(n_33190) );
na02f80 g779201 ( .a(n_1862), .b(n_1850), .o(n_1851) );
no02f80 g752806 ( .a(n_28297), .b(n_28257), .o(n_28379) );
in01f80 g769340 ( .a(n_11631), .o(n_11546) );
na02f80 g742396 ( .a(n_37765), .b(n_37764), .o(n_37766) );
in01f80 g760902 ( .a(n_19461), .o(n_19503) );
in01f80 g780593 ( .a(n_793), .o(n_794) );
no02f80 g754115 ( .a(n_26114), .b(n_26113), .o(n_26116) );
no02f80 g765382 ( .a(FE_OCP_RBN3620_n_15135), .b(n_14055), .o(n_15461) );
in01f80 newInst_2762 ( .a(newNet_2761), .o(newNet_2762) );
na02f80 g742500 ( .a(n_37563), .b(n_37561), .o(n_37562) );
na02f80 g752048 ( .a(n_28693), .b(n_28692), .o(n_28694) );
in01f80 newInst_3472 ( .a(newNet_3471), .o(newNet_3472) );
no02f80 g751341 ( .a(n_29511), .b(n_29510), .o(n_29512) );
no02f80 g736738 ( .a(n_43359), .b(n_43342), .o(n_43432) );
na02f80 g740918 ( .a(n_39286), .b(n_39285), .o(n_39287) );
in01f80 g746423 ( .a(n_34127), .o(n_33517) );
no02f80 g746709 ( .a(n_33083), .b(n_32998), .o(n_33112) );
no02f80 g749349 ( .a(n_30624), .b(n_30262), .o(n_30650) );
no02f80 g756243 ( .a(n_24737), .b(n_24736), .o(n_24738) );
no02f80 g777007 ( .a(n_3983), .b(n_3874), .o(n_4032) );
in01f80 FE_OCP_RBC2863_n_39523 ( .a(n_39523), .o(FE_OCP_RBN2863_n_39523) );
no02f80 g750434 ( .a(n_29577), .b(FE_OCP_DRV_N3741_n_29576), .o(n_29632) );
na02f80 g749921 ( .a(n_30077), .b(n_29327), .o(n_30119) );
na02f80 g780500 ( .a(n_869), .b(n_891), .o(n_930) );
in01f80 g773122 ( .a(n_7693), .o(n_7675) );
in01f80 FE_RC_4057_0 ( .a(n_26390), .o(FE_RN_1765_0) );
no02f80 g764242 ( .a(n_16376), .b(n_16405), .o(n_16445) );
in01f80 g774479 ( .a(n_6687), .o(n_6628) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_0_ ( .ck(newNet_373), .d(n_1314), .o(delay_xor_ln22_unr3_stage2_stallmux_q_0_) );
in01f80 FE_OCP_RBC3679_n_21051 ( .a(FE_OCP_RBN3678_n_21051), .o(FE_OCP_RBN3679_n_21051) );
no02f80 g763807 ( .a(n_17422), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n_17424) );
in01f80 newInst_756 ( .a(newNet_755), .o(newNet_756) );
in01f80 newInst_1557 ( .a(newNet_1556), .o(newNet_1557) );
in01f80 newInst_1000 ( .a(newNet_999), .o(newNet_1000) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_1_ ( .ck(newNet_2288), .d(n_39779), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_) );
in01f80 newInst_2504 ( .a(newNet_2503), .o(newNet_2504) );
oa22f80 g739935 ( .a(n_39961), .b(n_40322), .c(n_39962), .d(n_40323), .o(n_40410) );
oa22f80 g743661 ( .a(n_36391), .b(n_36359), .c(n_36390), .d(n_36360), .o(n_36440) );
na03f80 g784153 ( .a(n_1432), .b(n_1480), .c(n_1387), .o(n_45900) );
na02f80 g755709 ( .a(n_24326), .b(n_23886), .o(n_24408) );
na02f80 g744544 ( .a(n_35333), .b(n_35236), .o(n_35353) );
no02f80 g748792 ( .a(n_32445), .b(n_32459), .o(n_32556) );
in01f80 g769113 ( .a(n_11803), .o(n_11804) );
in01f80 newInst_3683 ( .a(newNet_2841), .o(newNet_3683) );
na02f80 g757900 ( .a(n_22884), .b(n_22783), .o(n_22954) );
in01f80 g769248 ( .a(n_11497), .o(n_11532) );
na02f80 g749365 ( .a(n_30672), .b(n_30671), .o(n_30673) );
in01f80 FE_OCP_RBC3605_n_8981 ( .a(FE_OCP_RBN3604_n_8981), .o(FE_OCP_RBN3605_n_8981) );
in01f80 FE_RC_126_0 ( .a(n_11993), .o(FE_RN_31_0) );
in01f80 FE_OCP_RBC3692_n_10852 ( .a(n_10852), .o(FE_OCP_RBN3692_n_10852) );
in01f80 newInst_342 ( .a(newNet_341), .o(newNet_342) );
in01f80 newInst_2107 ( .a(newNet_2106), .o(newNet_2107) );
in01f80 g773878 ( .a(n_7068), .o(n_7069) );
in01f80 g742255 ( .a(n_38266), .o(n_38267) );
na02f80 g776789 ( .a(n_4030), .b(n_3912), .o(n_4186) );
in01f80 g748775 ( .a(n_32587), .o(n_32532) );
in01f80 g777034 ( .a(n_3746), .o(n_3814) );
in01f80 g739955 ( .a(n_40409), .o(n_40436) );
na02f80 g777908 ( .a(n_3167), .b(n_3169), .o(n_3187) );
na02f80 g752348 ( .a(n_28457), .b(n_28445), .o(n_28446) );
in01f80 g776654 ( .a(n_4394), .o(n_4395) );
no02f80 g769076 ( .a(n_11436), .b(n_11458), .o(n_11604) );
in01f80 FE_OCPC847_n_3597 ( .a(n_3597), .o(FE_OCPN847_n_3597) );
na02f80 g764794 ( .a(n_15844), .b(n_15934), .o(n_16027) );
no02f80 g774347 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .o(n_6758) );
na02f80 g776252 ( .a(n_4792), .b(FE_OCP_RBN2578_n_47017), .o(n_4917) );
na02f80 g772604 ( .a(n_8390), .b(n_8389), .o(n_8484) );
in01f80 FE_OCP_RBC2656_FE_RN_1288_0 ( .a(FE_RN_1288_0), .o(FE_OCP_RBN2656_FE_RN_1288_0) );
in01f80 newInst_1768 ( .a(newNet_1767), .o(newNet_1768) );
in01f80 g739404 ( .a(n_40983), .o(n_40984) );
na02f80 g748036 ( .a(n_32107), .b(n_32024), .o(n_32108) );
no02f80 g745891 ( .a(n_35336), .b(n_34759), .o(n_35373) );
in01f80 g779463 ( .a(n_1773), .o(n_1774) );
in01f80 g777058 ( .a(n_3753), .o(n_3754) );
na02f80 g770887 ( .a(n_10013), .b(n_9820), .o(n_10071) );
in01f80 g756465 ( .a(n_23848), .o(n_23849) );
no02f80 g756896 ( .a(n_23384), .b(n_23095), .o(n_23387) );
no02f80 g764154 ( .a(n_16533), .b(n_16332), .o(n_16534) );
in01f80 FE_RC_3603_0 ( .a(FE_RN_1575_0), .o(n_20760) );
oa22f80 g757877 ( .a(n_22168), .b(n_22095), .c(n_22204), .d(n_22094), .o(n_22392) );
in01f80 FE_OCP_RBC2629_n_14590 ( .a(FE_OCP_RBN2628_n_14590), .o(FE_OCP_RBN2629_n_14590) );
na02f80 g748929 ( .a(n_31132), .b(n_31050), .o(n_31241) );
in01f80 FE_RC_1311_0 ( .a(n_3744), .o(FE_RN_385_0) );
in01f80 g744381 ( .a(n_46211), .o(n_36859) );
in01f80 FE_OCPC1398_n_21973 ( .a(FE_OCPN1397_n_21973), .o(FE_OCPN1398_n_21973) );
no02f80 g743768 ( .a(n_36074), .b(n_36075), .o(n_36110) );
in01f80 g739644 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_29_), .o(n_40891) );
oa12f80 g764343 ( .a(n_16181), .b(n_16366), .c(n_16271), .o(n_16394) );
na02f80 g751368 ( .a(n_28770), .b(n_28631), .o(n_28746) );
na02f80 g749424 ( .a(n_30515), .b(n_30502), .o(n_30580) );
na02f80 g742365 ( .a(n_37838), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37783) );
no02f80 g759509 ( .a(n_20650), .b(n_45010), .o(n_20774) );
in01f80 g772280 ( .a(n_8621), .o(n_8611) );
na02f80 g761867 ( .a(n_18368), .b(n_18367), .o(n_18406) );
na02f80 g764781 ( .a(n_15734), .b(n_14419), .o(n_15800) );
ao22s80 FE_RC_1980_0 ( .a(FE_RN_642_0), .b(n_19799), .c(FE_RN_643_0), .d(n_19722), .o(n_19915) );
na02f80 g742008 ( .a(n_38073), .b(n_37906), .o(n_38071) );
ao12f80 g780332 ( .a(n_879), .b(n_937), .c(n_878), .o(n_957) );
na02f80 g779061 ( .a(n_2085), .b(n_2084), .o(n_2518) );
na02f80 g751442 ( .a(n_28509), .b(n_28508), .o(n_28526) );
no02f80 g784758 ( .a(n_8889), .b(n_47235), .o(n_47244) );
in01f80 g779482 ( .a(n_1717), .o(n_1718) );
in01f80 g738188 ( .a(n_42006), .o(n_42007) );
in01f80 g773057 ( .a(n_7754), .o(n_7796) );
ao12f80 g757410 ( .a(n_23391), .b(n_44068), .c(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .o(n_23095) );
in01f80 g755564 ( .a(n_24717), .o(n_24794) );
in01f80 g746331 ( .a(n_33594), .o(n_33581) );
no02f80 g758042 ( .a(n_22690), .b(n_22729), .o(n_22763) );
in01f80 fopt783524 ( .a(n_45136), .o(n_45135) );
in01f80 g759956 ( .a(n_20251), .o(n_20271) );
in01f80 g752109 ( .a(n_28781), .o(n_28793) );
no02f80 g770984 ( .a(n_9582), .b(n_9461), .o(n_9581) );
no02f80 g772575 ( .a(n_8335), .b(FE_OCP_RBN3463_n_7886), .o(n_8398) );
no02f80 g776778 ( .a(n_4126), .b(n_3909), .o(n_4179) );
no02f80 g737506 ( .a(n_42535), .b(n_42534), .o(n_42536) );
in01f80 newInst_169 ( .a(newNet_168), .o(newNet_169) );
in01f80 g766841 ( .a(n_13601), .o(n_13631) );
no02f80 g764786 ( .a(n_15734), .b(n_14419), .o(n_15735) );
in01f80 g742172 ( .a(n_38307), .o(n_38308) );
in01f80 g756838 ( .a(n_23836), .o(n_23837) );
in01f80 g771101 ( .a(n_9637), .o(n_9713) );
in01f80 FE_OCP_RBC3130_n_17591 ( .a(n_17591), .o(FE_OCP_RBN3130_n_17591) );
oa22f80 FE_RC_3361_0 ( .a(FE_RN_699_0), .b(n_35078), .c(FE_RN_700_0), .d(FE_RN_701_0), .o(n_35198) );
in01f80 g740769 ( .a(n_39386), .o(n_39497) );
na02f80 g756044 ( .a(n_25032), .b(n_25027), .o(n_25081) );
na02f80 g774720 ( .a(n_6271), .b(n_6277), .o(n_6376) );
na02f80 g747825 ( .a(n_33392), .b(n_33437), .o(n_33495) );
in01f80 FE_OCP_RBC1378_n_20889 ( .a(FE_OCP_RBN1377_n_20889), .o(FE_OCP_RBN1378_n_20889) );
in01f80 newInst_1369 ( .a(newNet_1368), .o(newNet_1369) );
in01f80 g748095 ( .a(n_31853), .o(n_31876) );
no02f80 g751162 ( .a(n_29944), .b(n_29993), .o(n_30096) );
in01f80 FE_RC_2278_0 ( .a(n_28175), .o(FE_RN_850_0) );
na02f80 g740006 ( .a(n_40068), .b(n_40003), .o(n_40150) );
in01f80 g745563 ( .a(n_34745), .o(n_34746) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_6_ ( .ck(newNet_1069), .d(n_9917), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_) );
in01f80 g775232 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_19_), .o(n_5984) );
na02f80 g764293 ( .a(n_16278), .b(FE_OCPN3775_n_14730), .o(n_16377) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_9_ ( .ck(newNet_534), .d(n_17552), .o(delay_xor_ln22_unr12_stage5_stallmux_q_9_) );
oa12f80 g780340 ( .a(n_915), .b(n_955), .c(n_580), .o(n_1023) );
no02f80 FE_RC_2206_0 ( .a(FE_OCPN3186_FE_OCP_RBN1140_n_25816), .b(n_27120), .o(FE_RN_793_0) );
in01f80 FE_OCP_RBC3627_n_38870 ( .a(FE_OCP_RBN3625_n_38870), .o(FE_OCP_RBN3627_n_38870) );
na02f80 g736876 ( .a(n_43187), .b(n_43502), .o(n_43605) );
in01f80 g760796 ( .a(n_19621), .o(n_19622) );
ao22s80 FE_RC_931_0 ( .a(n_27246), .b(FE_OCP_RBN2911_n_30908), .c(n_27366), .d(n_30908), .o(n_31023) );
in01f80 g752680 ( .a(n_27532), .o(n_27533) );
in01f80 newInst_2385 ( .a(newNet_2384), .o(newNet_2385) );
no02f80 g744054 ( .a(n_44223), .b(n_34751), .o(n_35827) );
in01f80 newInst_409 ( .a(newNet_408), .o(newNet_409) );
na02f80 g766229 ( .a(n_14335), .b(n_14152), .o(n_14414) );
na02f80 g751911 ( .a(n_28988), .b(n_28987), .o(n_28989) );
in01f80 FE_RC_2700_0 ( .a(n_8303), .o(FE_RN_1133_0) );
in01f80 FE_OCP_RBC2734_n_4219 ( .a(FE_OCP_RBN2732_n_4219), .o(FE_OCP_RBN2734_n_4219) );
in01f80 g766487 ( .a(n_14093), .o(n_14094) );
no02f80 g774881 ( .a(n_6145), .b(n_6158), .o(n_6328) );
no02f80 g780758 ( .a(n_547), .b(n_543), .o(n_544) );
in01f80 g759360 ( .a(n_21754), .o(n_21755) );
ao22s80 FE_RC_4257_0 ( .a(FE_RN_1873_0), .b(n_22187), .c(FE_RN_1874_0), .d(n_22288), .o(n_22470) );
oa12f80 g738159 ( .a(n_42000), .b(n_41999), .c(n_41998), .o(n_42035) );
in01f80 newInst_2177 ( .a(newNet_2176), .o(newNet_2177) );
in01f80 g770256 ( .a(n_10848), .o(n_10814) );
no02f80 g749691 ( .a(n_31455), .b(n_31454), .o(n_31482) );
ao12f80 g747289 ( .a(n_32751), .b(n_32770), .c(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n_32811) );
oa12f80 g761364 ( .a(n_19826), .b(n_19980), .c(n_19793), .o(n_20515) );
in01f80 FE_OCP_RBC2358_n_13818 ( .a(n_13818), .o(FE_OCP_RBN2358_n_13818) );
na02f80 g753301 ( .a(n_27120), .b(FE_OCPN3797_n_26115), .o(n_27355) );
in01f80 newInst_291 ( .a(newNet_290), .o(newNet_291) );
no02f80 g771353 ( .a(n_9208), .b(n_9163), .o(n_9353) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_12_ ( .ck(newNet_1650), .d(n_27015), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_) );
in01f80 FE_OCP_RBC3044_n_46337 ( .a(FE_OCP_RBN3041_n_46337), .o(FE_OCP_RBN3044_n_46337) );
in01f80 g776421 ( .a(n_4494), .o(n_4495) );
no02f80 g774589 ( .a(n_6371), .b(n_5754), .o(n_6385) );
no02f80 g762023 ( .a(n_18205), .b(n_16990), .o(n_18285) );
na02f80 g747382 ( .a(n_32630), .b(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n_32810) );
in01f80 g774163 ( .a(n_7515), .o(n_6859) );
ao22s80 g777255 ( .a(n_47018), .b(n_3029), .c(FE_OCP_RBN2532_n_47018), .d(n_2913), .o(n_3689) );
in01f80 g762821 ( .a(n_17758), .o(n_17894) );
na02f80 g746238 ( .a(n_33706), .b(n_33768), .o(n_33820) );
na02f80 g750508 ( .a(n_29527), .b(FE_OFN788_n_25834), .o(n_29528) );
in01f80 g779001 ( .a(n_2181), .o(n_2182) );
oa22f80 g740124 ( .a(FE_OCP_RBN3055_n_39913), .b(n_39840), .c(FE_OCP_RBN3721_n_39913), .d(n_39460), .o(n_40318) );
in01f80 newInst_1716 ( .a(newNet_1715), .o(newNet_1716) );
ao12f80 g781257 ( .a(n_122), .b(n_7), .c(beta_18), .o(n_232) );
in01f80 FE_OCP_RBC2552_n_44921 ( .a(n_44921), .o(FE_OCP_RBN2552_n_44921) );
in01f80 newInst_2589 ( .a(newNet_2588), .o(newNet_2589) );
na02f80 g746812 ( .a(n_33377), .b(n_33376), .o(n_33402) );
no02f80 g743277 ( .a(n_37959), .b(n_37958), .o(n_37960) );
oa12f80 g767298 ( .a(n_13500), .b(n_13468), .c(n_13451), .o(n_13612) );
no02f80 g754490 ( .a(n_25518), .b(n_25517), .o(n_25519) );
na02f80 g748111 ( .a(n_31549), .b(n_31563), .o(n_31667) );
na02f80 FE_RC_2061_0 ( .a(n_23590), .b(FE_RN_698_0), .o(n_26797) );
na02f80 g743932 ( .a(n_35981), .b(n_44222), .o(n_36038) );
in01f80 newInst_2954 ( .a(newNet_2953), .o(newNet_2954) );
in01f80 g751733 ( .a(n_28355), .o(n_28356) );
na02f80 g763540 ( .a(n_16763), .b(n_16792), .o(n_16916) );
in01f80 g764087 ( .a(FE_OCP_RBN3358_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17256) );
in01f80 g740948 ( .a(n_39088), .o(n_39114) );
in01f80 g749590 ( .a(n_30405), .o(n_30424) );
na02f80 g752570 ( .a(n_27634), .b(n_27429), .o(n_27646) );
in01f80 g741221 ( .a(n_39322), .o(n_39323) );
na02f80 g746151 ( .a(n_33665), .b(n_33676), .o(n_33735) );
na02f80 g757391 ( .a(n_46964), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_), .o(n_23186) );
oa12f80 g764123 ( .a(n_16065), .b(n_16852), .c(n_16021), .o(n_16928) );
na02f80 g761492 ( .a(n_19787), .b(n_19399), .o(n_19930) );
na03f80 FE_RC_3971_0 ( .a(n_24345), .b(n_24411), .c(FE_OCP_RBN1060_n_24473), .o(n_24578) );
ao12f80 g748054 ( .a(n_31499), .b(n_31614), .c(n_31521), .o(n_31708) );
in01f80 newInst_1213 ( .a(newNet_1015), .o(newNet_1213) );
in01f80 g741151 ( .a(n_39203), .o(n_39204) );
in01f80 FE_OCPC866_n_45697 ( .a(FE_OCP_RBN2115_n_45224), .o(FE_OCPN866_n_45697) );
na02f80 g780559 ( .a(n_679), .b(n_678), .o(n_698) );
no02f80 FE_RC_711_0 ( .a(FE_RN_225_0), .b(FE_RN_226_0), .o(FE_RN_227_0) );
in01f80 g771179 ( .a(n_9822), .o(n_9924) );
in01f80 g760702 ( .a(n_19739), .o(n_19740) );
na02f80 g775509 ( .a(n_5755), .b(n_5697), .o(n_5698) );
ao12f80 g763211 ( .a(n_17272), .b(n_17472), .c(n_17393), .o(n_17433) );
in01f80 newInst_1498 ( .a(newNet_1497), .o(newNet_1498) );
in01f80 newInst_1796 ( .a(newNet_1795), .o(newNet_1796) );
oa22f80 g757860 ( .a(n_22237), .b(n_22183), .c(n_22316), .d(n_22184), .o(n_22479) );
oa12f80 g748566 ( .a(n_32657), .b(n_32658), .c(n_32656), .o(n_33370) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_30_ ( .ck(newNet_3201), .d(n_36669), .o(delay_add_ln22_unr23_stage9_stallmux_q_30_) );
in01f80 g758583 ( .a(n_22064), .o(n_22145) );
no02f80 g749844 ( .a(FE_OCP_RBN3013_n_31117), .b(n_31116), .o(n_31143) );
in01f80 g738069 ( .a(n_42130), .o(n_42131) );
in01f80 FE_OCP_RBC3478_n_13756 ( .a(n_13756), .o(FE_OCP_RBN3478_n_13756) );
no02f80 g767904 ( .a(FE_OCPN3757_n_13889), .b(n_12724), .o(n_12725) );
oa12f80 g751070 ( .a(n_30065), .b(n_30156), .c(n_29992), .o(n_30689) );
in01f80 fopt783427 ( .a(n_45024), .o(n_45023) );
no02f80 g746900 ( .a(FE_OCP_RBN3384_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_25_), .o(n_33264) );
in01f80 g749319 ( .a(n_30652), .o(n_30653) );
na02f80 g752179 ( .a(FE_OCPN878_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .o(n_28360) );
in01f80 g769850 ( .a(n_11278), .o(n_11232) );
oa22f80 FE_RC_72_0 ( .a(n_18238), .b(n_18475), .c(n_18239), .d(n_18476), .o(n_18678) );
in01f80 newInst_833 ( .a(newNet_832), .o(newNet_833) );
na02f80 g738144 ( .a(n_42066), .b(n_42065), .o(n_42064) );
oa22f80 g747642 ( .a(n_32143), .b(n_31834), .c(n_32144), .d(n_31833), .o(n_32255) );
no03m80 FE_RC_1074_0 ( .a(n_1543), .b(n_1422), .c(n_1521), .o(n_1557) );
in01f80 newInst_2419 ( .a(newNet_2418), .o(newNet_2419) );
na02f80 g755419 ( .a(n_24662), .b(n_24698), .o(n_24760) );
no02f80 g740936 ( .a(n_39194), .b(n_38937), .o(n_39261) );
na02f80 g758009 ( .a(n_22261), .b(n_22300), .o(n_22340) );
na02f80 g747126 ( .a(n_32953), .b(n_32952), .o(n_33007) );
na03f80 g746451 ( .a(n_33276), .b(n_33275), .c(n_32895), .o(n_33346) );
no02f80 g771188 ( .a(n_9195), .b(n_9145), .o(n_9359) );
in01f80 FE_RC_3988_0 ( .a(n_29832), .o(FE_RN_1729_0) );
ao12f80 g777390 ( .a(n_3467), .b(n_3466), .c(n_3465), .o(n_5166) );
no02f80 g760045 ( .a(n_20162), .b(n_20216), .o(n_20250) );
no02f80 FE_RC_2644_0 ( .a(n_23172), .b(n_23173), .o(FE_RN_1103_0) );
in01f80 newInst_1959 ( .a(newNet_1039), .o(newNet_1959) );
na02f80 g777753 ( .a(n_3392), .b(n_3376), .o(n_3503) );
na02f80 g767800 ( .a(n_13315), .b(n_13167), .o(n_13316) );
in01f80 g780554 ( .a(n_845), .o(n_736) );
in01f80 FE_RC_2047_0 ( .a(n_25626), .o(FE_RN_689_0) );
in01f80 newInst_3395 ( .a(newNet_1906), .o(newNet_3395) );
in01f80 newInst_2538 ( .a(newNet_1524), .o(newNet_2538) );
no02f80 g745307 ( .a(n_35581), .b(n_35187), .o(n_35606) );
in01f80 FE_OCP_RBC2207_n_12907 ( .a(FE_OCP_RBN2206_n_12907), .o(FE_OCP_RBN2207_n_12907) );
in01f80 g738471 ( .a(n_41414), .o(n_41428) );
na02f80 g751213 ( .a(n_29783), .b(n_29769), .o(n_29770) );
na02f80 g780522 ( .a(n_771), .b(n_747), .o(n_1145) );
na02f80 g766799 ( .a(n_13827), .b(n_13800), .o(n_13801) );
na02f80 g760789 ( .a(n_19563), .b(FE_OCP_DRV_N1562_n_19562), .o(n_19656) );
no02f80 g779291 ( .a(n_1712), .b(n_1711), .o(n_1713) );
na02f80 g765639 ( .a(n_15324), .b(n_14424), .o(n_15366) );
na02f80 g744087 ( .a(n_35595), .b(FE_OCP_DRV_N1586_n_35594), .o(n_35650) );
in01f80 newInst_1604 ( .a(newNet_1603), .o(newNet_1604) );
no02f80 g775465 ( .a(n_5441), .b(n_5340), .o(n_5503) );
na02f80 g776981 ( .a(n_4035), .b(n_4034), .o(n_4087) );
ao12f80 g780637 ( .a(n_745), .b(n_809), .c(n_808), .o(n_768) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_5_ ( .ck(newNet_1685), .d(n_21932), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_) );
no02f80 g761032 ( .a(n_19992), .b(n_20010), .o(n_20896) );
oa12f80 g772909 ( .a(n_7898), .b(n_7897), .c(n_7896), .o(n_7978) );
in01f80 g773371 ( .a(n_7721), .o(n_7743) );
na02f80 g778538 ( .a(n_2438), .b(n_3084), .o(n_2548) );
in01f80 newInst_1653 ( .a(newNet_1652), .o(newNet_1653) );
in01f80 newInst_3627 ( .a(newNet_3626), .o(newNet_3627) );
no03m80 FE_RC_2434_0 ( .a(n_6749), .b(FE_RN_969_0), .c(n_7332), .o(n_47176) );
in01f80 FE_OCP_RBC1347_n_19270 ( .a(FE_OCP_RBN1346_n_19270), .o(FE_OCP_RBN1347_n_19270) );
oa12f80 g749720 ( .a(n_31175), .b(n_31174), .c(n_186), .o(n_31226) );
na02f80 g758054 ( .a(n_22783), .b(n_22620), .o(n_22784) );
ao12f80 g747946 ( .a(n_33093), .b(n_33092), .c(n_33091), .o(n_33683) );
in01f80 g744796 ( .a(n_35204), .o(n_35172) );
in01f80 newInst_2140 ( .a(newNet_2139), .o(newNet_2140) );
in01f80 g776816 ( .a(n_4152), .o(n_4190) );
oa12f80 g760249 ( .a(n_20896), .b(n_20834), .c(n_20040), .o(n_21050) );
in01f80 g760183 ( .a(n_20703), .o(n_20704) );
in01f80 newInst_2692 ( .a(newNet_2691), .o(newNet_2692) );
na02f80 g746414 ( .a(n_33331), .b(n_33038), .o(n_33409) );
no02f80 g739359 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_22_), .o(n_40908) );
in01f80 newInst_3098 ( .a(newNet_3097), .o(newNet_3098) );
in01f80 g763571 ( .a(n_17128), .o(n_17061) );
no02f80 g775114 ( .a(n_5831), .b(n_5885), .o(n_5946) );
in01f80 g755466 ( .a(n_24857), .o(n_24872) );
na02f80 g780409 ( .a(n_935), .b(n_784), .o(n_1155) );
in01f80 newInst_1927 ( .a(newNet_493), .o(newNet_1927) );
na02f80 g753866 ( .a(n_26226), .b(FE_OCP_RBN1203_n_26121), .o(n_26304) );
in01f80 newInst_687 ( .a(newNet_686), .o(newNet_687) );
in01f80 FE_OCP_RBC3520_n_19663 ( .a(n_19663), .o(FE_OCP_RBN3520_n_19663) );
in01f80 g773014 ( .a(n_7756), .o(n_7784) );
na02f80 g748346 ( .a(n_31759), .b(n_31725), .o(n_31829) );
in01f80 newInst_2570 ( .a(newNet_2569), .o(newNet_2570) );
no02f80 g762624 ( .a(FE_OCP_RBN2142_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .o(n_18051) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_28_ ( .ck(newNet_1086), .d(n_11402), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_) );
no02f80 g765287 ( .a(n_15967), .b(n_15868), .o(n_15968) );
no02f80 g760390 ( .a(n_20701), .b(n_20700), .o(n_20702) );
in01f80 g748618 ( .a(n_31646), .o(n_31647) );
in01f80 g737087 ( .a(n_43013), .o(n_43017) );
ao12f80 g775847 ( .a(n_4962), .b(n_5283), .c(n_5017), .o(n_5332) );
in01f80 FE_OCP_DRV_C1548_n_17643 ( .a(FE_OCP_DRV_N1547_n_17643), .o(FE_OCP_DRV_N1548_n_17643) );
in01f80 g765487 ( .a(n_16173), .o(n_16174) );
na02f80 g740666 ( .a(n_39587), .b(n_39601), .o(n_40011) );
na02f80 g767979 ( .a(n_13162), .b(n_12993), .o(n_13733) );
no02f80 g748131 ( .a(n_32782), .b(n_32418), .o(n_32809) );
oa22f80 FE_RC_1173_0 ( .a(n_7514), .b(n_8476), .c(n_8461), .d(n_7513), .o(n_8599) );
na02f80 g761020 ( .a(n_19178), .b(n_18459), .o(n_19215) );
na02f80 g768387 ( .a(n_12463), .b(n_12462), .o(n_12506) );
in01f80 g773614 ( .a(n_7395), .o(n_7396) );
in01f80 g747557 ( .a(n_32310), .o(n_32285) );
in01f80 g760344 ( .a(n_20871), .o(n_21595) );
in01f80 g778029 ( .a(n_3047), .o(n_3048) );
in01f80 g754593 ( .a(n_26924), .o(n_26925) );
in01f80 FE_OCP_RBC2550_n_44944 ( .a(FE_OCP_RBN2545_n_44944), .o(FE_OCP_RBN2550_n_44944) );
no02f80 g745654 ( .a(n_34308), .b(n_34366), .o(n_34450) );
na03f80 FE_RC_3764_0 ( .a(n_24231), .b(n_24319), .c(n_24320), .o(n_24347) );
no02f80 g761463 ( .a(n_19647), .b(n_19794), .o(n_20234) );
in01f80 g739034 ( .a(n_41098), .o(n_41114) );
in01f80 g756567 ( .a(n_23711), .o(n_23712) );
no02f80 g770135 ( .a(n_11502), .b(n_44463), .o(n_10729) );
no02f80 g741962 ( .a(n_38164), .b(n_38131), .o(n_38165) );
no02f80 g776865 ( .a(n_3723), .b(n_2849), .o(n_3812) );
no02f80 g748143 ( .a(n_47271), .b(n_31967), .o(n_31990) );
in01f80 g748013 ( .a(n_32060), .o(n_32079) );
na02f80 g744253 ( .a(n_44180), .b(n_34893), .o(n_36138) );
na02f80 g779391 ( .a(n_1551), .b(n_1393), .o(n_1552) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_1_ ( .ck(newNet_3625), .d(n_15033), .o(delay_add_ln22_unr11_stage5_stallmux_q_1_) );
in01f80 g736836 ( .a(n_43258), .o(n_43259) );
in01f80 g761107 ( .a(n_19177), .o(n_19204) );
in01f80 g736796 ( .a(n_43145), .o(n_43146) );
na02f80 g757809 ( .a(n_23027), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_7_), .o(n_23028) );
no02f80 g771003 ( .a(n_9796), .b(n_8388), .o(n_9891) );
no02f80 g770462 ( .a(n_10437), .b(n_44490), .o(n_10508) );
oa22f80 FE_RC_1551_0 ( .a(n_45508), .b(n_40627), .c(FE_OCP_RBN2133_n_45508), .d(n_40628), .o(n_40676) );
in01f80 g752140 ( .a(n_28179), .o(n_28180) );
na02f80 g780843 ( .a(n_561), .b(n_570), .o(n_571) );
ao22s80 FE_RC_3778_0 ( .a(n_19686), .b(n_19964), .c(n_19687), .d(n_19963), .o(n_20072) );
in01f80 g773581 ( .a(n_7437), .o(n_7438) );
in01f80 FE_RC_3664_0 ( .a(FE_RN_1609_0), .o(n_26532) );
no02f80 g766598 ( .a(n_13890), .b(FE_OFN747_n_13889), .o(n_13922) );
in01f80 FE_OCP_RBC2871_n_39542 ( .a(n_39542), .o(FE_OCP_RBN2871_n_39542) );
na02f80 g760678 ( .a(n_19691), .b(FE_OCP_RBN1699_n_19353), .o(n_19745) );
in01f80 g770800 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_4_), .o(n_12127) );
ms00f80 sin_out_reg_4_ ( .ck(newNet_25), .d(n_43685), .o(sin_out_4) );
in01f80 FE_OCP_RBC2381_n_3502 ( .a(n_3502), .o(FE_OCP_RBN2381_n_3502) );
oa12f80 g744975 ( .a(n_35795), .b(n_36386), .c(n_35807), .o(n_36403) );
na02f80 g737368 ( .a(n_42837), .b(n_42828), .o(n_42956) );
in01f80 g743123 ( .a(n_37040), .o(n_37041) );
na02f80 g773233 ( .a(n_7709), .b(n_7691), .o(n_7744) );
no02f80 g739114 ( .a(n_41030), .b(n_40780), .o(n_41058) );
na02f80 g736848 ( .a(n_43461), .b(n_43149), .o(n_43549) );
in01f80 newInst_2313 ( .a(newNet_850), .o(newNet_2313) );
in01f80 g778945 ( .a(n_2300), .o(n_2301) );
in01f80 g775212 ( .a(n_5790), .o(n_5852) );
no02f80 g780922 ( .a(n_457), .b(n_516), .o(n_542) );
na02f80 g765318 ( .a(n_15156), .b(FE_OCP_RBN3509_n_13860), .o(n_15272) );
no02f80 g752504 ( .a(n_27712), .b(n_27710), .o(n_27713) );
oa22f80 FE_RC_1227_0 ( .a(n_8940), .b(n_7597), .c(n_7596), .d(n_8939), .o(n_9082) );
in01f80 g747697 ( .a(n_33394), .o(n_33374) );
oa22f80 g784539 ( .a(n_11856), .b(FE_OFN803_n_46285), .c(n_11805), .d(FE_OCP_RBN3043_n_46337), .o(n_46360) );
oa22f80 g776274 ( .a(n_4271), .b(n_4226), .c(n_4272), .d(n_4227), .o(n_4459) );
in01f80 newInst_2340 ( .a(newNet_2339), .o(newNet_2340) );
na02f80 g743019 ( .a(n_37082), .b(n_36625), .o(n_37069) );
in01f80 g765219 ( .a(n_16256), .o(n_16257) );
in01f80 FE_RC_437_0 ( .a(n_17326), .o(FE_RN_123_0) );
in01f80 g769003 ( .a(n_11829), .o(n_11830) );
in01f80 g759109 ( .a(n_21351), .o(n_21352) );
no02f80 g752786 ( .a(n_27990), .b(n_27878), .o(n_27904) );
no02f80 g757218 ( .a(n_23530), .b(n_23529), .o(n_23531) );
in01f80 g754573 ( .a(n_26769), .o(n_26814) );
no02f80 g770286 ( .a(n_10781), .b(FE_OCP_RBN2718_n_9182), .o(n_10805) );
no02f80 g755168 ( .a(n_25714), .b(n_25689), .o(n_25690) );
no02f80 FE_RC_2229_0 ( .a(FE_RN_809_0), .b(FE_RN_810_0), .o(FE_RN_811_0) );
na02f80 g764421 ( .a(n_16169), .b(n_14650), .o(n_16200) );
in01f80 g766334 ( .a(n_14366), .o(n_14367) );
na02f80 g763426 ( .a(n_16986), .b(n_16943), .o(n_17176) );
na02f80 g760874 ( .a(FE_OCP_RBN3841_n_19419), .b(n_19508), .o(n_19510) );
no02f80 g763456 ( .a(n_17165), .b(n_17117), .o(n_17313) );
na02f80 g765933 ( .a(n_14811), .b(n_14845), .o(n_14846) );
in01f80 g753017 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n_27721) );
in01f80 g760548 ( .a(n_20077), .o(n_19994) );
na02f80 g760133 ( .a(n_20456), .b(FE_OCP_RBN2427_n_19599), .o(n_20708) );
na02f80 FE_RC_4259_0 ( .a(FE_RN_1875_0), .b(n_22596), .o(FE_RN_1876_0) );
no03m80 FE_RC_664_0 ( .a(n_38034), .b(n_38011), .c(n_38124), .o(n_38172) );
na02f80 g758065 ( .a(n_22654), .b(n_22648), .o(n_23154) );
no02f80 g747686 ( .a(n_32265), .b(n_32106), .o(n_32324) );
na02f80 g749466 ( .a(n_30468), .b(n_30280), .o(n_30513) );
ao12f80 g738866 ( .a(n_41262), .b(n_41261), .c(n_41260), .o(n_41296) );
in01f80 g746224 ( .a(n_33771), .o(n_33803) );
ao12f80 g756634 ( .a(n_24191), .b(n_24190), .c(n_24189), .o(n_24275) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_1_ ( .ck(newNet_1912), .d(n_36741), .o(delay_sub_ln22_unr24_stage9_stallmux_q_1_) );
in01f80 g760980 ( .a(n_19380), .o(n_19381) );
no02f80 g769924 ( .a(n_10910), .b(n_10802), .o(n_10936) );
ao12f80 g775644 ( .a(n_5406), .b(n_5455), .c(n_5405), .o(n_5538) );
in01f80 g753318 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .o(n_26972) );
no02f80 g740721 ( .a(n_39416), .b(n_39415), .o(n_39417) );
in01f80 g780240 ( .a(n_1041), .o(n_1042) );
oa22f80 FE_RC_3234_0 ( .a(n_11742), .b(n_12022), .c(n_11741), .d(n_11986), .o(n_12217) );
oa22f80 FE_RC_1586_0 ( .a(n_17584), .b(n_17835), .c(n_16339), .d(n_47195), .o(n_17880) );
oa12f80 g743284 ( .a(n_46228), .b(n_37899), .c(n_46227), .o(n_37992) );
na02f80 g773850 ( .a(n_7111), .b(n_7110), .o(n_7112) );
oa12f80 g736450 ( .a(n_335), .b(n_43704), .c(FE_OFN3_n_43918), .o(n_43746) );
na02f80 g768128 ( .a(n_12716), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_), .o(n_12809) );
no02f80 g755532 ( .a(n_24621), .b(n_24620), .o(n_24622) );
na02f80 g753130 ( .a(n_27296), .b(n_26398), .o(n_27347) );
no02f80 FE_RC_1113_0 ( .a(FE_RN_335_0), .b(n_6716), .o(n_6598) );
na02f80 g776093 ( .a(n_4717), .b(n_4716), .o(n_4789) );
in01f80 g763214 ( .a(n_17199), .o(n_17142) );
in01f80 newInst_1247 ( .a(newNet_1246), .o(newNet_1247) );
no02f80 g771139 ( .a(n_9623), .b(FE_OCPN3769_FE_OCP_RBN2375_n_8221), .o(n_9663) );
in01f80 g766004 ( .a(n_14763), .o(n_14783) );
no03m80 g756165 ( .a(n_24162), .b(n_24164), .c(n_23763), .o(n_24177) );
oa22f80 g781278 ( .a(n_46055), .b(beta_28), .c(n_7), .d(n_88), .o(n_278) );
oa12f80 g744581 ( .a(n_35180), .b(FE_OCP_RBN1374_n_35275), .c(n_35294), .o(n_35319) );
in01f80 newInst_791 ( .a(newNet_62), .o(newNet_791) );
in01f80 g737045 ( .a(n_43205), .o(n_43206) );
in01f80 g750476 ( .a(n_29587), .o(n_29588) );
in01f80 FE_OCP_RBC2174_n_37559 ( .a(n_37559), .o(FE_OCP_RBN2174_n_37559) );
no02f80 FE_RC_4208_0 ( .a(FE_RN_1841_0), .b(n_19806), .o(FE_RN_1842_0) );
in01f80 newInst_1501 ( .a(newNet_577), .o(newNet_1501) );
in01f80 g742052 ( .a(n_37975), .o(n_38332) );
in01f80 newInst_3747 ( .a(newNet_2459), .o(newNet_3747) );
in01f80 g752238 ( .a(n_28037), .o(n_28096) );
ao22s80 FE_RC_4115_0 ( .a(n_35135), .b(n_35289), .c(n_35137), .d(n_35288), .o(n_35383) );
in01f80 g779197 ( .a(n_1887), .o(n_1888) );
in01f80 newInst_1184 ( .a(newNet_1183), .o(newNet_1184) );
no02f80 g755635 ( .a(n_24435), .b(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24626) );
in01f80 g741303 ( .a(n_38959), .o(n_38905) );
in01f80 g743982 ( .a(n_35916), .o(n_35864) );
in01f80 newInst_2423 ( .a(newNet_2422), .o(newNet_2423) );
in01f80 g757458 ( .a(n_23011), .o(n_23012) );
oa22f80 g779856 ( .a(n_44659), .b(n_973), .c(n_44623), .d(n_899), .o(n_1288) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_5_ ( .ck(newNet_1471), .d(n_31691), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_) );
na02f80 g750342 ( .a(n_30662), .b(n_30158), .o(n_30719) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_31_ ( .ck(newNet_1188), .d(FE_OFN775_n_46137), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01f80 g759337 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .o(n_22608) );
na02f80 g781061 ( .a(sin_out_31), .b(FE_OFN5_n_43918), .o(n_295) );
na02f80 g763324 ( .a(n_17178), .b(n_17215), .o(n_17382) );
oa12f80 g741904 ( .a(n_38260), .b(n_38320), .c(n_38228), .o(n_38380) );
no02f80 g758038 ( .a(n_22844), .b(n_22843), .o(n_22923) );
no02f80 g764327 ( .a(n_16418), .b(n_16422), .o(n_16426) );
na02f80 g765268 ( .a(n_15573), .b(n_15572), .o(n_15574) );
na02f80 g750859 ( .a(n_29055), .b(FE_OCP_RBN1153_n_29053), .o(n_29139) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_7_ ( .ck(newNet_431), .d(n_27836), .o(delay_xor_ln22_unr18_stage7_stallmux_q_7_) );
oa12f80 g776742 ( .a(n_3917), .b(n_4028), .c(n_3862), .o(n_4029) );
oa22f80 FE_RC_418_0 ( .a(n_14824), .b(n_14465), .c(n_14464), .d(n_14891), .o(n_14962) );
no02f80 g750599 ( .a(n_45760), .b(FE_OFN788_n_25834), .o(n_29423) );
in01f80 g742625 ( .a(n_37488), .o(n_37489) );
na02f80 g743817 ( .a(n_36335), .b(n_36306), .o(n_36308) );
ao12f80 g757227 ( .a(n_22954), .b(n_23495), .c(n_22809), .o(n_23521) );
in01f80 g772238 ( .a(n_8799), .o(n_8833) );
na02f80 g769261 ( .a(n_11455), .b(n_11012), .o(n_11485) );
oa22f80 FE_RC_261_0 ( .a(n_20208), .b(n_20266), .c(n_20265), .d(n_20207), .o(n_20299) );
na03f80 g779329 ( .a(n_1715), .b(n_1648), .c(n_1714), .o(n_1742) );
na02f80 g772851 ( .a(n_8071), .b(n_7802), .o(n_8072) );
in01f80 newInst_1667 ( .a(newNet_1582), .o(newNet_1667) );
no02f80 g759470 ( .a(n_21029), .b(n_21028), .o(n_21144) );
na02f80 FE_RC_3027_0 ( .a(n_20997), .b(n_20628), .o(FE_RN_1326_0) );
na02f80 g756173 ( .a(n_24145), .b(n_23771), .o(n_24183) );
in01f80 g759888 ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_21852) );
in01f80 FE_RC_597_0 ( .a(n_25479), .o(FE_RN_186_0) );
oa22f80 g779883 ( .a(n_44659), .b(n_1066), .c(n_44623), .d(n_1028), .o(n_1346) );
no02f80 g737707 ( .a(n_42394), .b(n_42390), .o(n_42420) );
oa12f80 g742776 ( .a(n_37074), .b(n_37281), .c(n_36958), .o(n_37320) );
in01f80 g769446 ( .a(n_11527), .o(n_11655) );
na02f80 g754720 ( .a(n_26541), .b(n_26605), .o(n_26641) );
in01f80 fopt782874 ( .a(n_44311), .o(n_44309) );
in01f80 g756400 ( .a(n_23691), .o(n_23692) );
na02f80 g779610 ( .a(n_1794), .b(n_1584), .o(n_1802) );
no02f80 g748903 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .o(n_32499) );
ao12f80 g747950 ( .a(n_33123), .b(n_33122), .c(n_33121), .o(n_33720) );
in01f80 g763344 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_17_), .o(n_16921) );
in01f80 FE_OCP_RBC2265_n_29033 ( .a(FE_OCP_RBN2264_n_29033), .o(FE_OCP_RBN2265_n_29033) );
in01f80 g740985 ( .a(n_39137), .o(n_39138) );
in01f80 FE_OCP_RBC1220_n_27835 ( .a(n_27835), .o(FE_OCP_RBN1220_n_27835) );
in01f80 g780309 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n_1633) );
in01f80 newInst_181 ( .a(newNet_110), .o(newNet_181) );
in01f80 newInst_1231 ( .a(newNet_1011), .o(newNet_1231) );
in01f80 g772678 ( .a(n_8344), .o(n_8345) );
in01f80 g765542 ( .a(n_46419), .o(n_15219) );
in01f80 g759231 ( .a(n_21381), .o(n_21382) );
in01f80 newInst_300 ( .a(newNet_86), .o(newNet_300) );
na02f80 g740273 ( .a(n_40051), .b(n_40170), .o(n_40212) );
in01f80 g743240 ( .a(n_36802), .o(n_36803) );
in01f80 FE_RC_3193_0 ( .a(n_7245), .o(FE_RN_1418_0) );
in01f80 g761640 ( .a(n_18797), .o(n_18761) );
no02f80 g755934 ( .a(n_24290), .b(n_24309), .o(n_24429) );
oa22f80 g743690 ( .a(n_36248), .b(n_36240), .c(n_36279), .d(n_36241), .o(n_36377) );
no02f80 g763405 ( .a(FE_OCP_RBN3724_n_16975), .b(FE_OCP_RBN3689_n_16146), .o(n_17179) );
na02f80 g740217 ( .a(n_39890), .b(n_39942), .o(n_39941) );
in01f80 g740039 ( .a(n_40293), .o(n_40294) );
no02f80 g761502 ( .a(n_19573), .b(n_19572), .o(n_19574) );
oa22f80 g757787 ( .a(n_22358), .b(n_22108), .c(n_22391), .d(n_22109), .o(n_22540) );
in01f80 newInst_3734 ( .a(newNet_456), .o(newNet_3734) );
in01f80 g770975 ( .a(n_9762), .o(n_9856) );
na02f80 g784397 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .o(n_46209) );
in01f80 g744029 ( .a(n_35596), .o(n_35597) );
oa12f80 g768908 ( .a(n_11843), .b(n_11842), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_), .o(n_12747) );
in01f80 g756606 ( .a(n_23683), .o(n_23657) );
no02f80 g780716 ( .a(n_622), .b(n_621), .o(n_623) );
na02f80 g771765 ( .a(n_8990), .b(FE_OCP_RBN3571_n_44563), .o(n_9040) );
oa12f80 g778776 ( .a(n_1935), .b(n_2189), .c(n_1903), .o(n_2240) );
in01f80 g762413 ( .a(n_18522), .o(n_18523) );
na02f80 g747483 ( .a(FE_OCP_RBN3333_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .o(n_32592) );
in01f80 g755543 ( .a(n_24778), .o(n_24746) );
oa12f80 g751924 ( .a(n_28905), .b(n_28919), .c(n_28862), .o(n_29254) );
in01f80 g744683 ( .a(n_35237), .o(n_35238) );
na02f80 g775003 ( .a(n_6108), .b(FE_OCP_RBN2930_n_5221), .o(n_6234) );
na02f80 g754940 ( .a(n_25150), .b(n_24055), .o(n_25277) );
na02f80 g778918 ( .a(n_2243), .b(n_2265), .o(n_2286) );
no02f80 g743619 ( .a(n_36467), .b(n_36009), .o(n_36502) );
na02f80 g745011 ( .a(n_36315), .b(n_35808), .o(n_36385) );
na02f80 g775011 ( .a(n_6098), .b(n_5844), .o(n_6133) );
oa12f80 g754445 ( .a(n_25397), .b(n_25597), .c(n_25331), .o(n_25655) );
na02f80 g738137 ( .a(n_42021), .b(n_42020), .o(n_42022) );
in01f80 g740779 ( .a(n_39531), .o(n_39546) );
na02f80 g756910 ( .a(n_23648), .b(n_23647), .o(n_23649) );
na02f80 g745880 ( .a(n_33986), .b(n_34041), .o(n_34101) );
in01f80 newInst_1865 ( .a(newNet_1864), .o(newNet_1865) );
na02f80 g768088 ( .a(FE_OCPN860_n_12880), .b(n_13073), .o(n_13109) );
na02f80 g768253 ( .a(n_12571), .b(n_12371), .o(n_12589) );
oa12f80 g773959 ( .a(n_6901), .b(n_6900), .c(n_6899), .o(n_7690) );
oa22f80 g742169 ( .a(FE_OCP_RBN2240_n_44881), .b(n_37838), .c(FE_OCP_RBN3427_n_44881), .d(n_37823), .o(n_38211) );
no02f80 g769660 ( .a(n_11248), .b(n_46424), .o(n_11296) );
na02f80 g757989 ( .a(n_22305), .b(n_22220), .o(n_22306) );
oa12f80 g751918 ( .a(n_28160), .b(n_28186), .c(n_28112), .o(n_28255) );
in01f80 g772455 ( .a(n_8381), .o(n_8382) );
no02f80 g757246 ( .a(n_23132), .b(n_23226), .o(n_23210) );
in01f80 g741497 ( .a(n_38744), .o(n_38745) );
in01f80 g767874 ( .a(n_12823), .o(n_12929) );
no02f80 g749913 ( .a(n_29960), .b(n_30018), .o(n_30406) );
na02f80 g736965 ( .a(n_43120), .b(n_43250), .o(n_43350) );
in01f80 g738558 ( .a(n_41740), .o(n_41741) );
ao12f80 g776391 ( .a(n_4019), .b(n_4154), .c(n_4149), .o(n_4323) );
na02f80 g749453 ( .a(n_30500), .b(n_27014), .o(n_30537) );
no02f80 g756635 ( .a(n_24190), .b(n_24037), .o(n_24078) );
in01f80 g739723 ( .a(n_40503), .o(n_40504) );
in01f80 g765840 ( .a(n_14925), .o(n_14926) );
no02f80 g778048 ( .a(n_3042), .b(n_3028), .o(n_3128) );
no02f80 g767432 ( .a(n_13494), .b(n_13208), .o(n_13545) );
no02f80 g755878 ( .a(n_25055), .b(n_25033), .o(n_25471) );
in01f80 FE_OCP_RBC3385_n_33108 ( .a(n_33108), .o(FE_OCP_RBN3385_n_33108) );
no02f80 g753217 ( .a(n_27120), .b(n_26011), .o(n_27223) );
no02f80 g757976 ( .a(n_22481), .b(n_44287), .o(n_22347) );
in01f80 newInst_1125 ( .a(newNet_1124), .o(newNet_1125) );
in01f80 FE_OCP_RBC3028_n_39942 ( .a(FE_OCP_RBN3024_n_39942), .o(FE_OCP_RBN3028_n_39942) );
na02f80 g773415 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .o(n_7695) );
in01f80 newInst_1146 ( .a(newNet_1145), .o(newNet_1146) );
oa22f80 FE_RC_1090_0 ( .a(n_34394), .b(n_34880), .c(n_34395), .d(n_34881), .o(n_34982) );
in01f80 g744889 ( .a(n_35136), .o(n_35096) );
in01f80 g752132 ( .a(n_28093), .o(n_28094) );
ao12f80 g740202 ( .a(n_39772), .b(n_39753), .c(n_39750), .o(n_39824) );
in01f80 FE_OCP_RBC2902_n_44174 ( .a(FE_OCP_RBN2901_n_44174), .o(FE_OCP_RBN2902_n_44174) );
na02f80 g737867 ( .a(n_42406), .b(n_42383), .o(n_42480) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_6_ ( .ck(newNet_614), .d(n_46372), .o(delay_xor_ln21_unr9_stage4_stallmux_q_6_) );
oa22f80 FE_RC_1478_0 ( .a(n_28336), .b(n_32358), .c(n_32287), .d(n_32384), .o(n_32431) );
no02f80 g761826 ( .a(n_19125), .b(n_18730), .o(n_19191) );
in01f80 FE_OCPC1780_n_24097 ( .a(FE_OCPN1779_n_24097), .o(FE_OCPN1780_n_24097) );
in01f80 g738179 ( .a(n_42066), .o(n_42048) );
in01f80 g778694 ( .a(n_2571), .o(n_2635) );
in01f80 g751499 ( .a(n_28676), .o(n_28677) );
no02f80 g779317 ( .a(n_1691), .b(n_1690), .o(n_1692) );
in01f80 g737981 ( .a(n_42270), .o(n_42547) );
oa12f80 g747140 ( .a(n_33391), .b(n_33952), .c(n_33884), .o(n_34000) );
oa22f80 g775472 ( .a(n_45322), .b(n_5098), .c(n_45321), .d(n_5099), .o(n_5444) );
ao12f80 g742790 ( .a(n_37332), .b(n_37331), .c(n_37330), .o(n_37384) );
no02f80 g755814 ( .a(n_24426), .b(FE_OCP_DRV_N3154_n_24425), .o(n_24494) );
na02f80 g771790 ( .a(n_9955), .b(n_9877), .o(n_9956) );
ao12f80 g742650 ( .a(n_37199), .b(n_37380), .c(n_37375), .o(n_37429) );
na02f80 g736749 ( .a(n_43197), .b(n_43144), .o(n_43224) );
oa12f80 g738940 ( .a(n_41236), .b(n_41235), .c(n_41234), .o(n_41626) );
na02f80 g745302 ( .a(n_35932), .b(n_35931), .o(n_35933) );
ao12f80 g742661 ( .a(n_37484), .b(n_37483), .c(n_37482), .o(n_37618) );
no02f80 g742179 ( .a(n_44887), .b(n_38269), .o(n_38303) );
in01f80 newInst_1903 ( .a(newNet_1447), .o(newNet_1903) );
no02f80 g738579 ( .a(n_41560), .b(n_41481), .o(n_41612) );
no02f80 g742801 ( .a(n_37256), .b(n_37120), .o(n_37287) );
no02f80 g755826 ( .a(n_25034), .b(n_25090), .o(n_25091) );
in01f80 newInst_645 ( .a(newNet_644), .o(newNet_645) );
na02f80 FE_RC_15_0 ( .a(FE_RN_3_0), .b(FE_RN_4_0), .o(FE_RN_5_0) );
no02f80 g739239 ( .a(n_40738), .b(n_40674), .o(n_41086) );
oa22f80 FE_RC_1224_0 ( .a(n_6555), .b(n_6453), .c(n_6454), .d(n_6581), .o(n_6719) );
ao12f80 g780248 ( .a(n_684), .b(n_786), .c(n_698), .o(n_837) );
in01f80 newInst_63 ( .a(newNet_62), .o(newNet_63) );
in01f80 newInst_1882 ( .a(newNet_481), .o(newNet_1882) );
na02f80 g773402 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n_7621) );
ao12f80 g750290 ( .a(n_29641), .b(n_29720), .c(n_29602), .o(n_29790) );
in01f80 g780445 ( .a(n_784), .o(n_1061) );
na02f80 FE_RC_2903_0 ( .a(n_20024), .b(FE_RN_1259_0), .o(FE_RN_1260_0) );
in01f80 newInst_922 ( .a(newNet_921), .o(newNet_922) );
in01f80 g740874 ( .a(n_39264), .o(n_39239) );
na02f80 g742247 ( .a(n_37848), .b(n_37847), .o(n_37867) );
no02f80 g745247 ( .a(n_34465), .b(n_34438), .o(n_34439) );
na02f80 g778489 ( .a(n_2320), .b(n_2870), .o(n_2372) );
na02f80 g744573 ( .a(n_35290), .b(n_35211), .o(n_35333) );
in01f80 g768456 ( .a(n_12391), .o(n_12392) );
na02f80 g773949 ( .a(n_6990), .b(n_5268), .o(n_7063) );
no02f80 g774834 ( .a(n_6315), .b(n_5439), .o(n_6345) );
na02f80 g749775 ( .a(n_31340), .b(n_31339), .o(n_31341) );
in01f80 g742479 ( .a(n_37657), .o(n_37658) );
no02f80 FE_RC_1822_0 ( .a(n_35118), .b(n_35294), .o(FE_RN_544_0) );
no02f80 g778111 ( .a(n_2760), .b(n_2875), .o(n_2925) );
na02f80 g754067 ( .a(n_26032), .b(n_26064), .o(n_26188) );
na02f80 g737030 ( .a(n_43020), .b(FE_OCPN3777_n_43019), .o(n_43051) );
oa22f80 g758656 ( .a(n_21833), .b(n_21838), .c(n_21834), .d(n_21839), .o(n_21915) );
no02f80 g762597 ( .a(n_18069), .b(n_18086), .o(n_18160) );
no02f80 g740247 ( .a(n_40273), .b(n_40193), .o(n_40314) );
in01f80 newInst_846 ( .a(newNet_845), .o(newNet_846) );
in01f80 newInst_3065 ( .a(newNet_2475), .o(newNet_3065) );
in01f80 g756701 ( .a(n_23551), .o(n_23572) );
in01f80 FE_OCP_RBC2609_n_3807 ( .a(FE_OCP_RBN2608_n_3807), .o(FE_OCP_RBN2609_n_3807) );
in01f80 newInst_1415 ( .a(newNet_1414), .o(newNet_1415) );
oa12f80 g756369 ( .a(n_24302), .b(n_24301), .c(n_24300), .o(n_25085) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_11_ ( .ck(newNet_2495), .d(n_31955), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_) );
oa22f80 g758374 ( .a(n_21966), .b(n_21894), .c(n_21965), .d(n_21893), .o(n_22016) );
oa12f80 g739691 ( .a(n_40373), .b(n_40524), .c(n_40191), .o(n_40532) );
in01f80 g766400 ( .a(n_14533), .o(n_14496) );
na02f80 g739821 ( .a(n_40300), .b(n_39944), .o(n_40406) );
in01f80 g740822 ( .a(n_39538), .o(n_39488) );
na02f80 g755271 ( .a(n_25144), .b(n_25094), .o(n_25279) );
no02f80 g754692 ( .a(FE_OCPN928_n_26231), .b(n_26509), .o(n_26548) );
no02f80 FE_RC_2736_0 ( .a(FE_RN_1159_0), .b(n_44954), .o(n_39063) );
in01f80 g776404 ( .a(n_4809), .o(n_4810) );
ao12f80 g738271 ( .a(n_41673), .b(n_41844), .c(n_41577), .o(n_41928) );
ao12f80 g746187 ( .a(n_34615), .b(n_35087), .c(n_35041), .o(n_35111) );
in01f80 g753430 ( .a(n_27073), .o(n_27036) );
oa12f80 g751407 ( .a(n_28316), .b(n_28477), .c(n_28341), .o(n_28535) );
in01f80 g748665 ( .a(n_31488), .o(n_31484) );
in01f80 g742028 ( .a(n_38138), .o(n_38139) );
na02f80 g747094 ( .a(n_32928), .b(n_32682), .o(n_32929) );
in01f80 newInst_2725 ( .a(newNet_2724), .o(newNet_2725) );
no02f80 g779618 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .o(n_1945) );
ao12f80 g748060 ( .a(n_32883), .b(n_32882), .c(n_32881), .o(n_33512) );
no02f80 g738537 ( .a(n_41379), .b(n_41430), .o(n_41380) );
no02f80 g760001 ( .a(n_20667), .b(FE_OCP_RBN3662_n_20750), .o(n_20749) );
no02f80 g768355 ( .a(n_12459), .b(n_12053), .o(n_12514) );
no02f80 g738367 ( .a(n_41705), .b(n_41678), .o(n_41978) );
in01f80 g736537 ( .a(n_43665), .o(n_43670) );
ao12f80 g740844 ( .a(n_39244), .b(n_39310), .c(n_39304), .o(n_39349) );
in01f80 g752934 ( .a(n_27949), .o(n_28025) );
na02f80 g747225 ( .a(n_33798), .b(n_33797), .o(n_33799) );
na02f80 g773136 ( .a(n_7817), .b(n_7723), .o(n_7857) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_13_ ( .ck(newNet_462), .d(n_27838), .o(delay_xor_ln22_unr18_stage7_stallmux_q_13_) );
in01f80 FE_OCP_RBC2253_n_13017 ( .a(FE_OCP_RBN2251_n_13017), .o(FE_OCP_RBN2253_n_13017) );
no02f80 g765789 ( .a(FE_OCP_RBN3609_n_14905), .b(n_14215), .o(n_14957) );
in01f80 newInst_3216 ( .a(newNet_3215), .o(newNet_3216) );
no02f80 g754489 ( .a(n_25629), .b(n_25628), .o(n_25630) );
na02f80 g748595 ( .a(n_32723), .b(n_32491), .o(n_32724) );
in01f80 g747847 ( .a(n_32061), .o(n_32062) );
na02f80 g755891 ( .a(n_25254), .b(FE_RN_865_0), .o(n_25905) );
in01f80 FE_OCP_RBC2231_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2231_n_13141) );
no02f80 g770238 ( .a(n_10619), .b(n_10305), .o(n_10668) );
in01f80 g767466 ( .a(n_13501), .o(n_13502) );
no02f80 g739908 ( .a(n_40374), .b(n_40111), .o(n_40376) );
in01f80 FE_RC_2209_0 ( .a(n_20345), .o(FE_RN_795_0) );
in01f80 g776444 ( .a(n_4578), .o(n_4579) );
in01f80 fopt783577 ( .a(n_17689), .o(n_45205) );
in01f80 g766671 ( .a(n_13883), .o(n_13913) );
na02f80 g752917 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .o(n_27951) );
ao12f80 g750023 ( .a(n_29957), .b(FE_OCPN1786_n_30134), .c(FE_OCP_RBN1905_n_29080), .o(n_30493) );
in01f80 FE_RC_2447_0 ( .a(n_13109), .o(FE_RN_977_0) );
ao12f80 g777711 ( .a(n_3352), .b(n_3367), .c(n_3351), .o(n_4970) );
no02f80 g760707 ( .a(n_19666), .b(FE_OCP_DRV_N1564_n_19665), .o(n_19750) );
no02f80 g777288 ( .a(n_3788), .b(n_3771), .o(n_3815) );
na02f80 g764282 ( .a(n_16286), .b(n_16221), .o(n_16405) );
in01f80 g763373 ( .a(n_17081), .o(n_17082) );
in01f80 g757460 ( .a(n_22937), .o(n_22938) );
in01f80 g748552 ( .a(n_31449), .o(n_31466) );
na02f80 g766556 ( .a(FE_OCP_RBN2413_n_13960), .b(FE_OCP_RBN3507_n_13860), .o(n_14056) );
na02f80 g752024 ( .a(n_28072), .b(n_28101), .o(n_28188) );
in01f80 g771737 ( .a(n_8870), .o(n_8871) );
no02f80 g750108 ( .a(n_29857), .b(n_30136), .o(n_30470) );
in01f80 g740434 ( .a(n_39750), .o(n_39797) );
in01f80 g742490 ( .a(n_37646), .o(n_37626) );
na02f80 g769061 ( .a(n_11689), .b(FE_OCP_RBN3266_n_45224), .o(n_11993) );
ao12f80 g755668 ( .a(n_25439), .b(n_25438), .c(n_25437), .o(n_26419) );
in01f80 g767034 ( .a(n_13974), .o(n_14042) );
na02f80 g775248 ( .a(n_6011), .b(n_6002), .o(n_6116) );
ao22s80 FE_RC_621_0 ( .a(n_25395), .b(n_25634), .c(n_25394), .d(n_25655), .o(n_25763) );
in01f80 newInst_2430 ( .a(newNet_1576), .o(newNet_2430) );
ms00f80 cos_out_reg_18_ ( .ck(newNet_3733), .d(n_43851), .o(cos_out_18) );
na02f80 g743335 ( .a(n_36705), .b(n_36717), .o(n_36736) );
in01f80 g768271 ( .a(n_12585), .o(n_12586) );
in01f80 g750094 ( .a(n_29893), .o(n_29920) );
no02f80 g738113 ( .a(n_42105), .b(n_42083), .o(n_42084) );
in01f80 g764757 ( .a(FE_OCP_RBN2802_n_15706), .o(n_16940) );
no02f80 g753815 ( .a(n_26433), .b(n_23509), .o(n_26434) );
ao12f80 g737749 ( .a(n_42206), .b(n_42205), .c(n_42204), .o(n_43016) );
na02f80 g766681 ( .a(n_13774), .b(n_13279), .o(n_13857) );
no02f80 g771659 ( .a(n_8919), .b(n_8968), .o(n_8970) );
na02f80 g743049 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_36954) );
na02f80 g772904 ( .a(n_7791), .b(n_7804), .o(n_9003) );
no02f80 g760860 ( .a(n_19391), .b(n_19364), .o(n_19513) );
no02f80 g760658 ( .a(n_19702), .b(n_19750), .o(n_19810) );
in01f80 FE_OCP_RBC2607_n_3807 ( .a(n_3807), .o(FE_OCP_RBN2607_n_3807) );
na02f80 g775702 ( .a(n_5450), .b(n_5411), .o(n_5556) );
in01f80 FE_RC_3570_0 ( .a(n_24419), .o(FE_RN_1552_0) );
in01f80 g755371 ( .a(n_24896), .o(n_24915) );
no02f80 g761082 ( .a(n_19112), .b(n_19017), .o(n_19213) );
in01f80 FE_OCPUNCOC1807_n_31435 ( .a(n_31435), .o(FE_OCPUNCON1807_n_31435) );
na02f80 g746041 ( .a(n_33833), .b(n_33733), .o(n_33834) );
na02f80 g778286 ( .a(n_2529), .b(n_2085), .o(n_2638) );
na02f80 g761892 ( .a(n_18405), .b(n_18404), .o(n_18481) );
in01f80 fopt784007 ( .a(n_45739), .o(n_45738) );
na02f80 g771553 ( .a(n_9276), .b(n_9355), .o(n_9397) );
na02f80 g770951 ( .a(n_10043), .b(n_8427), .o(n_10165) );
no02f80 g777688 ( .a(n_3332), .b(n_2640), .o(n_3377) );
na02f80 g742031 ( .a(n_38001), .b(n_44875), .o(n_38118) );
in01f80 newInst_1566 ( .a(newNet_1302), .o(newNet_1566) );
na02f80 g770711 ( .a(n_10058), .b(n_9984), .o(n_10198) );
in01f80 newInst_249 ( .a(newNet_248), .o(newNet_249) );
no02f80 g780763 ( .a(n_523), .b(n_522), .o(n_524) );
no02f80 g754029 ( .a(n_26911), .b(n_26484), .o(n_26976) );
ao12f80 g737624 ( .a(n_42368), .b(n_42303), .c(n_42202), .o(n_42398) );
no03m80 g742476 ( .a(n_37605), .b(FE_OCP_RBN2184_FE_RN_464_0), .c(n_37659), .o(n_37717) );
in01f80 g756212 ( .a(n_24181), .o(n_24161) );
in01f80 g739769 ( .a(n_40462), .o(n_40463) );
no02f80 g741587 ( .a(n_38604), .b(n_38590), .o(n_38655) );
na02f80 g760400 ( .a(n_20167), .b(FE_OCPN1438_FE_OCP_RBN1330_n_18866), .o(n_20224) );
na02f80 FE_RC_3129_0 ( .a(n_30703), .b(n_30944), .o(FE_RN_1387_0) );
in01f80 FE_OCP_RBC2362_n_13785 ( .a(n_13785), .o(FE_OCP_RBN2362_n_13785) );
in01f80 g775031 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_24_), .o(n_6142) );
ao12f80 g762852 ( .a(n_17747), .b(n_17771), .c(n_17746), .o(n_19138) );
na02f80 FE_RC_1861_0 ( .a(n_14000), .b(FE_RN_570_0), .o(FE_RN_571_0) );
na02f80 g738402 ( .a(n_41830), .b(n_41808), .o(n_41856) );
na02f80 g749299 ( .a(n_30608), .b(n_27062), .o(n_30629) );
no02f80 FE_RC_2621_0 ( .a(n_44797), .b(FE_RN_1092_0), .o(n_40963) );
in01f80 g761612 ( .a(n_19647), .o(n_19787) );
no02f80 FE_RC_3591_0 ( .a(n_13514), .b(n_14321), .o(FE_RN_1567_0) );
na02f80 g738385 ( .a(n_41470), .b(n_41825), .o(n_41549) );
no02f80 g777744 ( .a(n_3350), .b(n_3325), .o(n_3403) );
na02f80 g776947 ( .a(n_3584), .b(n_3510), .o(n_3642) );
no02f80 g760608 ( .a(n_19783), .b(FE_OCPN1790_n_18119), .o(n_19816) );
oa12f80 g736272 ( .a(n_290), .b(n_43863), .c(FE_OFN3_n_43918), .o(n_43899) );
na02f80 g748070 ( .a(n_32844), .b(n_46107), .o(n_32880) );
na02f80 FE_RC_4060_0 ( .a(n_35640), .b(FE_RN_1766_0), .o(FE_RN_1767_0) );
in01f80 newInst_1065 ( .a(newNet_1064), .o(newNet_1065) );
na02f80 g750743 ( .a(n_29318), .b(n_29317), .o(n_29389) );
in01f80 newInst_2512 ( .a(newNet_818), .o(newNet_2512) );
na02f80 g742521 ( .a(n_37534), .b(n_37709), .o(n_37580) );
oa22f80 FE_RC_3424_0 ( .a(n_27366), .b(n_30888), .c(n_30708), .d(n_30943), .o(n_30965) );
no02f80 g767642 ( .a(n_13019), .b(n_13018), .o(n_13020) );
in01f80 g773000 ( .a(n_7999), .o(n_8000) );
na02f80 g742139 ( .a(n_38347), .b(n_38308), .o(n_38440) );
no02f80 g740122 ( .a(n_40217), .b(n_39872), .o(n_40320) );
oa22f80 g752206 ( .a(n_27871), .b(FE_OCP_RBN3308_n_44722), .c(n_44723), .d(delay_xor_ln22_unr18_stage7_stallmux_q_5_), .o(n_28011) );
in01f80 g779844 ( .a(n_1379), .o(n_1377) );
na02f80 g770036 ( .a(n_10806), .b(n_44511), .o(n_10886) );
na02f80 g750505 ( .a(n_29449), .b(n_29561), .o(n_29506) );
na02f80 FE_RC_3144_0 ( .a(n_31050), .b(FE_RN_1395_0), .o(n_31070) );
no02f80 g770969 ( .a(n_9848), .b(n_9803), .o(n_9992) );
in01f80 g758211 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n_22656) );
in01f80 g755519 ( .a(n_24874), .o(n_24797) );
in01f80 newInst_678 ( .a(newNet_677), .o(newNet_678) );
in01f80 g779512 ( .a(n_1453), .o(n_1454) );
in01f80 newInst_2748 ( .a(newNet_2747), .o(newNet_2748) );
na02f80 g749125 ( .a(n_30913), .b(n_30852), .o(n_30937) );
ao12f80 g773039 ( .a(n_7769), .b(n_7802), .c(n_7768), .o(n_7770) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_19_ ( .ck(newNet_241), .d(n_46183), .o(delay_xor_ln22_unr6_stage3_stallmux_q_19_) );
na02f80 FE_RC_3471_0 ( .a(n_39013), .b(n_39012), .o(FE_RN_1491_0) );
in01f80 g780909 ( .a(n_404), .o(n_405) );
in01f80 g746838 ( .a(n_33250), .o(n_33251) );
no02f80 g777356 ( .a(n_4556), .b(FE_OFN822_n_4597), .o(n_4622) );
in01f80 newInst_3700 ( .a(newNet_1625), .o(newNet_3700) );
in01f80 FE_RC_4093_0 ( .a(n_22187), .o(n_22249) );
in01f80 g745001 ( .a(n_34836), .o(n_34835) );
oa12f80 g781260 ( .a(n_107), .b(n_110), .c(n_46055), .o(n_144) );
na02f80 g775462 ( .a(n_5879), .b(n_5842), .o(n_5897) );
no02f80 g765017 ( .a(n_15789), .b(n_15721), .o(n_15933) );
in01f80 newInst_2622 ( .a(newNet_2621), .o(newNet_2622) );
in01f80 g768733 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n_12834) );
na02f80 g761312 ( .a(n_18918), .b(n_18945), .o(n_19030) );
ao12f80 g741774 ( .a(n_38401), .b(n_38400), .c(n_38399), .o(n_38471) );
in01f80 newInst_2843 ( .a(newNet_2552), .o(newNet_2843) );
na02f80 g738834 ( .a(n_44428), .b(n_41348), .o(n_41356) );
no02f80 g766545 ( .a(n_14018), .b(n_13437), .o(n_14057) );
in01f80 g754246 ( .a(n_25962), .o(n_25963) );
in01f80 g738764 ( .a(n_41374), .o(n_41375) );
in01f80 newInst_731 ( .a(newNet_20), .o(newNet_731) );
na02f80 g779251 ( .a(n_1795), .b(n_1768), .o(n_1769) );
no02f80 g767349 ( .a(n_13636), .b(n_13255), .o(n_13622) );
no02f80 g765154 ( .a(n_15455), .b(FE_OCPN3767_n_14439), .o(n_15456) );
no02f80 g771999 ( .a(FE_OCP_RBN3644_n_44490), .b(n_9598), .o(n_9772) );
in01f80 g749204 ( .a(n_30930), .o(n_30931) );
in01f80 newInst_579 ( .a(newNet_100), .o(newNet_579) );
no02f80 g742202 ( .a(n_44869), .b(n_37869), .o(n_37887) );
in01f80 newInst_2088 ( .a(newNet_2087), .o(newNet_2088) );
oa12f80 g764627 ( .a(n_15639), .b(n_15661), .c(n_15810), .o(n_15818) );
oa12f80 g760854 ( .a(n_19507), .b(n_19506), .c(n_19514), .o(n_21343) );
no02f80 g756556 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .o(n_23736) );
in01f80 newInst_854 ( .a(newNet_853), .o(newNet_854) );
na02f80 g740099 ( .a(n_40186), .b(n_39953), .o(n_40287) );
in01f80 fopt783780 ( .a(FE_OCP_RBN3212_n_44365), .o(n_45450) );
no02f80 g766876 ( .a(n_14304), .b(n_14210), .o(n_14343) );
oa12f80 g751267 ( .a(n_29748), .b(n_29747), .c(n_29746), .o(n_30063) );
in01f80 fopt783159 ( .a(n_40532), .o(n_44692) );
no02f80 g743968 ( .a(n_35827), .b(n_35785), .o(n_35786) );
no02f80 g736854 ( .a(n_43280), .b(n_43511), .o(n_43619) );
no02f80 g763695 ( .a(n_16719), .b(FE_OCP_RBN2741_n_15206), .o(n_16759) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_3_ ( .ck(newNet_1692), .d(n_21930), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_) );
in01f80 g780515 ( .a(n_1054), .o(n_1055) );
in01f80 g761054 ( .a(n_19372), .o(n_20523) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_12_ ( .ck(newNet_1427), .d(n_36496), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_) );
in01f80 FE_OCP_RBC1723_n_21004 ( .a(FE_OCP_RBN1722_n_21004), .o(FE_OCP_RBN1723_n_21004) );
in01f80 FE_OCP_RBC2700_n_4238 ( .a(FE_OCP_RBN2699_n_4238), .o(FE_OCP_RBN2700_n_4238) );
no02f80 g771211 ( .a(n_9092), .b(n_8309), .o(n_9195) );
no02f80 FE_RC_3081_0 ( .a(FE_RN_1358_0), .b(n_16518), .o(n_16570) );
na02f80 g770558 ( .a(n_10193), .b(FE_OFN756_n_44461), .o(n_10332) );
na02f80 g742643 ( .a(n_37420), .b(n_37419), .o(n_37421) );
in01f80 newInst_283 ( .a(newNet_282), .o(newNet_283) );
in01f80 FE_OCP_RBC2190_n_7346 ( .a(n_7346), .o(FE_OCP_RBN2190_n_7346) );
in01f80 newInst_1395 ( .a(newNet_1190), .o(newNet_1395) );
in01f80 g743693 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_13_), .o(n_36466) );
in01f80 newInst_1437 ( .a(newNet_1436), .o(newNet_1437) );
in01f80 g772617 ( .a(n_8396), .o(n_8419) );
in01f80 FE_RC_3967_0 ( .a(n_18548), .o(FE_RN_1719_0) );
no04s80 FE_RC_2334_0 ( .a(n_11844), .b(n_11737), .c(n_11881), .d(n_11882), .o(n_11956) );
in01f80 newInst_3021 ( .a(newNet_3020), .o(newNet_3021) );
no02f80 g743368 ( .a(n_37813), .b(n_37814), .o(n_37840) );
in01f80 g739468 ( .a(n_40802), .o(n_40803) );
no02f80 g760837 ( .a(n_19466), .b(n_19532), .o(n_19592) );
in01f80 g771468 ( .a(n_9166), .o(n_9167) );
ao12f80 g759801 ( .a(n_20244), .b(n_20379), .c(n_20285), .o(n_20476) );
no02f80 FE_RC_174_0 ( .a(FE_RN_54_0), .b(n_355), .o(n_379) );
no02f80 g759578 ( .a(n_20511), .b(n_20481), .o(n_20621) );
in01f80 g765659 ( .a(n_14987), .o(n_15014) );
na02f80 g751700 ( .a(n_28368), .b(n_28367), .o(n_28420) );
oa12f80 g744943 ( .a(n_36117), .b(n_36386), .c(n_35630), .o(n_36405) );
in01f80 g772641 ( .a(n_8321), .o(n_8322) );
no02f80 g748445 ( .a(n_31720), .b(n_31719), .o(n_31754) );
na02f80 g738330 ( .a(n_41862), .b(n_41699), .o(n_41863) );
in01f80 FE_OCP_RBC3508_n_13860 ( .a(FE_OCP_RBN3506_n_13860), .o(FE_OCP_RBN3508_n_13860) );
in01f80 g755775 ( .a(FE_OCP_RBN2366_n_24372), .o(n_24529) );
oa22f80 FE_RC_1703_0 ( .a(n_14618), .b(n_46982), .c(FE_OCP_RBN3669_n_46982), .d(n_14452), .o(n_15761) );
na02f80 g756482 ( .a(n_23684), .b(n_23656), .o(n_23685) );
in01f80 g760909 ( .a(n_20057), .o(n_20017) );
in01f80 g736558 ( .a(n_43573), .o(n_43574) );
no02f80 g745463 ( .a(n_34315), .b(n_34325), .o(n_34384) );
no02f80 g757090 ( .a(n_23263), .b(n_23322), .o(n_23324) );
no02f80 g755741 ( .a(n_24494), .b(n_24444), .o(n_24550) );
oa22f80 g758196 ( .a(n_22585), .b(n_21866), .c(n_22586), .d(n_21865), .o(n_22659) );
in01f80 g774403 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .o(n_6518) );
in01f80 g781397 ( .a(beta_20), .o(n_18) );
no02f80 g777401 ( .a(n_3627), .b(n_3626), .o(n_3749) );
in01f80 g764257 ( .a(n_16824), .o(n_16848) );
na02f80 FE_RC_2796_0 ( .a(n_33708), .b(n_34200), .o(FE_RN_1195_0) );
ao12f80 g738614 ( .a(n_41912), .b(n_41716), .c(n_41613), .o(n_42078) );
in01f80 FE_OCPC1396_n_7881 ( .a(FE_OCPN1395_n_7881), .o(FE_OCPN1396_n_7881) );
oa12f80 g739878 ( .a(n_40080), .b(n_40260), .c(n_39997), .o(n_40380) );
na02f80 g746214 ( .a(n_33820), .b(n_33917), .o(n_33822) );
in01f80 g744644 ( .a(n_35358), .o(n_35359) );
in01f80 g771248 ( .a(n_9788), .o(n_9789) );
na02f80 g738482 ( .a(n_41381), .b(n_41407), .o(n_41416) );
na02f80 g770331 ( .a(n_10541), .b(n_10241), .o(n_10573) );
in01f80 newInst_2134 ( .a(newNet_2133), .o(newNet_2134) );
in01f80 FE_RC_3143_0 ( .a(n_31025), .o(FE_RN_1395_0) );
na02f80 g745742 ( .a(n_34119), .b(n_34118), .o(n_34120) );
in01f80 g766511 ( .a(n_14032), .o(n_14002) );
no02f80 g767985 ( .a(n_12958), .b(n_12855), .o(n_13305) );
in01f80 g755981 ( .a(n_24251), .o(n_24252) );
in01f80 g742850 ( .a(n_37286), .o(n_37266) );
oa12f80 g751317 ( .a(n_28421), .b(n_28684), .c(n_28387), .o(n_28747) );
no02f80 g755893 ( .a(n_24362), .b(n_24361), .o(n_24442) );
in01f80 g754568 ( .a(n_26928), .o(n_26929) );
no02f80 g760725 ( .a(n_19637), .b(n_19463), .o(n_19640) );
na02f80 g759911 ( .a(n_21053), .b(n_21052), .o(n_21107) );
oa12f80 g739018 ( .a(n_41104), .b(n_41103), .c(n_41102), .o(n_41141) );
in01f80 g776029 ( .a(n_4800), .o(n_4801) );
na02f80 g740269 ( .a(n_40030), .b(n_40028), .o(n_40056) );
in01f80 newInst_2707 ( .a(newNet_2706), .o(newNet_2707) );
in01f80 g738096 ( .a(n_42085), .o(n_42086) );
na02f80 g736753 ( .a(n_43184), .b(n_43217), .o(n_43185) );
in01f80 g746428 ( .a(n_33426), .o(n_34343) );
na02f80 g762833 ( .a(n_17906), .b(n_17867), .o(n_17940) );
no02f80 g745264 ( .a(n_35806), .b(FE_OCP_RBN2988_n_35539), .o(n_35968) );
in01f80 g762702 ( .a(n_17918), .o(n_17919) );
na02f80 FE_RC_2494_0 ( .a(FE_RN_1010_0), .b(n_1387), .o(n_1433) );
ao22s80 g771903 ( .a(FE_OCP_RBN2520_n_8762), .b(n_8671), .c(n_8762), .d(FE_OCPN1400_n_8670), .o(n_8904) );
in01f80 newInst_132 ( .a(newNet_131), .o(newNet_132) );
in01f80 g778611 ( .a(n_2817), .o(n_2762) );
in01f80 newInst_2855 ( .a(newNet_2854), .o(newNet_2855) );
ms00f80 sin_out_reg_2_ ( .ck(newNet_33), .d(n_43337), .o(sin_out_2) );
no02f80 g743899 ( .a(n_36270), .b(n_36200), .o(n_36271) );
no02f80 g773063 ( .a(n_7696), .b(n_7227), .o(n_7742) );
ao12f80 g757527 ( .a(n_23297), .b(n_23298), .c(n_23296), .o(n_23978) );
no02f80 g761474 ( .a(n_19845), .b(n_19844), .o(n_19953) );
oa12f80 g751504 ( .a(n_28718), .b(FE_OCP_RBN2192_n_28597), .c(n_28646), .o(n_28732) );
na02f80 g767755 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_), .o(n_13203) );
no02f80 g770435 ( .a(n_10452), .b(n_10449), .o(n_10582) );
no02f80 g781290 ( .a(n_46055), .b(beta_7), .o(n_63) );
in01f80 newInst_1828 ( .a(newNet_1827), .o(newNet_1828) );
no02f80 g767947 ( .a(n_12782), .b(n_12781), .o(n_12783) );
in01f80 newInst_2256 ( .a(newNet_2255), .o(newNet_2256) );
in01f80 g749839 ( .a(n_31185), .o(n_31186) );
oa12f80 g740212 ( .a(n_39774), .b(n_39792), .c(n_39758), .o(n_39861) );
na02f80 g763755 ( .a(n_16727), .b(n_16726), .o(n_16825) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_8_ ( .ck(newNet_1275), .d(n_1112), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_) );
in01f80 g767380 ( .a(n_13298), .o(n_13299) );
in01f80 g780159 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .o(n_1174) );
ao22s80 g774193 ( .a(n_6542), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN1986_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(delay_xor_ln21_unr6_stage3_stallmux_q_2_), .o(n_6616) );
no02f80 FE_RC_2748_0 ( .a(FE_RN_1167_0), .b(n_39106), .o(n_39165) );
no02f80 g773206 ( .a(n_7721), .b(n_7723), .o(n_7913) );
no02f80 g754051 ( .a(n_26070), .b(n_26105), .o(n_26173) );
oa22f80 FE_RC_1089_0 ( .a(n_36797), .b(n_36842), .c(n_36796), .d(n_36831), .o(n_36885) );
no02f80 g744215 ( .a(n_35900), .b(n_36001), .o(n_36093) );
in01f80 g750848 ( .a(n_29141), .o(n_29142) );
ao22s80 FE_RC_3864_0 ( .a(FE_RN_1687_0), .b(n_21847), .c(FE_RN_1688_0), .d(n_21736), .o(n_21953) );
na02f80 g740154 ( .a(n_39781), .b(n_39562), .o(n_39953) );
na02f80 g769128 ( .a(n_11579), .b(n_11619), .o(n_11743) );
in01f80 g765033 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_4_), .o(n_17478) );
no02f80 g756235 ( .a(n_24740), .b(n_24739), .o(n_24741) );
ao22s80 g784423 ( .a(n_36497), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_), .o(n_46235) );
no02f80 g779028 ( .a(n_2054), .b(n_2053), .o(n_2055) );
in01f80 FE_OCP_RBC2479_n_8530 ( .a(n_8530), .o(FE_OCP_RBN2479_n_8530) );
ao12f80 g770438 ( .a(n_10561), .b(n_10572), .c(n_10560), .o(n_10631) );
ao12f80 g756356 ( .a(n_24384), .b(n_24417), .c(n_24383), .o(n_25109) );
oa22f80 FE_RC_3359_0 ( .a(n_34745), .b(n_35050), .c(n_34746), .d(n_35049), .o(n_35130) );
no02f80 g766869 ( .a(n_13557), .b(FE_OCPN860_n_12880), .o(n_13574) );
in01f80 g740260 ( .a(n_40102), .o(n_40103) );
in01f80 g764956 ( .a(n_15545), .o(n_15546) );
no02f80 g753197 ( .a(n_27087), .b(n_25963), .o(n_27188) );
na02f80 g750546 ( .a(n_29378), .b(n_29379), .o(n_29406) );
oa12f80 g767828 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .c(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_12967) );
na02f80 g765007 ( .a(n_15321), .b(FE_OCP_RBN2356_n_13858), .o(n_15320) );
in01f80 g774937 ( .a(n_6176), .o(n_6177) );
ao12f80 g751023 ( .a(n_29837), .b(n_29884), .c(n_29935), .o(n_30001) );
no02f80 g744826 ( .a(n_35015), .b(n_35039), .o(n_35102) );
in01f80 g757830 ( .a(n_22569), .o(n_22590) );
oa12f80 g757416 ( .a(n_22867), .b(n_22940), .c(n_22994), .o(n_23071) );
na02f80 g747108 ( .a(n_34000), .b(n_33999), .o(n_34001) );
oa12f80 g749734 ( .a(n_29874), .b(n_29875), .c(n_29873), .o(n_31583) );
in01f80 g737784 ( .a(n_42641), .o(n_42642) );
no02f80 g743127 ( .a(n_36540), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_36949) );
in01f80 g746400 ( .a(n_33518), .o(n_33559) );
oa12f80 g776202 ( .a(n_4535), .b(n_4630), .c(n_4568), .o(n_4855) );
no02f80 g744277 ( .a(n_44174), .b(n_35659), .o(n_35740) );
in01f80 g774981 ( .a(n_6138), .o(n_6139) );
in01f80 g770597 ( .a(n_10274), .o(n_10292) );
na02f80 g755058 ( .a(n_25613), .b(n_25645), .o(n_25661) );
in01f80 newInst_2028 ( .a(newNet_2027), .o(newNet_2028) );
no02f80 g736644 ( .a(n_43374), .b(n_43271), .o(n_43375) );
in01f80 fopt783277 ( .a(n_14508), .o(n_44849) );
in01f80 FE_OCP_RBC3699_n_43015 ( .a(n_43015), .o(FE_OCP_RBN3699_n_43015) );
na02f80 g770551 ( .a(n_10527), .b(n_10491), .o(n_10492) );
oa12f80 g769301 ( .a(n_11425), .b(n_11405), .c(n_11476), .o(n_11477) );
no02f80 FE_RC_2713_0 ( .a(FE_RN_1141_0), .b(FE_RN_1143_0), .o(n_13098) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_2_ ( .ck(newNet_1968), .d(n_9916), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_2_) );
no02f80 g752988 ( .a(n_27086), .b(n_27154), .o(n_27234) );
in01f80 newInst_330 ( .a(newNet_291), .o(newNet_330) );
oa12f80 g773908 ( .a(n_7014), .b(n_7013), .c(n_7012), .o(n_7714) );
in01f80 g754549 ( .a(n_26903), .o(n_26904) );
oa12f80 g745112 ( .a(n_34176), .b(n_34683), .c(n_34618), .o(n_34717) );
no02f80 g779096 ( .a(n_2051), .b(n_1797), .o(n_2067) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_7_ ( .ck(newNet_1066), .d(n_10044), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_) );
in01f80 FE_OCP_RBC3848_FE_RN_1548_0 ( .a(FE_RN_1548_0), .o(FE_OCP_RBN3848_FE_RN_1548_0) );
in01f80 g753233 ( .a(n_27296), .o(n_27336) );
no02f80 g741842 ( .a(n_38386), .b(n_38385), .o(n_38387) );
no02f80 g742370 ( .a(n_37801), .b(n_37800), .o(n_37832) );
oa12f80 g757704 ( .a(n_22311), .b(n_22543), .c(n_22344), .o(n_22544) );
ao12f80 g757099 ( .a(n_23079), .b(n_44068), .c(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .o(n_23144) );
in01f80 g777194 ( .a(n_5415), .o(n_5416) );
no02f80 g770695 ( .a(n_10375), .b(n_10374), .o(n_10417) );
na02f80 g774987 ( .a(n_6083), .b(n_5983), .o(n_6144) );
oa22f80 g757677 ( .a(n_22625), .b(n_22419), .c(n_44322), .d(n_22416), .o(n_22819) );
na02f80 g769284 ( .a(n_11585), .b(n_11039), .o(n_11557) );
no02f80 g762918 ( .a(n_17994), .b(n_17464), .o(n_18013) );
na02f80 g752181 ( .a(n_27942), .b(n_27895), .o(n_28008) );
in01f80 g752015 ( .a(n_29187), .o(n_29267) );
ao12f80 FE_RC_3651_0 ( .a(FE_RN_1602_0), .b(n_21956), .c(n_21923), .o(n_22005) );
in01f80 newInst_1638 ( .a(newNet_1637), .o(newNet_1638) );
in01f80 g748278 ( .a(n_47271), .o(n_32068) );
in01f80 newInst_1725 ( .a(newNet_1724), .o(newNet_1725) );
in01f80 g768999 ( .a(n_11765), .o(n_11766) );
na02f80 g748308 ( .a(n_31475), .b(n_31502), .o(n_31503) );
in01f80 g766886 ( .a(n_14339), .o(n_14456) );
in01f80 FE_OCP_RBC2661_n_9292 ( .a(n_9292), .o(FE_OCP_RBN2661_n_9292) );
na02f80 g773398 ( .a(n_7562), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_), .o(n_7594) );
in01f80 g762067 ( .a(n_18224), .o(n_18225) );
na02f80 g780095 ( .a(n_1153), .b(n_1145), .o(n_1146) );
na02f80 g777595 ( .a(n_3415), .b(n_3452), .o(n_3817) );
oa22f80 g736904 ( .a(n_43242), .b(n_42967), .c(FE_OCPN1247_n_43120), .d(FE_OCP_RBN3000_n_42959), .o(n_43533) );
in01f80 g748881 ( .a(n_32454), .o(n_32417) );
in01f80 g745378 ( .a(n_35929), .o(n_35883) );
no02f80 g748387 ( .a(n_31518), .b(n_31448), .o(n_31605) );
in01f80 FE_OFC822_n_4597 ( .a(FE_OFN839_n_4597), .o(FE_OFN822_n_4597) );
no02f80 g755788 ( .a(n_24314), .b(n_24040), .o(n_24346) );
in01f80 g749162 ( .a(n_30933), .o(n_30954) );
na02f80 g764495 ( .a(n_16003), .b(FE_OCPN3775_n_14730), .o(n_16056) );
na02f80 g772801 ( .a(n_8141), .b(n_8140), .o(n_8142) );
in01f80 newInst_943 ( .a(newNet_488), .o(newNet_943) );
na02f80 g757607 ( .a(n_22583), .b(n_22276), .o(n_22720) );
na02f80 g739194 ( .a(n_40703), .b(n_45149), .o(n_40795) );
in01f80 fopt783282 ( .a(n_11853), .o(n_44859) );
na02f80 g776482 ( .a(n_4314), .b(n_3029), .o(n_4547) );
no02f80 g745732 ( .a(n_34365), .b(n_34364), .o(n_34396) );
in01f80 newInst_713 ( .a(newNet_429), .o(newNet_713) );
in01f80 FE_OCP_RBC2580_n_3734 ( .a(n_3734), .o(FE_OCP_RBN2580_n_3734) );
ao12f80 g773867 ( .a(n_7043), .b(n_7052), .c(n_7042), .o(n_7103) );
no02f80 g774789 ( .a(n_6240), .b(n_6230), .o(n_6231) );
in01f80 g772948 ( .a(n_7887), .o(n_7929) );
na02f80 g749892 ( .a(FE_OCP_RBN3013_n_31117), .b(n_30432), .o(n_31169) );
na02f80 g738241 ( .a(n_41931), .b(n_41930), .o(n_41932) );
in01f80 g755477 ( .a(n_24803), .o(n_24802) );
no02f80 g751190 ( .a(n_29800), .b(n_29799), .o(n_29819) );
in01f80 g770840 ( .a(n_9970), .o(n_9971) );
in01f80 newInst_2688 ( .a(newNet_2687), .o(newNet_2688) );
ao12f80 g764638 ( .a(n_15944), .b(n_46980), .c(n_16111), .o(n_16109) );
in01f80 g752981 ( .a(n_27075), .o(n_27088) );
in01f80 g775149 ( .a(n_6051), .o(n_6052) );
oa12f80 g753741 ( .a(n_26414), .b(n_26413), .c(n_26412), .o(n_26477) );
no02f80 g746898 ( .a(FE_OCP_RBN3384_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_26_), .o(n_33259) );
na02f80 g773035 ( .a(n_7951), .b(n_7998), .o(n_8061) );
in01f80 g736601 ( .a(n_43378), .o(n_43379) );
ao12f80 g745550 ( .a(n_34354), .b(FE_OCPN1732_n_34369), .c(n_34323), .o(n_34762) );
na02f80 g768653 ( .a(n_12187), .b(n_12251), .o(n_12287) );
no02f80 g763241 ( .a(n_17126), .b(n_17189), .o(n_17277) );
na02f80 g753455 ( .a(n_26914), .b(n_26982), .o(n_27004) );
na02f80 g751967 ( .a(n_28793), .b(n_28664), .o(n_28940) );
ao12f80 g767743 ( .a(n_12932), .b(n_12929), .c(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_13045) );
no02f80 g751411 ( .a(n_28531), .b(n_28571), .o(n_28581) );
ao12f80 g742628 ( .a(n_37153), .b(n_37373), .c(n_37296), .o(n_37427) );
in01f80 FE_OCP_RBC3504_n_38592 ( .a(FE_OCP_RBN3503_n_38592), .o(FE_OCP_RBN3504_n_38592) );
in01f80 g776459 ( .a(n_4346), .o(n_4347) );
na02f80 g780112 ( .a(n_1029), .b(n_1012), .o(n_1013) );
in01f80 g772480 ( .a(n_8537), .o(n_8538) );
in01f80 FE_OCP_RBC3265_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3265_n_45224) );
na02f80 g767412 ( .a(n_13359), .b(n_13403), .o(n_13449) );
no02f80 g743206 ( .a(n_38129), .b(n_38094), .o(n_38173) );
na02f80 g761188 ( .a(FE_OCP_RBN1685_n_18986), .b(n_17732), .o(n_19045) );
na02f80 g740542 ( .a(n_39644), .b(n_39647), .o(n_39667) );
no02f80 g760310 ( .a(FE_OCP_RBN3847_FE_RN_1548_0), .b(n_20223), .o(n_20279) );
ao12f80 g779447 ( .a(n_1599), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_10_), .o(n_1649) );
na03f80 FE_RC_3390_0 ( .a(n_16170), .b(n_16205), .c(n_16172), .o(n_16290) );
no02f80 g739910 ( .a(n_40374), .b(n_40227), .o(n_40373) );
in01f80 newInst_3149 ( .a(newNet_3148), .o(newNet_3149) );
na02f80 g773579 ( .a(n_7420), .b(n_7419), .o(n_7421) );
in01f80 g772752 ( .a(n_8138), .o(n_8139) );
oa22f80 g741097 ( .a(FE_OCP_RBN3629_n_38870), .b(n_38526), .c(FE_OCPN957_n_39096), .d(n_38510), .o(n_39362) );
oa12f80 g784072 ( .a(n_1002), .b(n_1194), .c(n_45812), .o(n_45818) );
in01f80 FE_OCP_RBC3503_n_38592 ( .a(FE_OCP_RBN3502_n_38592), .o(FE_OCP_RBN3503_n_38592) );
no02f80 g766830 ( .a(n_14426), .b(n_14425), .o(n_15442) );
ao22s80 FE_RC_3910_0 ( .a(n_47187), .b(n_21578), .c(n_21543), .d(n_47186), .o(n_21791) );
no02f80 FE_RC_3932_0 ( .a(FE_OCP_RBN3268_n_45224), .b(FE_RN_1700_0), .o(FE_RN_1701_0) );
na02f80 g780829 ( .a(n_582), .b(n_581), .o(n_627) );
oa12f80 g749226 ( .a(n_31283), .b(n_32156), .c(n_31368), .o(n_32201) );
in01f80 FE_RC_4203_0 ( .a(n_19561), .o(FE_RN_1840_0) );
no02f80 g760535 ( .a(n_19915), .b(FE_OFN814_n_18287), .o(n_19969) );
no02f80 g756802 ( .a(n_23370), .b(n_23407), .o(n_23519) );
in01f80 FE_OCP_RBC3402_n_28597 ( .a(FE_OCP_RBN2192_n_28597), .o(FE_OCP_RBN3402_n_28597) );
in01f80 newInst_572 ( .a(newNet_354), .o(newNet_572) );
na02f80 g748922 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .o(n_32491) );
na02f80 g767296 ( .a(n_13696), .b(n_13036), .o(n_13734) );
in01f80 newInst_3200 ( .a(newNet_44), .o(newNet_3200) );
oa12f80 g773514 ( .a(n_7478), .b(n_7477), .c(n_7476), .o(n_7522) );
no02f80 g779634 ( .a(n_1471), .b(n_1470), .o(n_1504) );
ao12f80 g756788 ( .a(n_23911), .b(n_23723), .c(n_23743), .o(n_23938) );
oa12f80 g756625 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_20_), .c(delay_add_ln22_unr14_stage6_stallmux_q_21_), .o(n_23734) );
in01f80 g774800 ( .a(n_6299), .o(n_6322) );
in01f80 newInst_973 ( .a(newNet_875), .o(newNet_973) );
in01f80 FE_RC_89_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .o(FE_RN_27_0) );
oa12f80 g747590 ( .a(n_31727), .b(n_45517), .c(FE_OCPN977_n_31594), .o(n_32226) );
na02f80 g751158 ( .a(n_30156), .b(n_29993), .o(n_30431) );
no02f80 g772888 ( .a(n_7987), .b(n_7932), .o(n_8064) );
ms00f80 mux_while_ln12_psv_q_reg_4_ ( .ck(newNet_112), .d(n_204), .o(mux_while_ln12_psv_q_4_) );
na02f80 g750737 ( .a(n_29215), .b(n_29111), .o(n_29235) );
in01f80 newInst_391 ( .a(newNet_390), .o(newNet_391) );
na02f80 g751616 ( .a(n_28467), .b(n_27711), .o(n_28509) );
na02f80 g766353 ( .a(n_14158), .b(n_14189), .o(n_14326) );
in01f80 g745964 ( .a(n_34076), .o(n_34077) );
in01f80 g754202 ( .a(n_26118), .o(n_26079) );
in01f80 newInst_3430 ( .a(newNet_3429), .o(newNet_3430) );
no02f80 g757019 ( .a(n_24059), .b(n_23061), .o(n_24149) );
na02f80 g777628 ( .a(n_3393), .b(n_3210), .o(n_3395) );
no02f80 g737913 ( .a(FE_OCPN1231_n_42201), .b(n_42478), .o(n_42545) );
in01f80 newInst_3709 ( .a(newNet_216), .o(newNet_3709) );
in01f80 FE_OCP_RBC1702_n_19560 ( .a(n_19560), .o(FE_OCP_RBN1702_n_19560) );
no02f80 g774791 ( .a(n_6324), .b(n_6219), .o(n_6354) );
no02f80 g764677 ( .a(n_15765), .b(n_14650), .o(n_15856) );
in01f80 FE_OCPC1853_n_13366 ( .a(n_13366), .o(FE_OCPN1853_n_13366) );
in01f80 FE_OCP_RBC3439_n_33803 ( .a(n_33803), .o(FE_OCP_RBN3439_n_33803) );
in01f80 g759741 ( .a(n_21863), .o(n_21864) );
na02f80 g749406 ( .a(n_31981), .b(n_31276), .o(n_31979) );
no02f80 g755116 ( .a(n_25315), .b(n_25318), .o(n_25415) );
na02f80 g775260 ( .a(n_5799), .b(n_5583), .o(n_5895) );
na03f80 FE_RC_615_0 ( .a(FE_OCP_RBN2139_n_17547), .b(n_17642), .c(n_17579), .o(n_17797) );
in01f80 g739002 ( .a(n_41185), .o(n_41205) );
na02f80 g766952 ( .a(n_14758), .b(n_14253), .o(n_14390) );
na02f80 g769227 ( .a(n_11556), .b(FE_OCP_RBN2870_n_10480), .o(n_11678) );
in01f80 g760279 ( .a(n_20372), .o(n_20404) );
na02f80 g780820 ( .a(n_361), .b(n_367), .o(n_382) );
no02f80 g754541 ( .a(n_26609), .b(n_26608), .o(n_26610) );
oa12f80 g771642 ( .a(n_8855), .b(n_8872), .c(n_8856), .o(n_8922) );
na02f80 g769708 ( .a(n_11270), .b(n_11291), .o(n_11369) );
oa12f80 g748698 ( .a(n_32495), .b(n_32532), .c(n_32499), .o(n_32606) );
na02f80 g775918 ( .a(n_4936), .b(FE_OCP_RBN2722_n_4219), .o(n_5013) );
oa22f80 g763041 ( .a(n_17294), .b(n_17584), .c(n_17290), .d(n_17753), .o(n_17418) );
oa22f80 FE_RC_1222_0 ( .a(FE_OFN84_n_46137), .b(n_6646), .c(FE_OFN806_n_46196), .d(n_6670), .o(n_46190) );
no02f80 g768072 ( .a(n_12709), .b(n_12699), .o(n_12749) );
na02f80 g750461 ( .a(n_29585), .b(n_29603), .o(n_29620) );
oa22f80 FE_RC_3737_0 ( .a(n_16396), .b(n_16609), .c(n_16397), .d(n_16626), .o(n_16719) );
na02f80 FE_RC_3504_0 ( .a(FE_OCP_RBN3309_n_44722), .b(FE_RN_1512_0), .o(n_27802) );
in01f80 newInst_1859 ( .a(newNet_566), .o(newNet_1859) );
na02f80 g768555 ( .a(n_12231), .b(n_10611), .o(n_12335) );
in01f80 newInst_224 ( .a(newNet_223), .o(newNet_224) );
ao12f80 g738174 ( .a(n_41878), .b(n_41995), .c(n_41901), .o(n_42021) );
in01f80 g738899 ( .a(n_41285), .o(n_41310) );
na02f80 FE_RC_1974_0 ( .a(FE_OCP_RBN1190_n_14911), .b(n_16622), .o(FE_RN_640_0) );
in01f80 g762006 ( .a(n_18935), .o(n_19733) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_7_ ( .ck(newNet_3363), .d(n_26881), .o(delay_add_ln22_unr17_stage7_stallmux_q_7_) );
na04m80 g739192 ( .a(n_40878), .b(n_40934), .c(n_41208), .d(n_40928), .o(n_40935) );
no02f80 g759670 ( .a(n_20477), .b(n_45066), .o(n_20615) );
na02f80 g745032 ( .a(n_34927), .b(n_34705), .o(n_34928) );
in01f80 g752779 ( .a(n_27434), .o(n_27433) );
oa12f80 g756089 ( .a(n_24352), .b(n_24864), .c(n_24045), .o(n_24908) );
in01f80 g759270 ( .a(n_20949), .o(n_20950) );
na02f80 g744746 ( .a(n_35223), .b(FE_OCP_RBN3650_n_35169), .o(n_35225) );
no02f80 FE_RC_1239_0 ( .a(n_8807), .b(n_8825), .o(FE_RN_372_0) );
na02f80 g762412 ( .a(FE_OCP_RBN3410_n_45120), .b(n_18420), .o(n_19400) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_25_ ( .ck(newNet_3300), .d(n_32290), .o(delay_add_ln22_unr20_stage8_stallmux_q_25_) );
na02f80 g737914 ( .a(FE_OCPN1231_n_42201), .b(n_42478), .o(n_42582) );
no02f80 g777863 ( .a(n_3166), .b(n_3141), .o(n_4336) );
na02f80 g780895 ( .a(n_374), .b(n_387), .o(n_389) );
oa22f80 FE_RC_3157_0 ( .a(n_17336), .b(n_17630), .c(n_16338), .d(n_17628), .o(n_17731) );
ao12f80 g780353 ( .a(n_901), .b(n_955), .c(n_46055), .o(n_956) );
ao12f80 g772698 ( .a(n_8052), .b(n_8197), .c(n_8122), .o(n_8255) );
ao12f80 g756436 ( .a(n_23471), .b(n_23666), .c(n_23512), .o(n_23742) );
no02f80 g771239 ( .a(n_9568), .b(n_9555), .o(n_9701) );
no02f80 FE_RC_2801_0 ( .a(FE_RN_1197_0), .b(n_9342), .o(FE_RN_1198_0) );
in01f80 g753015 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27722) );
in01f80 newInst_1168 ( .a(newNet_1167), .o(newNet_1168) );
no02f80 g749665 ( .a(n_31512), .b(n_31392), .o(n_31513) );
oa22f80 g779848 ( .a(n_44652), .b(n_1206), .c(n_44637), .d(n_1201), .o(n_1312) );
in01f80 g774137 ( .a(n_6648), .o(n_6618) );
na02f80 g741659 ( .a(n_38522), .b(n_38374), .o(n_38555) );
no02f80 g751821 ( .a(n_28230), .b(n_28229), .o(n_28231) );
oa22f80 FE_RC_1594_0 ( .a(FE_OCP_RBN2263_n_29033), .b(n_29142), .c(n_29141), .d(FE_OCP_RBN2264_n_29033), .o(n_29299) );
oa12f80 g775197 ( .a(n_5589), .b(n_5811), .c(n_5566), .o(n_5927) );
in01f80 FE_RC_2619_0 ( .a(n_40822), .o(FE_RN_1091_0) );
in01f80 g768871 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_23_), .o(n_11785) );
in01f80 FE_OCP_RBC3094_n_11475 ( .a(FE_OCP_RBN3091_n_11475), .o(FE_OCP_RBN3094_n_11475) );
na02f80 g761066 ( .a(n_19173), .b(n_18785), .o(n_19212) );
in01f80 g779825 ( .a(n_1377), .o(n_1686) );
na02f80 g747380 ( .a(n_32615), .b(n_44962), .o(n_32636) );
no02f80 g763583 ( .a(n_17575), .b(n_17574), .o(n_17611) );
in01f80 g758408 ( .a(n_23447), .o(FE_RN_1667_0) );
na02f80 g738527 ( .a(n_41582), .b(n_41545), .o(n_41622) );
ao12f80 g771022 ( .a(n_9596), .b(n_10001), .c(n_9516), .o(n_10131) );
no02f80 g778683 ( .a(n_2438), .b(FE_OFN813_n_2540), .o(n_2634) );
na02f80 g743344 ( .a(n_36731), .b(n_36750), .o(n_36765) );
in01f80 g779643 ( .a(n_1487), .o(n_1488) );
no02f80 g776445 ( .a(n_4529), .b(FE_OCP_RBN3577_n_4528), .o(n_4578) );
in01f80 g753690 ( .a(n_27201), .o(n_27202) );
no02f80 g778496 ( .a(n_2344), .b(n_1980), .o(n_2337) );
na02f80 g771458 ( .a(n_9520), .b(n_8025), .o(n_9633) );
no02f80 g759053 ( .a(n_21390), .b(n_45072), .o(n_21424) );
no02f80 g746445 ( .a(n_33382), .b(n_33380), .o(n_33424) );
in01f80 g764930 ( .a(n_15394), .o(n_15395) );
in01f80 g736911 ( .a(n_43630), .o(n_43631) );
na02f80 g772479 ( .a(n_8415), .b(n_8464), .o(n_10137) );
na02f80 g759300 ( .a(FE_OCP_RBN3676_n_21039), .b(n_21077), .o(n_21153) );
na02f80 g739752 ( .a(n_40513), .b(n_40367), .o(n_40528) );
in01f80 newInst_2802 ( .a(newNet_2801), .o(newNet_2802) );
no02f80 g773421 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n_8840) );
na02f80 g753267 ( .a(n_27110), .b(n_25889), .o(n_27256) );
no02f80 g777392 ( .a(n_3466), .b(n_3465), .o(n_3467) );
in01f80 g751516 ( .a(n_28824), .o(n_28825) );
in01f80 g752514 ( .a(n_27728), .o(n_27706) );
no02f80 g737537 ( .a(n_42529), .b(n_42470), .o(n_42530) );
no02f80 g756818 ( .a(n_24029), .b(n_23934), .o(n_24031) );
in01f80 g770781 ( .a(n_10057), .o(n_10072) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_24_ ( .ck(newNet_324), .d(n_1308), .o(delay_xor_ln22_unr3_stage2_stallmux_q_24_) );
in01f80 g746507 ( .a(n_33221), .o(n_33222) );
in01f80 g776715 ( .a(n_4160), .o(n_5529) );
in01f80 g775493 ( .a(n_5684), .o(n_5685) );
oa22f80 FE_RC_1456_0 ( .a(n_32287), .b(n_32338), .c(n_28336), .d(n_44432), .o(n_32373) );
no02f80 g760751 ( .a(n_20138), .b(n_19649), .o(n_20181) );
na02f80 g749657 ( .a(n_30154), .b(n_30012), .o(n_30155) );
in01f80 newInst_2142 ( .a(newNet_1222), .o(newNet_2142) );
na02f80 g761058 ( .a(n_19248), .b(n_19212), .o(n_19342) );
no02f80 g771227 ( .a(n_9658), .b(n_9404), .o(n_9739) );
no02f80 g780770 ( .a(n_558), .b(n_557), .o(n_559) );
no02f80 g743098 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n_37093) );
in01f80 g775813 ( .a(n_5420), .o(n_5421) );
in01f80 newInst_3049 ( .a(newNet_903), .o(newNet_3049) );
na02f80 g737038 ( .a(n_43046), .b(n_42598), .o(n_43144) );
no02f80 g780870 ( .a(n_354), .b(beta_3), .o(n_360) );
na02f80 g749828 ( .a(FE_OCP_RBN3016_n_31117), .b(n_31253), .o(n_31572) );
na02f80 g767682 ( .a(n_13213), .b(n_13099), .o(n_13172) );
in01f80 g748906 ( .a(n_32391), .o(n_32447) );
in01f80 newInst_1166 ( .a(newNet_1165), .o(newNet_1166) );
no02f80 g771054 ( .a(n_9417), .b(n_8362), .o(n_9582) );
in01f80 g753634 ( .a(n_26628), .o(n_26629) );
na02f80 g759641 ( .a(n_20616), .b(n_20302), .o(n_20684) );
na02f80 g754854 ( .a(n_25624), .b(n_25625), .o(n_25650) );
oa12f80 g738355 ( .a(n_41521), .b(n_41551), .c(n_41520), .o(n_42241) );
in01f80 FE_OCP_DRV_C3168_FE_RN_1789_0 ( .a(FE_OCP_DRV_N3167_FE_RN_1789_0), .o(FE_OCP_DRV_N3168_FE_RN_1789_0) );
no02f80 g777111 ( .a(n_3929), .b(FE_OCP_RBN2582_n_3734), .o(n_3959) );
in01f80 g770019 ( .a(n_10910), .o(n_10935) );
in01f80 g780119 ( .a(n_1211), .o(n_1204) );
in01f80 FE_OCPC1022_n_23195 ( .a(FE_OCPN1021_n_23195), .o(FE_OCPN1022_n_23195) );
in01f80 g750436 ( .a(n_29609), .o(n_29610) );
in01f80 FE_OCP_RBC2579_n_3734 ( .a(n_3734), .o(FE_OCP_RBN2579_n_3734) );
in01f80 g773452 ( .a(n_7925), .o(n_7900) );
in01f80 newInst_1583 ( .a(newNet_1433), .o(newNet_1583) );
in01f80 g737068 ( .a(n_43165), .o(n_43214) );
no02f80 g776150 ( .a(n_4914), .b(n_4941), .o(n_5110) );
no02f80 g764112 ( .a(n_16588), .b(FE_OCP_RBN2697_n_14814), .o(n_16603) );
na02f80 g770828 ( .a(n_9931), .b(n_10016), .o(n_10032) );
na02f80 g771253 ( .a(n_9457), .b(n_9453), .o(n_9623) );
in01f80 g769894 ( .a(n_11052), .o(n_11029) );
ao22s80 g742692 ( .a(n_37379), .b(n_37123), .c(n_37317), .d(n_37122), .o(n_37411) );
oa12f80 g769117 ( .a(n_11424), .b(n_11582), .c(n_11581), .o(n_11652) );
ao12f80 g781096 ( .a(n_105), .b(n_245), .c(n_155), .o(n_255) );
ao12f80 g761636 ( .a(n_18940), .b(n_18887), .c(n_18822), .o(n_18971) );
in01f80 g760839 ( .a(n_19441), .o(n_19442) );
no02f80 g751455 ( .a(n_28574), .b(n_28605), .o(n_28628) );
no02f80 g747749 ( .a(n_33496), .b(n_33461), .o(n_33800) );
na02f80 g740182 ( .a(FE_OCP_RBN3715_n_39913), .b(n_39945), .o(n_40073) );
in01f80 g779353 ( .a(n_1787), .o(n_1648) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_22_ ( .ck(newNet_2554), .d(n_27693), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_) );
in01f80 FE_OCP_RBC1924_cordic_combinational_sub_ln23_0_unr12_z_0__ ( .a(FE_OCP_RBN1922_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__) );
na02f80 g765590 ( .a(n_15366), .b(n_15397), .o(n_15748) );
in01f80 newInst_1988 ( .a(newNet_1987), .o(newNet_1988) );
in01f80 FE_RC_3569_0 ( .a(n_24462), .o(FE_RN_1551_0) );
na02f80 g740522 ( .a(n_39690), .b(FE_OCP_RBN2945_FE_RN_1269_0), .o(n_39711) );
in01f80 g770798 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .o(n_10387) );
in01f80 FE_OCP_RBC3045_n_5881 ( .a(n_5881), .o(FE_OCP_RBN3045_n_5881) );
na02f80 g737009 ( .a(FE_OCP_RBN3073_n_43230), .b(n_42991), .o(n_43429) );
na02f80 g774938 ( .a(n_6110), .b(n_6104), .o(n_6176) );
ao22s80 g736354 ( .a(n_43840), .b(n_43600), .c(n_43841), .d(n_43599), .o(n_43868) );
in01f80 g762865 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n_17700) );
ao22s80 g762048 ( .a(FE_OCP_RBN2205_n_18242), .b(n_18331), .c(n_18355), .d(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n_18537) );
in01f80 g749086 ( .a(n_31048), .o(n_31049) );
no02f80 FE_RC_3689_0 ( .a(n_12395), .b(FE_RN_1621_0), .o(n_12463) );
na02f80 g746689 ( .a(n_34277), .b(n_33816), .o(n_34390) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_3_ ( .ck(newNet_1006), .d(n_16789), .o(delay_xor_ln21_unr12_stage5_stallmux_q_3_) );
no02f80 g760786 ( .a(n_19626), .b(n_19625), .o(n_19627) );
no02f80 g755533 ( .a(n_24638), .b(n_22207), .o(n_24685) );
na02f80 g749851 ( .a(FE_OCP_RBN3013_n_31117), .b(n_30417), .o(n_31222) );
in01f80 g746551 ( .a(n_34803), .o(n_34804) );
in01f80 newInst_3228 ( .a(newNet_1021), .o(newNet_3228) );
oa12f80 g781144 ( .a(n_127), .b(n_208), .c(n_92), .o(n_211) );
na02f80 g749972 ( .a(n_30196), .b(n_30113), .o(n_30220) );
in01f80 g780656 ( .a(n_779), .o(n_890) );
in01f80 g752692 ( .a(n_28082), .o(n_28136) );
na02f80 g770129 ( .a(n_10810), .b(FE_OCP_RBN3637_n_44490), .o(n_10897) );
na02f80 g761018 ( .a(n_19264), .b(FE_OFN780_n_17093), .o(n_19321) );
in01f80 g757945 ( .a(n_22235), .o(n_22314) );
in01f80 g779416 ( .a(n_1495), .o(n_1496) );
no02f80 g763816 ( .a(n_16853), .b(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n_16854) );
in01f80 newInst_3133 ( .a(newNet_706), .o(newNet_3133) );
no02f80 g757080 ( .a(n_23549), .b(n_23548), .o(n_23550) );
in01f80 g772558 ( .a(n_8428), .o(n_8429) );
in01f80 g736679 ( .a(n_43075), .o(n_43095) );
in01f80 newInst_1701 ( .a(newNet_1700), .o(newNet_1701) );
oa12f80 g738216 ( .a(n_41945), .b(n_41944), .c(n_41943), .o(n_41983) );
no02f80 g744725 ( .a(n_35204), .b(n_35133), .o(n_35253) );
in01f80 FE_OCP_RBC3599_FE_OCPN1243_n_44460 ( .a(FE_OCP_RBN3598_FE_OCPN1243_n_44460), .o(FE_OCP_RBN3599_FE_OCPN1243_n_44460) );
na02f80 g739373 ( .a(n_40823), .b(n_40719), .o(n_41282) );
in01f80 newInst_3578 ( .a(newNet_3577), .o(newNet_3578) );
na02f80 g763751 ( .a(n_46978), .b(FE_OCP_RBN2735_n_14985), .o(n_16706) );
in01f80 g738357 ( .a(n_41476), .o(n_41477) );
in01f80 g769596 ( .a(n_11337), .o(n_11479) );
in01f80 newInst_3088 ( .a(newNet_2319), .o(newNet_3088) );
na02f80 g753561 ( .a(n_26674), .b(n_26705), .o(n_26675) );
na02f80 g756399 ( .a(n_24259), .b(n_24240), .o(n_24241) );
in01f80 g778014 ( .a(n_4719), .o(n_3113) );
na02f80 g738708 ( .a(n_41435), .b(n_41122), .o(n_41577) );
in01f80 g758757 ( .a(n_21682), .o(n_21683) );
no02f80 g771397 ( .a(n_9643), .b(n_9642), .o(n_9787) );
in01f80 newInst_2187 ( .a(newNet_2186), .o(newNet_2187) );
na02f80 g775287 ( .a(n_5656), .b(n_4875), .o(n_5669) );
in01f80 g774144 ( .a(n_6866), .o(n_6867) );
in01f80 g745726 ( .a(n_35451), .o(n_35452) );
na02f80 g776223 ( .a(n_4706), .b(n_4699), .o(n_4734) );
in01f80 fopt783993 ( .a(n_45717), .o(n_45716) );
na02f80 g738485 ( .a(n_41381), .b(n_41406), .o(n_41391) );
in01f80 newInst_3264 ( .a(newNet_3263), .o(newNet_3264) );
no02f80 g741028 ( .a(n_39028), .b(n_39004), .o(n_39079) );
oa22f80 FE_RC_3253_0 ( .a(n_11501), .b(n_11553), .c(FE_RN_1435_0), .d(n_11523), .o(n_11778) );
oa22f80 FE_RC_1628_0 ( .a(n_6443), .b(n_6554), .c(n_6442), .d(n_6572), .o(n_6739) );
in01f80 FE_OCP_RBC3211_n_44365 ( .a(FE_OCP_RBN3213_n_44365), .o(FE_OCP_RBN3211_n_44365) );
in01f80 FE_RC_3638_0 ( .a(n_30224), .o(FE_RN_1596_0) );
na02f80 g770271 ( .a(n_10690), .b(n_10724), .o(n_10772) );
in01f80 FE_OCP_RBC2838_n_4692 ( .a(n_4692), .o(FE_OCP_RBN2838_n_4692) );
in01f80 FE_OCP_RBC2366_n_24372 ( .a(n_24372), .o(FE_OCP_RBN2366_n_24372) );
no02f80 g759779 ( .a(n_21697), .b(n_21450), .o(n_21715) );
no02f80 g752301 ( .a(FE_OCP_RBN2180_FE_RN_526_0), .b(n_28155), .o(n_28539) );
na02f80 g751982 ( .a(n_28782), .b(n_27958), .o(n_28811) );
ao22s80 FE_RC_242_0 ( .a(n_13515), .b(n_14328), .c(n_14327), .d(FE_OCP_RBN2252_n_13017), .o(n_14462) );
in01f80 newInst_233 ( .a(newNet_100), .o(newNet_233) );
in01f80 g759162 ( .a(n_21093), .o(n_21143) );
no02f80 g754502 ( .a(n_25513), .b(n_25232), .o(n_25601) );
na02f80 g764639 ( .a(n_15986), .b(n_15943), .o(n_16144) );
in01f80 g768008 ( .a(n_12683), .o(n_12635) );
in01f80 FE_OCP_RBC1327_n_36489 ( .a(FE_OCP_RBN1326_n_36489), .o(FE_OCP_RBN1327_n_36489) );
no02f80 g747827 ( .a(n_33392), .b(n_33437), .o(n_33461) );
no02f80 g770899 ( .a(n_9904), .b(n_8562), .o(n_9978) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_13_ ( .ck(newNet_1343), .d(n_1187), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_) );
oa22f80 g744203 ( .a(FE_OCPN1510_n_44174), .b(n_34899), .c(n_44180), .d(FE_OCPN1422_n_35611), .o(n_36291) );
in01f80 g780323 ( .a(n_45816), .o(n_863) );
oa22f80 FE_RC_4106_0 ( .a(n_22377), .b(n_22687), .c(n_22378), .d(n_22721), .o(n_22875) );
no02f80 g760935 ( .a(n_19454), .b(n_20523), .o(n_19455) );
na02f80 g738514 ( .a(n_41540), .b(n_41698), .o(n_41679) );
in01f80 newInst_1678 ( .a(newNet_617), .o(newNet_1678) );
no02f80 g747298 ( .a(n_32770), .b(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n_32751) );
in01f80 g775012 ( .a(n_6162), .o(n_6163) );
no02f80 g749263 ( .a(n_30678), .b(n_30403), .o(n_30712) );
in01f80 g756467 ( .a(n_23689), .o(n_23690) );
na02f80 g754151 ( .a(FE_OCP_RBN2815_n_25986), .b(n_23353), .o(n_26053) );
no02f80 g766954 ( .a(n_13903), .b(n_13902), .o(n_14083) );
in01f80 g759536 ( .a(n_20907), .o(n_20908) );
in01f80 newInst_3613 ( .a(newNet_1905), .o(newNet_3613) );
in01f80 g761129 ( .a(n_19238), .o(n_20343) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_31_ ( .ck(newNet_3199), .d(n_36629), .o(delay_add_ln22_unr23_stage9_stallmux_q_31_) );
oa12f80 g738930 ( .a(n_41245), .b(n_41244), .c(n_41243), .o(n_41628) );
na02f80 g766037 ( .a(n_14760), .b(n_14781), .o(n_14915) );
na02f80 g766554 ( .a(n_14049), .b(n_14141), .o(n_14222) );
in01f80 newInst_1633 ( .a(newNet_1632), .o(newNet_1633) );
na02f80 g775414 ( .a(n_5543), .b(n_4182), .o(n_5558) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_1_ ( .ck(newNet_419), .d(n_32467), .o(delay_xor_ln22_unr21_stage8_stallmux_q_1_) );
in01f80 FE_OCP_RBC1352_n_19148 ( .a(FE_OCP_RBN1351_n_19148), .o(FE_OCP_RBN1352_n_19148) );
na02f80 g742122 ( .a(n_37862), .b(n_37275), .o(n_38073) );
in01f80 newInst_1278 ( .a(newNet_1277), .o(newNet_1278) );
na02f80 g775657 ( .a(n_5215), .b(n_4556), .o(n_5358) );
oa12f80 g770254 ( .a(n_10753), .b(n_10752), .c(n_10751), .o(n_10815) );
no02f80 g768470 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_20_), .o(n_12400) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_27_ ( .ck(newNet_1386), .d(n_36729), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_) );
in01f80 fopt783329 ( .a(n_44877), .o(n_44875) );
in01f80 g757271 ( .a(n_23045), .o(n_23046) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_1_ ( .ck(newNet_2954), .d(n_4491), .o(delay_add_ln22_unr5_stage3_stallmux_q_1_) );
na02f80 g742951 ( .a(n_37103), .b(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37183) );
no03m80 g754960 ( .a(n_25693), .b(n_25750), .c(n_25749), .o(n_25751) );
in01f80 FE_OCPC1394_n_962 ( .a(FE_OCPN1393_n_962), .o(FE_OCPN1394_n_962) );
na02f80 g741859 ( .a(n_38434), .b(n_38432), .o(n_38433) );
no02f80 g770327 ( .a(FE_OCP_RBN2869_n_10480), .b(n_44463), .o(n_10520) );
na02f80 g746444 ( .a(n_33277), .b(n_33274), .o(n_33351) );
na02f80 g760158 ( .a(n_20537), .b(n_20528), .o(n_20529) );
no02f80 g748167 ( .a(n_31706), .b(n_31680), .o(n_31743) );
in01f80 g745434 ( .a(n_34326), .o(n_34386) );
oa12f80 g770294 ( .a(n_9915), .b(n_10720), .c(n_9824), .o(n_10817) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_7_ ( .ck(newNet_2141), .d(n_1004), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_) );
in01f80 newInst_1124 ( .a(newNet_1123), .o(newNet_1124) );
no02f80 g775718 ( .a(n_5255), .b(n_4556), .o(n_5313) );
na02f80 g744290 ( .a(n_44180), .b(FE_OCP_RBN2645_n_34980), .o(n_35857) );
na02f80 g742367 ( .a(n_37791), .b(n_37240), .o(n_37815) );
no02f80 g756587 ( .a(n_23606), .b(n_23605), .o(n_23607) );
in01f80 FE_OCP_RBC3693_n_10852 ( .a(n_10852), .o(FE_OCP_RBN3693_n_10852) );
in01f80 g737497 ( .a(n_42635), .o(n_42636) );
na02f80 g739466 ( .a(FE_OCPN898_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .o(n_41077) );
no02f80 g780919 ( .a(n_521), .b(n_549), .o(n_560) );
na02f80 FE_RC_2808_0 ( .a(FE_RN_1201_0), .b(FE_OCP_RBN2348_n_13702), .o(n_13788) );
no02f80 g760580 ( .a(n_19836), .b(n_19887), .o(n_19948) );
na02f80 g776462 ( .a(n_4502), .b(n_4230), .o(n_4661) );
in01f80 g757487 ( .a(n_22959), .o(n_23226) );
in01f80 g768563 ( .a(n_12325), .o(n_12326) );
in01f80 g741456 ( .a(n_38811), .o(n_38812) );
in01f80 newInst_1780 ( .a(newNet_597), .o(newNet_1780) );
in01f80 newInst_2326 ( .a(newNet_2325), .o(newNet_2326) );
in01f80 newInst_1766 ( .a(newNet_1765), .o(newNet_1766) );
in01f80 g738073 ( .a(n_42459), .o(n_42483) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_15_ ( .ck(newNet_1638), .d(n_27134), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_) );
in01f80 newInst_2199 ( .a(newNet_2198), .o(newNet_2199) );
in01f80 newInst_2992 ( .a(newNet_2991), .o(newNet_2992) );
ao12f80 g756352 ( .a(n_23955), .b(n_24417), .c(n_24215), .o(n_24455) );
na02f80 g763738 ( .a(n_17428), .b(n_17468), .o(n_18234) );
in01f80 newInst_1694 ( .a(newNet_1693), .o(newNet_1694) );
no02f80 g758059 ( .a(n_22760), .b(n_22839), .o(n_23526) );
no02f80 g750258 ( .a(n_30840), .b(n_30232), .o(n_30895) );
in01f80 g752770 ( .a(n_28152), .o(n_28153) );
no02f80 g737508 ( .a(n_42498), .b(n_42497), .o(n_42538) );
no02f80 g741007 ( .a(n_39102), .b(n_39157), .o(n_39253) );
no02f80 FE_RC_127_0 ( .a(FE_RN_30_0), .b(FE_RN_31_0), .o(FE_RN_32_0) );
in01f80 newInst_2664 ( .a(newNet_2663), .o(newNet_2664) );
in01f80 FE_OFC838_n_4632 ( .a(n_4632), .o(FE_OFN838_n_4632) );
in01f80 g761825 ( .a(n_19191), .o(n_19158) );
ao12f80 g743473 ( .a(n_37676), .b(n_37713), .c(n_46238), .o(n_37750) );
ao12f80 g747973 ( .a(n_33044), .b(n_33043), .c(n_33042), .o(n_33438) );
no02f80 FE_RC_2985_0 ( .a(FE_RN_1302_0), .b(n_10828), .o(FE_RN_1303_0) );
in01f80 newInst_1597 ( .a(newNet_1596), .o(newNet_1597) );
in01f80 newInst_3504 ( .a(newNet_3503), .o(newNet_3504) );
no02f80 g745744 ( .a(n_34128), .b(n_34127), .o(n_34129) );
na02f80 FE_RC_2832_0 ( .a(FE_RN_1217_0), .b(n_24285), .o(n_24307) );
in01f80 g746814 ( .a(n_33303), .o(n_33304) );
na02f80 g770931 ( .a(n_10131), .b(n_10086), .o(n_10087) );
ao12f80 g746763 ( .a(n_33108), .b(n_33199), .c(n_32336), .o(n_33202) );
in01f80 newInst_362 ( .a(newNet_361), .o(newNet_362) );
no02f80 FE_RC_2581_0 ( .a(FE_RN_1063_0), .b(FE_RN_1064_0), .o(FE_RN_1065_0) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_30_ ( .ck(newNet_2448), .d(n_32519), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_) );
ao12f80 g738604 ( .a(n_41724), .b(n_41716), .c(n_41339), .o(n_42056) );
in01f80 g758897 ( .a(n_21473), .o(n_21474) );
oa12f80 g746632 ( .a(n_33760), .b(n_34300), .c(n_33703), .o(n_34442) );
no02f80 g744056 ( .a(n_44222), .b(n_35785), .o(n_36331) );
in01f80 newInst_3729 ( .a(newNet_1271), .o(newNet_3729) );
na02f80 g770693 ( .a(n_10375), .b(n_10374), .o(n_10489) );
no02f80 g769901 ( .a(n_11045), .b(n_10989), .o(n_11080) );
no02f80 g748421 ( .a(n_31518), .b(n_46958), .o(n_31704) );
in01f80 g747633 ( .a(n_32219), .o(n_32220) );
na02f80 g771365 ( .a(n_9188), .b(n_8232), .o(n_9254) );
no02f80 g742153 ( .a(n_38131), .b(n_38079), .o(n_38153) );
oa22f80 g779852 ( .a(n_44652), .b(n_1025), .c(n_44623), .d(n_989), .o(n_1300) );
no02f80 g744004 ( .a(n_36192), .b(n_36097), .o(n_36193) );
in01f80 g745184 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_36354) );
na02f80 g773021 ( .a(n_7704), .b(n_7729), .o(n_7820) );
ao22s80 FE_RC_3238_0 ( .a(n_9170), .b(n_9293), .c(n_9242), .d(n_9215), .o(n_9494) );
in01f80 g749173 ( .a(n_32227), .o(n_32245) );
na02f80 g737319 ( .a(n_42840), .b(n_42408), .o(n_42873) );
in01f80 g781177 ( .a(n_368), .o(n_372) );
in01f80 newInst_2847 ( .a(newNet_2367), .o(newNet_2847) );
in01f80 g759196 ( .a(n_22156), .o(n_21413) );
no02f80 g759183 ( .a(n_21384), .b(FE_OCPN1524_n_45072), .o(n_21463) );
ao12f80 g756440 ( .a(n_23606), .b(n_23761), .c(n_23773), .o(n_23774) );
no02f80 g748261 ( .a(n_31835), .b(FE_OCP_RBN2804_n_30534), .o(n_31846) );
no02f80 g781318 ( .a(beta_29), .b(beta_31), .o(n_56) );
in01f80 g747833 ( .a(n_33667), .o(n_33668) );
na02f80 g740545 ( .a(n_39657), .b(n_39616), .o(n_39677) );
in01f80 g751460 ( .a(n_28679), .o(n_28680) );
in01f80 newInst_1911 ( .a(newNet_1910), .o(newNet_1911) );
in01f80 FE_RC_2058_0 ( .a(n_24823), .o(FE_RN_697_0) );
no02f80 g767292 ( .a(n_13535), .b(n_13489), .o(n_13537) );
no02f80 g764236 ( .a(n_16446), .b(n_16199), .o(n_16495) );
in01f80 g778922 ( .a(n_2191), .o(n_2225) );
in01f80 g765483 ( .a(n_15108), .o(n_15109) );
in01f80 g780517 ( .a(n_1070), .o(n_1071) );
in01f80 g755186 ( .a(n_25715), .o(n_25688) );
na02f80 FE_RC_2610_0 ( .a(FE_RN_1085_0), .b(n_18096), .o(n_18113) );
in01f80 g739686 ( .a(n_40536), .o(n_40537) );
na02f80 g762928 ( .a(n_17990), .b(n_17989), .o(n_17991) );
in01f80 g773208 ( .a(n_7815), .o(n_7816) );
na02f80 g771605 ( .a(n_9238), .b(n_9265), .o(n_9365) );
no02f80 FE_RC_2288_0 ( .a(FE_RN_857_0), .b(n_17734), .o(FE_RN_858_0) );
na02f80 g759455 ( .a(FE_OCP_RBN1842_n_20910), .b(FE_RN_1585_0), .o(n_20968) );
no02f80 g750501 ( .a(n_29485), .b(FE_OCPN1406_n_25859), .o(n_29486) );
in01f80 g773055 ( .a(FE_OCPN915_n_7832), .o(n_8752) );
in01f80 g740963 ( .a(n_39194), .o(n_39195) );
in01f80 g763230 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(n_17394) );
in01f80 newInst_227 ( .a(newNet_226), .o(newNet_227) );
oa22f80 g771729 ( .a(n_8720), .b(n_8859), .c(n_8719), .d(n_8836), .o(n_9009) );
na02f80 FE_RC_2598_0 ( .a(n_2913), .b(FE_RN_1076_0), .o(FE_RN_1077_0) );
no02f80 g772758 ( .a(n_8134), .b(n_8078), .o(n_8213) );
na02f80 g777345 ( .a(n_4675), .b(n_5165), .o(n_5387) );
no02f80 g742821 ( .a(n_37243), .b(n_37242), .o(n_37244) );
oa22f80 g781280 ( .a(n_77), .b(n_46055), .c(n_7), .d(beta_8), .o(n_188) );
no02f80 g751583 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n_28608) );
in01f80 g765264 ( .a(n_15523), .o(n_15524) );
na02f80 g779237 ( .a(n_1796), .b(n_1666), .o(n_1847) );
in01f80 newInst_3148 ( .a(newNet_3147), .o(newNet_3148) );
no02f80 g769940 ( .a(n_11059), .b(n_9620), .o(n_11158) );
na02f80 g738917 ( .a(n_41270), .b(n_41269), .o(n_41271) );
na02f80 g736996 ( .a(n_43097), .b(n_42989), .o(n_43187) );
no02f80 g778429 ( .a(n_2734), .b(n_2657), .o(n_2764) );
in01f80 FE_OCP_RBC3217_n_19781 ( .a(n_19781), .o(FE_OCP_RBN3217_n_19781) );
na03f80 FE_RC_2247_0 ( .a(FE_RN_824_0), .b(n_37157), .c(FE_RN_825_0), .o(FE_RN_826_0) );
in01f80 g767037 ( .a(n_13900), .o(n_13901) );
ao12f80 g741854 ( .a(n_38284), .b(n_38286), .c(n_38271), .o(n_38391) );
in01f80 g774482 ( .a(n_6569), .o(n_6621) );
in01f80 g739688 ( .a(n_40534), .o(n_40535) );
no02f80 g764454 ( .a(n_16123), .b(n_16082), .o(n_16161) );
no02f80 g769183 ( .a(n_12080), .b(n_12079), .o(n_12081) );
oa12f80 g781101 ( .a(n_70), .b(n_244), .c(n_135), .o(n_247) );
na02f80 g750534 ( .a(n_29478), .b(n_29454), .o(n_29574) );
in01f80 g746845 ( .a(n_33262), .o(n_33263) );
na02f80 g745449 ( .a(n_34436), .b(n_34307), .o(n_34437) );
in01f80 g739271 ( .a(n_40929), .o(n_40930) );
na02f80 g768358 ( .a(n_12427), .b(n_12363), .o(n_12466) );
na02f80 g761257 ( .a(n_18952), .b(n_18512), .o(n_18989) );
na02f80 g746320 ( .a(n_33613), .b(n_33534), .o(n_33614) );
na02f80 g742251 ( .a(n_37853), .b(n_37845), .o(n_37846) );
no02f80 g747619 ( .a(n_32223), .b(n_32197), .o(n_32198) );
na02f80 g767474 ( .a(n_13462), .b(n_12999), .o(n_13505) );
na02f80 g765148 ( .a(n_15343), .b(FE_OCP_DRV_N3156_n_15342), .o(n_15460) );
na02f80 g759358 ( .a(n_21069), .b(n_20665), .o(n_21071) );
na02f80 g754569 ( .a(n_26898), .b(n_26897), .o(n_26928) );
oa12f80 g767325 ( .a(n_12914), .b(n_13407), .c(n_13453), .o(n_13535) );
no02f80 g763025 ( .a(n_17939), .b(n_17471), .o(n_17959) );
no02f80 g774340 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_13_), .o(n_6951) );
oa22f80 g749112 ( .a(n_32158), .b(n_31315), .c(n_32176), .d(n_31316), .o(n_32248) );
na02f80 g741906 ( .a(n_38126), .b(n_38125), .o(n_38127) );
na02f80 g777126 ( .a(n_3575), .b(n_3460), .o(n_3683) );
ao22s80 g778904 ( .a(n_2305), .b(n_2020), .c(n_2279), .d(n_2019), .o(n_2387) );
no02f80 g744628 ( .a(n_36603), .b(n_36084), .o(n_36621) );
no02f80 g778630 ( .a(n_2741), .b(n_2752), .o(n_2900) );
no02f80 g776703 ( .a(n_4310), .b(n_4256), .o(n_4368) );
in01f80 FE_RC_4218_0 ( .a(n_29896), .o(FE_RN_1847_0) );
na02f80 g779370 ( .a(n_1572), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_), .o(n_1657) );
na02f80 g758593 ( .a(n_21850), .b(n_21616), .o(n_21923) );
na02f80 g752390 ( .a(n_44763), .b(delay_xor_ln22_unr18_stage7_stallmux_q_1_), .o(n_27738) );
ao12f80 g778992 ( .a(n_2165), .b(n_2172), .c(n_2164), .o(n_2197) );
na02f80 g754690 ( .a(n_26856), .b(n_26679), .o(n_26897) );
in01f80 newInst_1053 ( .a(newNet_1052), .o(newNet_1053) );
in01f80 g768124 ( .a(n_12731), .o(n_12732) );
oa22f80 g753573 ( .a(n_27320), .b(n_26928), .c(n_27319), .d(n_26929), .o(n_27447) );
in01f80 g781009 ( .a(n_465), .o(n_274) );
no02f80 g767765 ( .a(n_13069), .b(n_12188), .o(n_13377) );
na02f80 g771525 ( .a(n_9470), .b(n_9387), .o(n_9471) );
in01f80 g771168 ( .a(n_9840), .o(n_9841) );
ao12f80 g739389 ( .a(n_40770), .b(FE_OCPN897_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n_41269) );
in01f80 g755527 ( .a(n_24581), .o(n_24582) );
in01f80 g763507 ( .a(n_16903), .o(n_16944) );
na02f80 FE_RC_531_0 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .b(FE_OCP_RBN3822_n_44061), .o(FE_RN_165_0) );
in01f80 newInst_2357 ( .a(newNet_330), .o(newNet_2357) );
na02f80 g764772 ( .a(n_15628), .b(n_15658), .o(n_15765) );
na02f80 g741518 ( .a(n_38703), .b(n_38697), .o(n_38733) );
na02f80 g748438 ( .a(n_31469), .b(n_31519), .o(n_31550) );
oa12f80 g763218 ( .a(n_16809), .b(n_16884), .c(n_16760), .o(n_17009) );
in01f80 newInst_2037 ( .a(newNet_2036), .o(newNet_2037) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_6_ ( .ck(newNet_3189), .d(n_35705), .o(delay_add_ln22_unr23_stage9_stallmux_q_6_) );
in01f80 FE_OCP_RBC3009_n_31117 ( .a(FE_OCP_RBN3701_n_31064), .o(FE_OCP_RBN3009_n_31117) );
ao12f80 g740912 ( .a(n_39339), .b(n_39338), .c(n_39337), .o(n_39808) );
na02f80 g747716 ( .a(n_32088), .b(n_31683), .o(n_32090) );
na02f80 g780606 ( .a(n_890), .b(n_905), .o(n_1053) );
na02f80 g741050 ( .a(n_38921), .b(n_38964), .o(n_38965) );
in01f80 newInst_3650 ( .a(newNet_3649), .o(newNet_3650) );
na02f80 g773811 ( .a(n_7091), .b(delay_add_ln22_unr5_stage3_stallmux_q_12_), .o(n_7147) );
in01f80 g754474 ( .a(n_25598), .o(n_25599) );
ms00f80 cos_out_reg_15_ ( .ck(newNet_3743), .d(n_43850), .o(cos_out_15) );
in01f80 g759679 ( .a(n_21796), .o(n_21797) );
oa22f80 g757703 ( .a(n_22513), .b(n_22312), .c(n_22543), .d(n_22346), .o(n_22635) );
na02f80 FE_RC_192_0 ( .a(FE_RN_65_0), .b(n_13851), .o(n_46984) );
no02f80 g775261 ( .a(n_5653), .b(n_5670), .o(n_5802) );
no02f80 g778721 ( .a(n_2365), .b(n_2357), .o(n_2390) );
in01f80 g754974 ( .a(n_25149), .o(n_25150) );
no02f80 g744304 ( .a(FE_OCP_RBN2903_n_44174), .b(n_35194), .o(n_36030) );
in01f80 g759730 ( .a(n_20420), .o(n_20443) );
no02f80 g740335 ( .a(n_40308), .b(n_40241), .o(n_40355) );
in01f80 FE_OCP_RBC1844_n_20910 ( .a(FE_OCP_RBN1843_n_20910), .o(FE_OCP_RBN1844_n_20910) );
no02f80 g776016 ( .a(n_5021), .b(n_4998), .o(n_5022) );
in01f80 g762405 ( .a(n_18655), .o(n_18728) );
oa22f80 g758704 ( .a(n_22247), .b(n_21716), .c(n_22248), .d(n_21715), .o(n_22361) );
in01f80 g750652 ( .a(n_29347), .o(n_29348) );
oa12f80 g736257 ( .a(n_293), .b(n_43908), .c(FE_OFN4_n_43918), .o(n_43917) );
no02f80 g746250 ( .a(n_33642), .b(n_47249), .o(n_33643) );
in01f80 FE_OCP_RBC3409_n_45120 ( .a(n_45120), .o(FE_OCP_RBN3409_n_45120) );
in01f80 g762034 ( .a(n_18591), .o(n_18592) );
na02f80 g747620 ( .a(n_32191), .b(n_31841), .o(n_32241) );
in01f80 newInst_3519 ( .a(newNet_3518), .o(newNet_3519) );
no02f80 g767274 ( .a(n_13716), .b(n_13700), .o(n_13701) );
no02f80 g740220 ( .a(n_39970), .b(FE_OCP_RBN3021_n_39942), .o(n_40107) );
in01f80 newInst_110 ( .a(newNet_109), .o(newNet_110) );
oa22f80 FE_RC_3263_0 ( .a(n_9306), .b(n_9229), .c(n_9230), .d(n_9307), .o(n_9506) );
na02f80 g749788 ( .a(n_31394), .b(n_31254), .o(n_31315) );
in01f80 FE_OCP_RBC3029_n_39942 ( .a(FE_OCP_RBN3025_n_39942), .o(FE_OCP_RBN3029_n_39942) );
na02f80 g771125 ( .a(n_47259), .b(n_9447), .o(n_9542) );
oa12f80 g770429 ( .a(n_9773), .b(n_10551), .c(n_9776), .o(n_10689) );
oa12f80 g738864 ( .a(n_41274), .b(n_41273), .c(n_41272), .o(n_41656) );
in01f80 g736284 ( .a(n_43892), .o(n_43893) );
in01f80 newInst_1555 ( .a(newNet_487), .o(newNet_1555) );
in01f80 newInst_3715 ( .a(newNet_3714), .o(newNet_3715) );
in01f80 g739835 ( .a(n_40446), .o(n_40447) );
na02f80 g743969 ( .a(n_35784), .b(n_35824), .o(n_35825) );
in01f80 g756907 ( .a(n_23420), .o(n_23386) );
na02f80 g751559 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_19_), .o(n_28520) );
no02f80 g777915 ( .a(n_3149), .b(n_2983), .o(n_3150) );
no02f80 g736340 ( .a(n_43788), .b(n_43468), .o(n_43816) );
na02f80 g776244 ( .a(n_4320), .b(n_4175), .o(n_4462) );
ao12f80 g773691 ( .a(n_7334), .b(n_7335), .c(n_7333), .o(n_7611) );
na02f80 g745065 ( .a(n_34855), .b(n_34854), .o(n_34856) );
in01f80 g736532 ( .a(n_43709), .o(n_43710) );
in01f80 g740597 ( .a(n_39616), .o(n_39621) );
in01f80 newInst_1816 ( .a(newNet_1274), .o(newNet_1816) );
na02f80 g740773 ( .a(n_39512), .b(n_39492), .o(n_39905) );
in01f80 newInst_2275 ( .a(newNet_2274), .o(newNet_2275) );
na02f80 g759728 ( .a(n_47174), .b(n_20348), .o(n_20477) );
in01f80 g736787 ( .a(n_43558), .o(n_43559) );
in01f80 newInst_679 ( .a(newNet_396), .o(newNet_679) );
no02f80 g774709 ( .a(n_6373), .b(n_6244), .o(n_6374) );
na02f80 g738418 ( .a(n_41696), .b(n_41695), .o(n_41697) );
in01f80 g755114 ( .a(n_25352), .o(n_25416) );
oa12f80 g765581 ( .a(n_14526), .b(n_15481), .c(n_14528), .o(n_15576) );
no02f80 g755800 ( .a(n_24267), .b(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24296) );
in01f80 FE_OCP_RBC3712_n_31466 ( .a(n_31466), .o(FE_OCP_RBN3712_n_31466) );
oa12f80 g758323 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n_23087) );
in01f80 FE_OCP_RBC2294_n_2438 ( .a(FE_OCP_RBN2290_n_2438), .o(FE_OCP_RBN2294_n_2438) );
ao12f80 g764117 ( .a(n_16524), .b(n_16552), .c(n_16580), .o(n_16624) );
na02f80 g766104 ( .a(n_14552), .b(FE_OCP_RBN2449_n_14114), .o(n_14583) );
in01f80 g778365 ( .a(n_2809), .o(n_2810) );
in01f80 g742041 ( .a(n_38214), .o(n_38215) );
in01f80 newInst_2506 ( .a(newNet_2505), .o(newNet_2506) );
na02f80 g778139 ( .a(n_2908), .b(n_2963), .o(n_2967) );
in01f80 g781337 ( .a(n_91), .o(n_92) );
no02f80 g743428 ( .a(n_44809), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36687) );
ao12f80 g741093 ( .a(n_38858), .b(n_38857), .c(n_38856), .o(n_39768) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_17_ ( .ck(newNet_574), .d(n_17770), .o(delay_xor_ln22_unr12_stage5_stallmux_q_17_) );
na02f80 g750777 ( .a(n_29120), .b(n_28805), .o(n_29196) );
in01f80 newInst_2670 ( .a(newNet_745), .o(newNet_2670) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_12_ ( .ck(newNet_3169), .d(n_40441), .o(delay_add_ln22_unr27_stage10_stallmux_q_12_) );
in01f80 newInst_3411 ( .a(newNet_3318), .o(newNet_3411) );
in01f80 FE_OCP_RBC1711_n_21087 ( .a(n_21087), .o(FE_OCP_RBN1711_n_21087) );
na02f80 g749865 ( .a(FE_OCP_RBN3011_n_31117), .b(n_31216), .o(n_31284) );
na02f80 g742430 ( .a(n_37668), .b(n_37696), .o(n_37745) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_4_ ( .ck(newNet_951), .d(n_22770), .o(delay_xor_ln21_unr15_stage6_stallmux_q_4_) );
in01f80 g779521 ( .a(n_1478), .o(n_1537) );
no02f80 g764701 ( .a(n_16415), .b(n_15882), .o(n_16449) );
na02f80 g751404 ( .a(n_29287), .b(n_29286), .o(n_29288) );
na02f80 g778759 ( .a(n_2298), .b(n_1177), .o(n_2385) );
na02f80 g763449 ( .a(n_17113), .b(n_17170), .o(n_17319) );
in01f80 g741186 ( .a(n_38987), .o(n_39037) );
in01f80 newInst_588 ( .a(newNet_587), .o(newNet_588) );
no03m80 g748773 ( .a(n_32411), .b(n_32501), .c(n_32444), .o(n_32533) );
no02f80 g742012 ( .a(n_38112), .b(n_38106), .o(n_38183) );
no02f80 g773089 ( .a(n_7886), .b(n_7950), .o(n_8081) );
na02f80 g781028 ( .a(cos_out_3), .b(FE_OFN2_n_43918), .o(n_301) );
na03f80 FE_RC_1038_0 ( .a(n_23237), .b(FE_RN_299_0), .c(n_23113), .o(n_23253) );
in01f80 g774943 ( .a(n_6301), .o(n_6280) );
no02f80 g742462 ( .a(n_37686), .b(n_37709), .o(n_37704) );
ao12f80 g763764 ( .a(n_17211), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n_17702) );
no02f80 g739105 ( .a(n_40999), .b(n_40998), .o(n_41000) );
in01f80 g771551 ( .a(n_9185), .o(n_9186) );
ao22s80 g771029 ( .a(n_9883), .b(n_9665), .c(n_9831), .d(n_9664), .o(n_10042) );
ao12f80 g761715 ( .a(n_19368), .b(n_19401), .c(n_19367), .o(n_19873) );
no02f80 g749457 ( .a(n_30597), .b(n_30466), .o(n_30639) );
na02f80 g741471 ( .a(n_38762), .b(n_38783), .o(n_38797) );
no02f80 g751176 ( .a(n_29837), .b(n_29940), .o(n_29995) );
in01f80 g739172 ( .a(n_40896), .o(n_40868) );
na02f80 g752141 ( .a(n_28113), .b(n_28160), .o(n_28179) );
ao12f80 g764945 ( .a(n_15643), .b(n_15676), .c(n_15606), .o(n_15677) );
na02f80 g757606 ( .a(FE_OCP_RBN2052_delay_xor_ln22_unr15_stage6_stallmux_q_2_), .b(n_44061), .o(n_22714) );
ao22s80 FE_RC_3246_0 ( .a(n_45070), .b(n_20950), .c(n_45032), .d(n_20949), .o(n_21084) );
no02f80 FE_RC_2207_0 ( .a(FE_RN_793_0), .b(n_27150), .o(FE_RN_794_0) );
in01f80 g774205 ( .a(n_6928), .o(n_6929) );
no02f80 g760515 ( .a(n_19967), .b(n_19945), .o(n_20043) );
in01f80 FE_OCP_RBC2002_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN2002_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
na02f80 g738400 ( .a(n_41677), .b(n_41635), .o(n_41703) );
oa22f80 g744587 ( .a(n_36601), .b(n_36219), .c(n_36577), .d(n_36220), .o(n_36663) );
no02f80 g770539 ( .a(n_10436), .b(n_10372), .o(n_10559) );
in01f80 g753403 ( .a(n_27024), .o(n_27025) );
no02f80 g775652 ( .a(n_5409), .b(n_5313), .o(n_5477) );
in01f80 g740578 ( .a(n_39693), .o(n_39694) );
na02f80 g771614 ( .a(n_9165), .b(FE_OCP_RBN3572_n_44563), .o(n_9243) );
in01f80 g757044 ( .a(n_23900), .o(n_23952) );
in01f80 g776336 ( .a(n_4949), .o(n_4950) );
oa22f80 g746182 ( .a(n_33750), .b(n_33752), .c(FE_OCP_RBN3437_n_33750), .d(n_33769), .o(n_33868) );
na02f80 g769375 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n_12115) );
in01f80 g768930 ( .a(n_12110), .o(n_12111) );
in01f80 g739695 ( .a(n_40565), .o(n_40566) );
in01f80 g737212 ( .a(n_43298), .o(n_42972) );
na02f80 g759507 ( .a(n_20912), .b(n_20911), .o(n_21035) );
oa12f80 g758820 ( .a(n_21366), .b(n_21477), .c(n_21397), .o(n_21558) );
na02f80 g748945 ( .a(n_31196), .b(n_31152), .o(n_31262) );
in01f80 newInst_516 ( .a(newNet_515), .o(newNet_516) );
in01f80 FE_OCP_RBC3367_n_44722 ( .a(FE_OCP_RBN3365_n_44722), .o(FE_OCP_RBN3367_n_44722) );
no02f80 g777761 ( .a(n_3312), .b(n_3333), .o(n_3407) );
na02f80 g774751 ( .a(n_6238), .b(n_6170), .o(n_6271) );
in01f80 g752927 ( .a(n_28212), .o(n_28213) );
in01f80 g747821 ( .a(n_33293), .o(n_33359) );
na02f80 g749912 ( .a(n_30384), .b(n_30423), .o(n_30444) );
in01f80 g745591 ( .a(n_34460), .o(n_34403) );
oa22f80 FE_RC_1521_0 ( .a(n_24350), .b(n_27804), .c(n_27845), .d(n_27774), .o(n_27862) );
na02f80 g738027 ( .a(n_42143), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42153) );
na02f80 g740609 ( .a(n_39634), .b(n_45841), .o(n_39660) );
no02f80 g756062 ( .a(n_24994), .b(n_24276), .o(n_24995) );
ao22s80 g739212 ( .a(n_45144), .b(n_40696), .c(n_45144), .d(n_40339), .o(n_40743) );
oa12f80 g741913 ( .a(n_38232), .b(n_38170), .c(n_38254), .o(n_38335) );
ao12f80 g745508 ( .a(n_34451), .b(n_34453), .c(n_44102), .o(n_34538) );
na02f80 g763513 ( .a(FE_OCP_RBN3082_n_16977), .b(n_16088), .o(n_17169) );
in01f80 g779714 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .o(n_1372) );
oa12f80 g754987 ( .a(n_25344), .b(n_25744), .c(n_25193), .o(n_25884) );
no02f80 g742308 ( .a(FE_OCP_RBN3423_n_37794), .b(n_37823), .o(n_37824) );
no02f80 g743387 ( .a(n_36689), .b(n_36672), .o(n_36718) );
na02f80 g746480 ( .a(n_34642), .b(n_34640), .o(n_34670) );
na02f80 g768256 ( .a(n_12697), .b(n_12657), .o(n_12714) );
na02f80 g747426 ( .a(n_33746), .b(n_33516), .o(n_33578) );
na02f80 g764880 ( .a(n_15395), .b(n_15266), .o(n_15477) );
na02f80 g748129 ( .a(n_31743), .b(n_31808), .o(n_31809) );
no02f80 g751863 ( .a(n_28188), .b(delay_add_ln22_unr17_stage7_stallmux_q_6_), .o(n_28210) );
no02f80 FE_RC_3404_0 ( .a(FE_RN_1472_0), .b(FE_RN_1473_0), .o(FE_RN_1474_0) );
in01f80 g743356 ( .a(n_36763), .o(n_36764) );
na02f80 g764912 ( .a(n_15552), .b(n_14452), .o(n_15551) );
no02f80 FE_RC_2306_0 ( .a(FE_RN_873_0), .b(n_25868), .o(FE_RN_874_0) );
no02f80 g745066 ( .a(n_34873), .b(n_34852), .o(n_34853) );
in01f80 FE_OCP_RBC1213_n_31847 ( .a(n_31847), .o(FE_OCP_RBN1213_n_31847) );
na02f80 g776577 ( .a(n_4360), .b(FE_OCP_RBN2528_n_3421), .o(n_4474) );
in01f80 g756219 ( .a(n_24218), .o(n_24219) );
no02f80 g761339 ( .a(n_20134), .b(n_20178), .o(n_20424) );
na02f80 g749838 ( .a(FE_OCP_RBN3012_n_31117), .b(n_31171), .o(n_31287) );
na02f80 g773938 ( .a(n_6993), .b(n_6992), .o(n_7079) );
in01f80 g742939 ( .a(n_37059), .o(n_37060) );
ao12f80 g754365 ( .a(n_25782), .b(n_25704), .c(n_25561), .o(n_25819) );
ao12f80 g752497 ( .a(n_28340), .b(n_28339), .c(n_28338), .o(n_28834) );
no02f80 g759546 ( .a(FE_OCP_RBN1367_n_20763), .b(n_45050), .o(n_20818) );
in01f80 g751388 ( .a(n_29361), .o(n_29362) );
in01f80 g738556 ( .a(n_41672), .o(n_41620) );
na02f80 g740429 ( .a(n_39777), .b(n_39806), .o(n_39829) );
no02f80 FE_RC_2345_0 ( .a(n_32507), .b(n_32408), .o(FE_RN_899_0) );
na02f80 g755051 ( .a(n_25349), .b(n_24422), .o(n_25381) );
oa22f80 g777828 ( .a(n_3192), .b(n_3004), .c(n_3236), .d(n_3005), .o(n_3697) );
in01f80 g763337 ( .a(n_17380), .o(n_17381) );
oa12f80 g784665 ( .a(n_6121), .b(n_6036), .c(n_5889), .o(n_46995) );
ao12f80 g765391 ( .a(n_14789), .b(n_14942), .c(n_14845), .o(n_15023) );
in01f80 FE_OCP_RBC2490_n_3338 ( .a(FE_OCP_RBN2489_n_3338), .o(FE_OCP_RBN2490_n_3338) );
no02f80 g763404 ( .a(FE_OCPN1756_n_16923), .b(FE_OCP_RBN3689_n_16146), .o(n_17076) );
in01f80 g752737 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_11_), .o(n_28367) );
in01f80 g763929 ( .a(n_17261), .o(n_17154) );
in01f80 FE_OCPC1434_n_30614 ( .a(FE_OCPN1433_n_30614), .o(FE_OCPN1434_n_30614) );
in01f80 newInst_2112 ( .a(newNet_1515), .o(newNet_2112) );
oa22f80 g747969 ( .a(n_31881), .b(n_31608), .c(n_31882), .d(n_31609), .o(n_31958) );
na02f80 g750701 ( .a(n_29392), .b(n_29391), .o(n_29413) );
no02f80 g741496 ( .a(n_38739), .b(n_38738), .o(n_38760) );
no02f80 g773673 ( .a(n_7267), .b(n_7141), .o(n_7306) );
oa22f80 FE_RC_2749_0 ( .a(n_8537), .b(n_8756), .c(n_8538), .d(n_8755), .o(n_8889) );
in01f80 FE_OCP_RBC1134_n_16041 ( .a(FE_OCP_RBN1133_n_16041), .o(FE_OCP_RBN1134_n_16041) );
in01f80 FE_RC_581_0 ( .a(n_23391), .o(FE_RN_178_0) );
in01f80 g772790 ( .a(n_8208), .o(n_8209) );
in01f80 g755930 ( .a(n_24457), .o(n_25390) );
in01f80 g752045 ( .a(n_28161), .o(n_28162) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_6_ ( .ck(newNet_486), .d(n_22758), .o(delay_xor_ln22_unr15_stage6_stallmux_q_6_) );
in01f80 newInst_602 ( .a(newNet_601), .o(newNet_602) );
na02f80 g772967 ( .a(n_7820), .b(n_7819), .o(n_7912) );
in01f80 fopt782976 ( .a(n_26208), .o(n_44443) );
no02f80 g778375 ( .a(n_2731), .b(n_3532), .o(n_2770) );
no02f80 g751482 ( .a(n_28736), .b(n_28735), .o(n_28768) );
ao12f80 g747604 ( .a(n_33571), .b(n_33704), .c(n_33762), .o(n_33763) );
in01f80 g748052 ( .a(n_31748), .o(n_31777) );
in01f80 newInst_3362 ( .a(newNet_3234), .o(newNet_3362) );
oa12f80 g739803 ( .a(n_40292), .b(n_40349), .c(n_40218), .o(n_40423) );
in01f80 g736825 ( .a(n_43344), .o(n_43345) );
in01f80 newInst_1180 ( .a(newNet_1179), .o(newNet_1180) );
in01f80 g757286 ( .a(n_23206), .o(n_23207) );
oa22f80 FE_RC_974_0 ( .a(n_32224), .b(n_31858), .c(n_31859), .d(n_32242), .o(n_32338) );
in01f80 g746617 ( .a(n_34496), .o(n_34550) );
oa12f80 g755263 ( .a(n_24966), .b(n_24971), .c(n_24937), .o(n_25038) );
no02f80 g736708 ( .a(n_43317), .b(n_43120), .o(n_43407) );
oa22f80 g742957 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(n_37082), .d(n_36486), .o(n_37423) );
no02f80 FE_RC_221_0 ( .a(FE_RN_74_0), .b(n_11882), .o(n_11763) );
ao12f80 g742166 ( .a(n_38326), .b(n_44887), .c(n_38325), .o(n_38501) );
in01f80 g778108 ( .a(n_3004), .o(n_3005) );
in01f80 FE_RC_4075_0 ( .a(n_44040), .o(FE_RN_1776_0) );
in01f80 g745884 ( .a(n_34124), .o(n_34113) );
ao12f80 g768557 ( .a(n_12323), .b(n_45659), .c(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .o(n_12541) );
no02f80 g751895 ( .a(n_28919), .b(n_29076), .o(n_29101) );
in01f80 newInst_3658 ( .a(newNet_3657), .o(newNet_3658) );
no02f80 g750707 ( .a(n_29279), .b(FE_OCP_RBN3404_n_28597), .o(n_29275) );
oa12f80 g756729 ( .a(n_23430), .b(n_23429), .c(n_23428), .o(n_24825) );
no02f80 g742985 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n_37002) );
in01f80 g737208 ( .a(n_46936), .o(n_42994) );
no02f80 g757179 ( .a(n_23231), .b(n_23228), .o(n_23305) );
na02f80 g742410 ( .a(n_37697), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37698) );
oa12f80 g750577 ( .a(n_29413), .b(n_29513), .c(n_29465), .o(n_29558) );
na02f80 g771649 ( .a(n_8886), .b(n_7573), .o(n_9010) );
na02f80 g759772 ( .a(n_21253), .b(n_21252), .o(n_21254) );
in01f80 g759064 ( .a(n_21391), .o(n_21279) );
na02f80 g755428 ( .a(n_25347), .b(n_25346), .o(n_25348) );
in01f80 newInst_1246 ( .a(newNet_1245), .o(newNet_1246) );
in01f80 g776312 ( .a(n_4616), .o(n_4617) );
in01f80 g738444 ( .a(n_41881), .o(n_41882) );
oa22f80 FE_RC_1476_0 ( .a(n_24350), .b(n_27755), .c(n_27845), .d(n_27729), .o(n_27780) );
no02f80 g759769 ( .a(n_20636), .b(n_18642), .o(n_20677) );
na02f80 g741166 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39232), .o(n_39304) );
no02f80 g772618 ( .a(n_8368), .b(n_8320), .o(n_8396) );
in01f80 g762751 ( .a(n_17847), .o(n_17848) );
na02f80 g741307 ( .a(FE_OCP_RBN2549_n_44944), .b(n_38495), .o(n_38904) );
na02f80 g743596 ( .a(n_36445), .b(n_36193), .o(n_36446) );
in01f80 g740691 ( .a(n_39481), .o(n_39482) );
na02f80 g766877 ( .a(n_14390), .b(n_14298), .o(n_15247) );
in01f80 g768993 ( .a(n_11877), .o(n_11878) );
no02f80 g738982 ( .a(n_41185), .b(n_40813), .o(n_41193) );
in01f80 fopt783676 ( .a(n_25964), .o(n_45329) );
in01f80 g769560 ( .a(n_11503), .o(n_11504) );
in01f80 g755759 ( .a(n_25286), .o(n_25287) );
oa12f80 g750407 ( .a(n_29630), .b(n_29594), .c(n_29545), .o(n_29631) );
in01f80 g736899 ( .a(n_43581), .o(n_43582) );
in01f80 g752629 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_), .o(n_28466) );
in01f80 FE_OCPC1017_n_23307 ( .a(FE_OCPN1016_n_23307), .o(FE_OCPN1017_n_23307) );
na02f80 g738344 ( .a(n_41793), .b(n_41711), .o(n_41794) );
oa12f80 g769659 ( .a(n_11142), .b(n_11247), .c(FE_OCP_RBN3037_n_47269), .o(n_11274) );
ao12f80 g739249 ( .a(n_40815), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_19_), .o(n_41168) );
in01f80 g741402 ( .a(n_38841), .o(n_38842) );
in01f80 g778662 ( .a(n_2544), .o(n_2545) );
in01f80 newInst_2937 ( .a(newNet_2936), .o(newNet_2937) );
na02f80 g756927 ( .a(n_24352), .b(n_24086), .o(n_24845) );
na02f80 FE_RC_2352_0 ( .a(n_1645), .b(n_1646), .o(FE_RN_905_0) );
na02f80 g751330 ( .a(n_29601), .b(n_29102), .o(n_29597) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_14_ ( .ck(newNet_2677), .d(n_22236), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_) );
no03m80 g742487 ( .a(n_37514), .b(n_37515), .c(n_37118), .o(n_37537) );
no02f80 g746029 ( .a(n_34007), .b(n_34006), .o(n_34008) );
na02f80 g764433 ( .a(FE_OCP_RBN2868_n_16088), .b(n_14588), .o(n_16164) );
oa12f80 g754741 ( .a(n_26231), .b(n_26230), .c(n_26307), .o(n_26383) );
ao12f80 g741977 ( .a(n_37952), .b(n_37951), .c(n_37950), .o(n_38817) );
na02f80 g773430 ( .a(n_7584), .b(n_6631), .o(n_8635) );
no02f80 g741070 ( .a(n_39039), .b(FE_OCP_RBN2546_n_44944), .o(n_39102) );
in01f80 newInst_1728 ( .a(newNet_1390), .o(newNet_1728) );
no02f80 g740389 ( .a(n_39803), .b(n_39520), .o(n_39937) );
na02f80 g745879 ( .a(n_34052), .b(n_34051), .o(n_34067) );
ao22s80 FE_RC_828_0 ( .a(n_24010), .b(n_24399), .c(n_24009), .d(n_24398), .o(n_24501) );
in01f80 newInst_2888 ( .a(newNet_2887), .o(newNet_2888) );
na02f80 g771814 ( .a(n_8962), .b(n_8961), .o(n_8963) );
in01f80 g780180 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_19_), .o(n_1101) );
na02f80 g753578 ( .a(n_26661), .b(n_26317), .o(n_26700) );
ao12f80 g743057 ( .a(n_36922), .b(n_36936), .c(n_36934), .o(n_36937) );
no02f80 g747725 ( .a(n_33671), .b(n_33626), .o(n_33479) );
oa12f80 g738989 ( .a(n_41077), .b(n_41192), .c(n_41107), .o(n_41226) );
in01f80 g778565 ( .a(FE_OFN817_n_2285), .o(n_2876) );
in01f80 newInst_2956 ( .a(newNet_2955), .o(newNet_2956) );
in01f80 g752216 ( .a(n_28987), .o(n_28557) );
in01f80 g757469 ( .a(n_23901), .o(n_23399) );
in01f80 g749568 ( .a(n_30436), .o(n_30437) );
in01f80 FE_OCP_RBC3336_n_44610 ( .a(n_44610), .o(FE_OCP_RBN3336_n_44610) );
oa12f80 g740497 ( .a(n_39767), .b(n_39766), .c(n_39765), .o(n_39786) );
no02f80 g756365 ( .a(n_23827), .b(n_23797), .o(n_23798) );
oa22f80 FE_RC_727_0 ( .a(n_7486), .b(n_8112), .c(n_8111), .d(n_7487), .o(n_8221) );
in01f80 FE_RC_3137_0 ( .a(FE_RN_1392_0), .o(n_16868) );
ao12f80 g774222 ( .a(n_6870), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .o(n_6926) );
in01f80 newInst_3744 ( .a(newNet_1449), .o(newNet_3744) );
in01f80 FE_OCP_RBC3517_n_8498 ( .a(FE_OCP_RBN3516_n_8498), .o(FE_OCP_RBN3517_n_8498) );
in01f80 g746524 ( .a(n_34529), .o(n_34500) );
na02f80 g765224 ( .a(n_15720), .b(n_15719), .o(n_15930) );
na02f80 g775338 ( .a(n_5700), .b(n_4875), .o(n_5735) );
na02f80 g754327 ( .a(n_25843), .b(n_25537), .o(n_25876) );
in01f80 g748924 ( .a(n_32403), .o(n_32404) );
oa12f80 g754204 ( .a(n_26745), .b(n_26744), .c(n_26743), .o(n_26796) );
na02f80 g741737 ( .a(n_38475), .b(n_38134), .o(n_38531) );
no02f80 g757993 ( .a(n_22413), .b(n_22438), .o(n_22442) );
na02f80 g777116 ( .a(n_3604), .b(n_3803), .o(n_3840) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_20_ ( .ck(newNet_1316), .d(n_1244), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_) );
in01f80 newInst_2252 ( .a(newNet_2251), .o(newNet_2252) );
in01f80 g750681 ( .a(n_30416), .o(n_30417) );
oa12f80 g749693 ( .a(n_30024), .b(n_30056), .c(n_30023), .o(n_31473) );
na02f80 g757332 ( .a(n_22971), .b(n_22938), .o(n_23020) );
in01f80 g774433 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_25_), .o(n_6509) );
na02f80 g741748 ( .a(n_38453), .b(n_38158), .o(n_38497) );
oa12f80 g756422 ( .a(n_23427), .b(n_23615), .c(n_23394), .o(n_23640) );
in01f80 g776824 ( .a(n_3822), .o(n_3894) );
in01f80 g758515 ( .a(n_21971), .o(n_21972) );
no02f80 g753185 ( .a(n_27207), .b(FE_OCP_RBN1142_n_25816), .o(n_27392) );
in01f80 newInst_3708 ( .a(newNet_3707), .o(newNet_3708) );
na02f80 g773594 ( .a(n_7350), .b(n_7382), .o(n_7399) );
in01f80 g769871 ( .a(n_11056), .o(n_11083) );
in01f80 g749939 ( .a(n_30145), .o(n_30146) );
na02f80 g744782 ( .a(n_45221), .b(n_35059), .o(n_35123) );
no02f80 g760577 ( .a(n_20354), .b(n_20353), .o(n_20450) );
in01f80 g743477 ( .a(n_36569), .o(n_36552) );
ao22s80 FE_RC_230_0 ( .a(n_13929), .b(n_13022), .c(n_13023), .d(n_13928), .o(n_14069) );
na02f80 FE_RC_3037_0 ( .a(n_11419), .b(n_11415), .o(FE_RN_1330_0) );
in01f80 g762372 ( .a(n_18575), .o(n_18576) );
na02f80 g753485 ( .a(n_26877), .b(n_26823), .o(n_26915) );
ao12f80 g748059 ( .a(n_31754), .b(n_31853), .c(n_31799), .o(n_31935) );
in01f80 g779003 ( .a(n_2186), .o(n_2201) );
na02f80 g761441 ( .a(n_19578), .b(n_19577), .o(n_19579) );
in01f80 g747561 ( .a(n_32517), .o(n_32466) );
na02f80 g769196 ( .a(n_12084), .b(n_12047), .o(n_12702) );
in01f80 g749405 ( .a(n_31979), .o(n_31980) );
in01f80 FE_OFC827_n_1941 ( .a(n_1941), .o(FE_OFN827_n_1941) );
no02f80 g750115 ( .a(FE_OCP_RBN2573_n_29922), .b(n_29398), .o(n_30279) );
ao12f80 g739986 ( .a(n_39907), .b(n_39871), .c(n_39816), .o(n_39987) );
in01f80 g763117 ( .a(n_17414), .o(n_17452) );
na02f80 g753980 ( .a(n_26249), .b(n_26248), .o(n_26278) );
no02f80 g756766 ( .a(n_23458), .b(n_23457), .o(n_23459) );
in01f80 g756657 ( .a(n_23821), .o(n_23783) );
na02f80 g770225 ( .a(n_10667), .b(n_10736), .o(n_10741) );
no02f80 g768541 ( .a(n_12333), .b(n_12311), .o(n_12352) );
oa22f80 g743660 ( .a(n_36325), .b(n_36291), .c(n_36326), .d(n_36292), .o(n_36396) );
in01f80 g765202 ( .a(n_15408), .o(n_15409) );
in01f80 fopt782743 ( .a(n_22677), .o(n_44155) );
oa22f80 g775116 ( .a(n_6024), .b(n_5258), .c(n_6062), .d(n_5259), .o(n_6085) );
in01f80 g765531 ( .a(n_15839), .o(n_15710) );
no04s80 g747182 ( .a(FE_OCPN1015_n_32820), .b(n_32818), .c(FE_OCP_RBN2154_n_32772), .d(n_32634), .o(n_32856) );
in01f80 g766084 ( .a(n_14709), .o(n_14710) );
in01f80 g751081 ( .a(n_28888), .o(n_28889) );
oa22f80 g779659 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .c(FE_OCPN946_n_1780), .d(n_756), .o(n_1626) );
in01f80 newInst_2342 ( .a(newNet_2341), .o(newNet_2342) );
no02f80 g763226 ( .a(n_17277), .b(n_17241), .o(n_17479) );
in01f80 newInst_29 ( .a(newNet_28), .o(newNet_29) );
na02f80 g759763 ( .a(n_21519), .b(n_21402), .o(n_21564) );
oa12f80 g762699 ( .a(n_17946), .b(n_17892), .c(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_18133) );
in01f80 newInst_735 ( .a(newNet_422), .o(newNet_735) );
no02f80 g766660 ( .a(n_13856), .b(n_13351), .o(n_13915) );
in01f80 g760888 ( .a(n_20198), .o(n_21819) );
in01f80 FE_OCPC1414_n_19715 ( .a(FE_OCPN1413_n_19715), .o(FE_OCPN1414_n_19715) );
no02f80 g773621 ( .a(n_7393), .b(n_7392), .o(n_7394) );
in01f80 g738997 ( .a(n_41576), .o(n_41219) );
no02f80 g755729 ( .a(n_25007), .b(n_25092), .o(n_25062) );
no02f80 g755876 ( .a(n_25217), .b(n_25216), .o(n_25799) );
no03m80 FE_RC_3832_0 ( .a(n_23126), .b(FE_RN_1671_0), .c(n_23226), .o(n_23246) );
in01f80 g739482 ( .a(n_40711), .o(n_40712) );
in01f80 g749093 ( .a(n_30885), .o(n_30886) );
in01f80 g780399 ( .a(n_789), .o(n_856) );
na02f80 g740444 ( .a(n_39727), .b(n_39668), .o(n_39729) );
ao12f80 g765217 ( .a(n_15110), .b(n_15136), .c(n_15195), .o(n_15243) );
in01f80 newInst_1650 ( .a(newNet_1649), .o(newNet_1650) );
na02f80 g755886 ( .a(n_25160), .b(n_25304), .o(n_25368) );
in01f80 newInst_3556 ( .a(newNet_3555), .o(newNet_3556) );
in01f80 g763497 ( .a(n_16984), .o(n_16985) );
no02f80 g771367 ( .a(n_9113), .b(n_9112), .o(n_9261) );
na02f80 g753310 ( .a(n_27110), .b(n_26213), .o(n_27297) );
in01f80 g764101 ( .a(n_16745), .o(n_16746) );
in01f80 fopt782845 ( .a(n_44275), .o(n_44267) );
in01f80 g739345 ( .a(n_40704), .o(n_40691) );
na02f80 g738376 ( .a(n_41547), .b(FE_OCP_RBN2312_n_41420), .o(n_41645) );
in01f80 newInst_3168 ( .a(newNet_3167), .o(newNet_3168) );
in01f80 g747520 ( .a(n_32340), .o(n_32309) );
no02f80 g754230 ( .a(n_46962), .b(n_23259), .o(n_25968) );
no02f80 g779200 ( .a(n_1924), .b(n_1923), .o(n_1925) );
in01f80 g744700 ( .a(n_35266), .o(n_35267) );
in01f80 g771686 ( .a(n_9237), .o(n_9286) );
na02f80 g748380 ( .a(FE_OCP_RBN3090_FE_OCPN1052_n_31674), .b(n_30505), .o(n_31793) );
na02f80 g763599 ( .a(n_17430), .b(n_17421), .o(n_17431) );
oa12f80 g745351 ( .a(n_34148), .b(n_34226), .c(n_34114), .o(n_34275) );
no02f80 g763207 ( .a(n_17283), .b(n_16982), .o(n_17285) );
in01f80 g751265 ( .a(n_30095), .o(n_29797) );
in01f80 g759341 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_), .o(n_22898) );
in01f80 g738126 ( .a(n_42072), .o(n_42093) );
in01f80 FE_OCP_RBC2436_n_14072 ( .a(FE_OCP_RBN2435_n_14072), .o(FE_OCP_RBN2436_n_14072) );
in01f80 g784728 ( .a(n_47212), .o(n_47213) );
no02f80 g776805 ( .a(n_4100), .b(n_2532), .o(n_4304) );
no02f80 g743160 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_5_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_5_), .o(n_36922) );
no03m80 g743205 ( .a(n_38076), .b(n_38128), .c(n_38093), .o(n_38174) );
no02f80 g744037 ( .a(n_44221), .b(n_34541), .o(n_35754) );
no02f80 g744804 ( .a(n_35249), .b(FE_OCPN1794_n_30612), .o(n_35250) );
na02f80 g764475 ( .a(n_16119), .b(n_16090), .o(n_16285) );
in01f80 g756672 ( .a(n_24132), .o(n_24192) );
no02f80 g774997 ( .a(n_5973), .b(n_6013), .o(n_6059) );
no02f80 g774808 ( .a(n_6228), .b(n_5640), .o(n_6272) );
in01f80 g771193 ( .a(n_9553), .o(n_9573) );
ao12f80 g749696 ( .a(n_29931), .b(n_29970), .c(n_29930), .o(n_31676) );
na02f80 g746128 ( .a(FE_OCP_RBN3440_n_33803), .b(n_33849), .o(n_33850) );
na02f80 g739156 ( .a(n_40896), .b(n_41007), .o(n_41011) );
in01f80 newInst_1471 ( .a(newNet_1470), .o(newNet_1471) );
in01f80 newInst_1473 ( .a(newNet_303), .o(newNet_1473) );
no02f80 g780377 ( .a(n_1155), .b(n_876), .o(n_877) );
no02f80 g764564 ( .a(n_16007), .b(n_14524), .o(n_16010) );
in01f80 FE_RC_3403_0 ( .a(n_19246), .o(FE_RN_1473_0) );
no02f80 g749359 ( .a(FE_OCP_RBN2806_n_30643), .b(FE_OCP_DRV_N3158_n_27062), .o(n_30701) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_12_ ( .ck(newNet_847), .d(n_1329), .o(delay_xor_ln21_unr3_stage2_stallmux_q_12_) );
oa22f80 FE_RC_3903_0 ( .a(FE_OCP_RBN2423_n_24501), .b(n_44423), .c(n_24555), .d(n_24990), .o(n_25102) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_24_ ( .ck(newNet_1394), .d(n_36663), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_) );
oa22f80 g745570 ( .a(n_34369), .b(n_34039), .c(n_34286), .d(n_46955), .o(n_34743) );
ao12f80 g760215 ( .a(n_20191), .b(n_20171), .c(n_20192), .o(n_20290) );
no02f80 g751039 ( .a(n_30157), .b(n_30085), .o(n_30158) );
in01f80 newInst_3641 ( .a(newNet_3640), .o(newNet_3641) );
in01f80 FE_OCP_RBC2803_n_15706 ( .a(FE_OCP_RBN2801_n_15706), .o(FE_OCP_RBN2803_n_15706) );
in01f80 g770251 ( .a(n_10795), .o(n_10796) );
in01f80 g741996 ( .a(n_38376), .o(n_38377) );
in01f80 g736828 ( .a(n_43551), .o(n_43552) );
ao12f80 g741776 ( .a(n_38452), .b(n_38451), .c(n_38450), .o(n_38512) );
in01f80 newInst_2971 ( .a(newNet_1170), .o(newNet_2971) );
no02f80 g741279 ( .a(n_44921), .b(n_46951), .o(n_39043) );
na02f80 g746734 ( .a(n_33188), .b(n_33107), .o(n_33220) );
na02f80 g766493 ( .a(n_13932), .b(FE_OCP_RBN2249_n_13017), .o(n_14005) );
no02f80 FE_RC_2356_0 ( .a(FE_RN_903_0), .b(FE_RN_908_0), .o(n_45718) );
na02f80 g761726 ( .a(n_19339), .b(n_18774), .o(n_19404) );
ao12f80 g744390 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .b(n_36785), .c(n_36784), .o(n_36793) );
oa22f80 g765410 ( .a(n_15874), .b(n_15631), .c(n_16245), .d(n_14391), .o(n_16355) );
no02f80 g758081 ( .a(n_22005), .b(FE_OCPN1416_FE_OCP_RBN1362_n_20504), .o(n_22027) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_2_ ( .ck(newNet_860), .d(n_40600), .o(delay_xor_ln21_unr28_stage10_stallmux_q_2_) );
oa12f80 g746017 ( .a(n_33778), .b(n_33877), .c(n_33829), .o(n_33925) );
oa12f80 g772688 ( .a(n_7432), .b(n_7986), .c(n_7395), .o(n_8101) );
in01f80 g761984 ( .a(n_18268), .o(n_18284) );
in01f80 newInst_397 ( .a(newNet_192), .o(newNet_397) );
ao12f80 g745782 ( .a(n_34141), .b(n_34140), .c(n_34139), .o(n_35367) );
ao12f80 g736390 ( .a(n_43684), .b(n_43822), .c(n_43429), .o(n_43840) );
in01f80 FE_OCP_RBC2965_n_26231 ( .a(FE_OCP_RBN2963_n_26231), .o(FE_OCP_RBN2965_n_26231) );
in01f80 g740210 ( .a(n_39898), .o(n_39899) );
no02f80 g775928 ( .a(n_5322), .b(n_3817), .o(n_5412) );
in01f80 g777450 ( .a(n_3637), .o(n_3734) );
na02f80 g770282 ( .a(n_10749), .b(n_10811), .o(n_10834) );
in01f80 g762342 ( .a(n_18451), .o(n_18452) );
no02f80 g761322 ( .a(n_19848), .b(n_19845), .o(n_20014) );
na02f80 g772409 ( .a(n_8421), .b(n_8466), .o(n_8520) );
no02f80 g744486 ( .a(n_35416), .b(n_35415), .o(n_35459) );
na02f80 FE_RC_2613_0 ( .a(n_14510), .b(n_14508), .o(FE_RN_1087_0) );
no02f80 g748983 ( .a(n_31126), .b(n_31125), .o(n_31151) );
na02f80 g737613 ( .a(n_42437), .b(n_42463), .o(n_42487) );
in01f80 newInst_1001 ( .a(newNet_675), .o(newNet_1001) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_23_ ( .ck(newNet_329), .d(n_1357), .o(delay_xor_ln22_unr3_stage2_stallmux_q_23_) );
no02f80 g760077 ( .a(n_20778), .b(n_20662), .o(n_20784) );
no02f80 g759008 ( .a(n_21279), .b(n_21323), .o(n_21471) );
no02f80 g753777 ( .a(n_26469), .b(n_26468), .o(n_26559) );
in01f80 g750038 ( .a(n_30347), .o(n_30348) );
in01f80 g776054 ( .a(n_5153), .o(n_5154) );
no02f80 g756922 ( .a(n_23704), .b(n_23908), .o(n_24672) );
na02f80 g763605 ( .a(n_16732), .b(n_16737), .o(n_16792) );
in01f80 g738349 ( .a(n_41646), .o(n_41647) );
no02f80 g771739 ( .a(n_8863), .b(n_8840), .o(n_8841) );
na02f80 g738387 ( .a(n_41621), .b(n_41638), .o(n_41710) );
in01f80 newInst_2777 ( .a(newNet_2776), .o(newNet_2777) );
no02f80 g774549 ( .a(n_6806), .b(FE_OCP_RBN1987_delay_xor_ln23_unr6_stage3_stallmux_q), .o(n_7070) );
in01f80 g768901 ( .a(n_11823), .o(n_11850) );
na02f80 g773742 ( .a(n_7240), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .o(n_7305) );
in01f80 g742609 ( .a(n_37551), .o(n_37567) );
in01f80 g764676 ( .a(n_15856), .o(n_15903) );
na03f80 FE_RC_1493_0 ( .a(n_16899), .b(n_16988), .c(n_16894), .o(n_17245) );
in01f80 g764243 ( .a(n_16443), .o(n_16444) );
oa12f80 g739079 ( .a(n_40971), .b(n_41051), .c(n_40988), .o(n_41075) );
no02f80 g760130 ( .a(n_20429), .b(n_19461), .o(n_20574) );
in01f80 g763060 ( .a(n_17639), .o(n_17640) );
oa22f80 FE_RC_1447_0 ( .a(n_32287), .b(FE_OCP_RBN3121_n_32239), .c(n_28336), .d(n_32239), .o(n_32288) );
na02f80 FE_RC_1336_0 ( .a(FE_RN_396_0), .b(FE_RN_397_0), .o(FE_RN_398_0) );
in01f80 newInst_2386 ( .a(newNet_614), .o(newNet_2386) );
no02f80 g764629 ( .a(n_15901), .b(n_15708), .o(n_15949) );
in01f80 g752327 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .o(n_27803) );
in01f80 g762340 ( .a(n_18453), .o(n_18581) );
in01f80 g741682 ( .a(n_38569), .o(n_38568) );
in01f80 FE_RC_2244_0 ( .a(n_37034), .o(FE_RN_823_0) );
na02f80 g755990 ( .a(n_24231), .b(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24232) );
in01f80 FE_OCPC1419_n_14003 ( .a(n_14003), .o(FE_OCPN1419_n_14003) );
na02f80 g758258 ( .a(n_22608), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22621) );
in01f80 g779025 ( .a(n_2187), .o(n_2188) );
na02f80 g740173 ( .a(FE_OCP_RBN3056_n_39913), .b(n_39627), .o(n_40074) );
na02f80 g744144 ( .a(n_35687), .b(n_35684), .o(n_35735) );
na02f80 g755626 ( .a(n_24471), .b(n_24502), .o(n_24472) );
na02f80 FE_RC_165_0 ( .a(FE_RN_50_0), .b(n_11999), .o(n_12100) );
in01f80 newInst_3150 ( .a(newNet_3149), .o(newNet_3150) );
in01f80 g762367 ( .a(n_18612), .o(n_18613) );
in01f80 g746942 ( .a(n_32920), .o(n_32895) );
no02f80 g779585 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_24_), .o(n_2026) );
in01f80 newInst_386 ( .a(newNet_385), .o(newNet_386) );
in01f80 g738256 ( .a(n_41949), .o(n_41923) );
no02f80 g768398 ( .a(n_12528), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .o(n_12539) );
na02f80 g776854 ( .a(n_4149), .b(n_4020), .o(n_4202) );
na02f80 g758050 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .o(n_23116) );
in01f80 FE_OCPC1737_n_19052 ( .a(n_19052), .o(FE_OCPN1737_n_19052) );
na02f80 g748605 ( .a(n_32611), .b(n_32562), .o(n_32658) );
no02f80 FE_RC_682_0 ( .a(FE_RN_219_0), .b(FE_RN_220_0), .o(FE_RN_221_0) );
in01f80 g772601 ( .a(n_8423), .o(n_8424) );
in01f80 g739641 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_25_), .o(n_40572) );
ao12f80 g774053 ( .a(n_7173), .b(n_7172), .c(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .o(n_7374) );
na02f80 g748719 ( .a(n_31441), .b(n_31377), .o(n_31419) );
in01f80 newInst_884 ( .a(newNet_58), .o(newNet_884) );
in01f80 g748973 ( .a(n_31132), .o(n_31153) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_25_ ( .ck(newNet_3517), .d(n_22818), .o(delay_add_ln22_unr14_stage6_stallmux_q_25_) );
no02f80 g777139 ( .a(n_3659), .b(n_3643), .o(n_3660) );
in01f80 g762612 ( .a(n_18045), .o(n_18046) );
no02f80 g777057 ( .a(n_3720), .b(n_3029), .o(n_3918) );
na02f80 g779773 ( .a(n_1780), .b(n_1392), .o(n_1393) );
na02f80 g778118 ( .a(n_2917), .b(n_2890), .o(n_3024) );
in01f80 g749206 ( .a(n_30914), .o(n_30939) );
na02f80 g758685 ( .a(n_21946), .b(n_20275), .o(n_21961) );
ao12f80 g778363 ( .a(n_2489), .b(n_2488), .c(n_2487), .o(n_2583) );
na02f80 g750978 ( .a(FE_OCP_RBN2631_n_29947), .b(n_30003), .o(n_30005) );
oa22f80 g739893 ( .a(n_40092), .b(n_40328), .c(n_40123), .d(n_40329), .o(n_40411) );
in01f80 FE_RC_3538_0 ( .a(FE_OFN779_n_17093), .o(FE_RN_1531_0) );
in01f80 FE_OCPC1516_n_35367 ( .a(FE_OCPN1515_n_35367), .o(FE_OCPN1516_n_35367) );
in01f80 newInst_22 ( .a(newNet_20), .o(newNet_22) );
in01f80 newInst_2260 ( .a(newNet_2259), .o(newNet_2260) );
na02f80 g774798 ( .a(n_45214), .b(n_6192), .o(n_6253) );
no02f80 g752125 ( .a(n_28709), .b(n_28216), .o(n_28729) );
no02f80 g760928 ( .a(n_19256), .b(n_18506), .o(n_19335) );
na02f80 g738263 ( .a(n_41870), .b(n_41869), .o(n_41871) );
in01f80 g751722 ( .a(n_28349), .o(n_28350) );
in01f80 FE_OCP_RBC2530_n_9044 ( .a(n_9044), .o(FE_OCP_RBN2530_n_9044) );
in01f80 g761280 ( .a(n_18955), .o(n_18956) );
oa22f80 FE_RC_117_0 ( .a(FE_OCP_RBN1341_n_19077), .b(n_19326), .c(n_19325), .d(FE_OCP_RBN1342_n_19077), .o(n_19419) );
in01f80 g757089 ( .a(n_23345), .o(n_23389) );
in01f80 g743181 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42196) );
no02f80 g754216 ( .a(n_25914), .b(n_23259), .o(n_25970) );
na02f80 g771087 ( .a(n_10029), .b(n_10028), .o(n_10070) );
in01f80 g756630 ( .a(n_23627), .o(n_23628) );
in01f80 g766452 ( .a(n_14266), .o(n_14267) );
oa22f80 g766203 ( .a(n_14384), .b(n_13514), .c(n_45521), .d(n_13515), .o(n_14539) );
ao12f80 g761167 ( .a(n_19188), .b(n_19187), .c(n_19186), .o(n_21007) );
in01f80 FE_OCP_RBC2230_n_13141 ( .a(n_13141), .o(FE_OCP_RBN2230_n_13141) );
in01f80 g774214 ( .a(n_7034), .o(n_7035) );
ao12f80 g756890 ( .a(n_23368), .b(n_23367), .c(n_23366), .o(n_24764) );
in01f80 g736784 ( .a(n_43427), .o(n_43428) );
oa12f80 g780146 ( .a(n_935), .b(n_1162), .c(n_1061), .o(n_1175) );
oa22f80 g775855 ( .a(n_4714), .b(n_4850), .c(n_4849), .d(n_4715), .o(n_5003) );
no02f80 g753150 ( .a(n_27378), .b(n_27332), .o(n_27488) );
no02f80 g737892 ( .a(n_42270), .b(n_42569), .o(n_42606) );
in01f80 newInst_46 ( .a(newNet_32), .o(newNet_46) );
in01f80 g750253 ( .a(n_29841), .o(n_29857) );
na02f80 g766253 ( .a(n_14461), .b(n_14497), .o(n_14590) );
in01f80 g776107 ( .a(n_5145), .o(n_5146) );
no02f80 g769351 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n_11709) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_25_ ( .ck(newNet_2547), .d(n_27782), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_25_) );
in01f80 newInst_2853 ( .a(newNet_404), .o(newNet_2853) );
no02f80 g777326 ( .a(n_4182), .b(FE_OFN820_n_4333), .o(n_4504) );
no02f80 g746824 ( .a(n_33063), .b(n_33104), .o(n_33080) );
na02f80 g757974 ( .a(n_22085), .b(n_22084), .o(n_22108) );
in01f80 g778589 ( .a(n_2732), .o(n_2733) );
na02f80 g738978 ( .a(n_41149), .b(n_40827), .o(n_41171) );
oa12f80 g775350 ( .a(n_5879), .b(n_5892), .c(n_5843), .o(n_5934) );
ao22s80 g784421 ( .a(n_36541), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n_46233) );
na02f80 g775577 ( .a(n_5477), .b(n_5472), .o(n_5515) );
na02f80 g738039 ( .a(n_42137), .b(n_42570), .o(n_42138) );
ao12f80 g742663 ( .a(n_37458), .b(n_37457), .c(n_37456), .o(n_37554) );
oa12f80 g781084 ( .a(n_89), .b(n_258), .c(n_120), .o(n_259) );
no02f80 g769007 ( .a(n_11690), .b(n_11737), .o(n_11991) );
in01f80 newInst_2283 ( .a(newNet_2282), .o(newNet_2283) );
in01f80 newInst_174 ( .a(newNet_173), .o(newNet_174) );
in01f80 g745205 ( .a(n_34572), .o(n_34656) );
no02f80 g744685 ( .a(n_35157), .b(n_35147), .o(n_35212) );
in01f80 g771660 ( .a(n_9025), .o(n_9026) );
in01f80 FE_RC_3626_0 ( .a(FE_RN_1588_0), .o(FE_RN_1585_0) );
in01f80 g757257 ( .a(n_23169), .o(n_23213) );
no02f80 g749317 ( .a(n_30650), .b(n_30261), .o(n_30735) );
in01f80 g771484 ( .a(n_9654), .o(n_9780) );
no02f80 g758281 ( .a(n_21951), .b(n_21812), .o(n_21974) );
in01f80 g742085 ( .a(n_38255), .o(n_38256) );
ao12f80 g742652 ( .a(n_37011), .b(n_37371), .c(n_37133), .o(n_37469) );
in01f80 newInst_882 ( .a(newNet_881), .o(newNet_882) );
no02f80 g737933 ( .a(n_42270), .b(n_42542), .o(n_42556) );
ao22s80 g747345 ( .a(n_32622), .b(n_44962), .c(FE_OCP_RBN2103_n_44962), .d(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .o(n_32680) );
in01f80 newInst_3119 ( .a(newNet_3118), .o(newNet_3119) );
no02f80 g765851 ( .a(n_14857), .b(n_14860), .o(n_14923) );
na02f80 g765155 ( .a(n_15416), .b(n_15415), .o(n_15417) );
na02f80 g779075 ( .a(n_2009), .b(n_1844), .o(n_2000) );
na02f80 g747541 ( .a(n_33397), .b(n_33396), .o(n_33398) );
ao12f80 g739255 ( .a(n_40909), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n_41230) );
in01f80 g744361 ( .a(n_46221), .o(n_36820) );
in01f80 newInst_407 ( .a(newNet_41), .o(newNet_407) );
na02f80 g762029 ( .a(n_18279), .b(n_18313), .o(n_18335) );
oa22f80 FE_RC_3721_0 ( .a(n_38678), .b(n_38653), .c(n_38666), .d(n_38679), .o(n_38739) );
in01f80 g752684 ( .a(n_27442), .o(n_27473) );
oa12f80 g774521 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n_6895) );
in01f80 newInst_2899 ( .a(newNet_2898), .o(newNet_2899) );
no02f80 g759751 ( .a(n_20713), .b(n_20631), .o(n_20714) );
no02f80 g745776 ( .a(n_34283), .b(n_34302), .o(n_34394) );
in01f80 g756773 ( .a(n_23426), .o(n_23441) );
no02f80 g755481 ( .a(n_24746), .b(n_24546), .o(n_24801) );
na02f80 g750459 ( .a(n_29530), .b(FE_OCPN1464_n_29630), .o(n_29550) );
in01f80 g780580 ( .a(n_814), .o(n_790) );
no02f80 g767937 ( .a(n_12694), .b(n_12693), .o(n_12722) );
no02f80 g781256 ( .a(n_66), .b(n_264), .o(n_98) );
oa12f80 g764858 ( .a(n_16354), .b(n_16353), .c(n_16352), .o(n_16412) );
in01f80 fopt782852 ( .a(n_21973), .o(n_44275) );
no02f80 g767700 ( .a(n_12800), .b(n_12677), .o(n_12801) );
na02f80 g770077 ( .a(n_10673), .b(n_10733), .o(n_10734) );
in01f80 g749395 ( .a(n_30697), .o(n_30729) );
no02f80 g777141 ( .a(n_3711), .b(FE_OCP_RBN2623_n_3631), .o(n_3750) );
no02f80 g760629 ( .a(n_20301), .b(n_19851), .o(n_20354) );
in01f80 g772293 ( .a(FE_OCP_RBN2475_n_8664), .o(n_8731) );
no02f80 g749643 ( .a(n_31396), .b(n_31143), .o(n_31433) );
na02f80 g765290 ( .a(n_16018), .b(n_15823), .o(n_15720) );
in01f80 g778623 ( .a(n_2768), .o(n_2769) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_22_ ( .ck(newNet_2471), .d(FE_OCP_RBN3137_n_32380), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_22_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_13_ ( .ck(newNet_2586), .d(n_27365), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_13_) );
in01f80 FE_OCP_RBC2707_n_15135 ( .a(FE_OCP_RBN3621_n_15135), .o(FE_OCP_RBN2707_n_15135) );
na02f80 g754512 ( .a(n_25515), .b(n_25514), .o(n_25516) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_22_ ( .ck(newNet_2280), .d(n_40506), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_) );
in01f80 newInst_536 ( .a(newNet_535), .o(newNet_536) );
ao12f80 g773727 ( .a(n_6718), .b(n_7280), .c(n_6767), .o(n_7314) );
in01f80 g763006 ( .a(n_17684), .o(n_17518) );
na02f80 g764485 ( .a(n_16008), .b(n_45332), .o(n_16171) );
no02f80 g752632 ( .a(n_28205), .b(n_27991), .o(n_28206) );
in01f80 g740112 ( .a(n_40249), .o(n_40250) );
in01f80 g755855 ( .a(n_24363), .o(n_24364) );
no02f80 g777851 ( .a(n_3176), .b(n_3027), .o(n_3177) );
na02f80 g776205 ( .a(n_4845), .b(n_4488), .o(n_4946) );
in01f80 newInst_1388 ( .a(newNet_1387), .o(newNet_1388) );
in01f80 g781191 ( .a(n_186), .o(n_179) );
oa12f80 g780731 ( .a(n_453), .b(n_608), .c(n_466), .o(n_609) );
ao22s80 FE_RC_1245_0 ( .a(FE_OCP_RBN2325_n_13616), .b(n_13713), .c(n_13746), .d(n_13616), .o(n_13849) );
no02f80 g775838 ( .a(n_47002), .b(n_5447), .o(n_5501) );
in01f80 g775065 ( .a(n_46995), .o(n_6175) );
in01f80 newInst_3188 ( .a(newNet_2416), .o(newNet_3188) );
no02f80 g752804 ( .a(n_28050), .b(n_28025), .o(n_28445) );
no02f80 g746935 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n_33252) );
in01f80 g738750 ( .a(n_41397), .o(n_41398) );
in01f80 newInst_2705 ( .a(newNet_487), .o(newNet_2705) );
ao22s80 FE_RC_1256_0 ( .a(n_4754), .b(n_4690), .c(n_4753), .d(n_4624), .o(n_4925) );
in01f80 newInst_320 ( .a(newNet_319), .o(newNet_320) );
oa12f80 g760790 ( .a(n_18633), .b(n_19479), .c(n_19478), .o(n_19519) );
oa22f80 FE_RC_4126_0 ( .a(n_35201), .b(n_35475), .c(n_35228), .d(n_35443), .o(n_35505) );
na02f80 g741150 ( .a(n_39183), .b(FE_OCP_RBN2485_n_38601), .o(n_39184) );
in01f80 g750063 ( .a(n_30172), .o(n_30138) );
in01f80 newInst_278 ( .a(newNet_277), .o(newNet_278) );
oa12f80 g761759 ( .a(n_18246), .b(n_18348), .c(n_18223), .o(n_18439) );
no02f80 g750740 ( .a(n_29316), .b(n_29167), .o(n_29319) );
in01f80 g754679 ( .a(FE_OCPN1410_n_27014), .o(n_30466) );
in01f80 g741468 ( .a(n_38802), .o(n_38803) );
na02f80 g742634 ( .a(n_37403), .b(n_37402), .o(n_37404) );
na02f80 g755545 ( .a(n_24476), .b(n_24512), .o(n_24623) );
na02f80 g773521 ( .a(n_7461), .b(n_7492), .o(n_7494) );
oa12f80 g737221 ( .a(n_42801), .b(n_42902), .c(n_42755), .o(n_42948) );
in01f80 FE_OCP_RBC2634_n_30213 ( .a(n_30213), .o(FE_OCP_RBN2634_n_30213) );
na03f80 g742884 ( .a(n_37542), .b(n_45897), .c(n_37308), .o(n_38371) );
oa22f80 g754608 ( .a(FE_OCP_RBN2960_n_26231), .b(n_26162), .c(n_26856), .d(n_26192), .o(n_26931) );
in01f80 g751525 ( .a(n_28845), .o(n_28846) );
in01f80 FE_OCP_RBC2113_n_45224 ( .a(FE_OCP_RBN3268_n_45224), .o(FE_OCP_RBN2113_n_45224) );
in01f80 g766295 ( .a(n_14779), .o(n_15779) );
in01f80 g760076 ( .a(n_20784), .o(n_20785) );
oa12f80 g742678 ( .a(n_37075), .b(n_37379), .c(n_36960), .o(n_37424) );
ao22s80 g737552 ( .a(n_42252), .b(n_42218), .c(n_42251), .d(n_42208), .o(n_43014) );
oa12f80 g760667 ( .a(n_19570), .b(n_19673), .c(n_19556), .o(n_19728) );
in01f80 g743648 ( .a(n_36382), .o(n_36383) );
na02f80 g755082 ( .a(n_25476), .b(n_25501), .o(n_25583) );
in01f80 g740240 ( .a(n_40316), .o(n_40317) );
in01f80 g745028 ( .a(n_34876), .o(n_34877) );
in01f80 newInst_3353 ( .a(newNet_3352), .o(newNet_3353) );
oa22f80 FE_RC_3291_0 ( .a(n_32128), .b(n_32383), .c(n_32129), .d(n_32382), .o(n_32546) );
oa12f80 g765232 ( .a(n_15664), .b(n_15834), .c(n_15833), .o(n_15835) );
na02f80 g749953 ( .a(n_30344), .b(n_30372), .o(n_30403) );
ao12f80 g774383 ( .a(n_6755), .b(n_6624), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .o(n_6922) );
na02f80 g773103 ( .a(n_7699), .b(n_7751), .o(n_7870) );
na02f80 FE_RC_2603_0 ( .a(FE_RN_1079_0), .b(FE_RN_1080_0), .o(FE_RN_1081_0) );
na02f80 g770401 ( .a(n_10444), .b(n_10408), .o(n_10537) );
no02f80 g769204 ( .a(n_12003), .b(n_11936), .o(n_12048) );
no02f80 g749244 ( .a(n_32094), .b(n_31456), .o(n_32114) );
no02f80 g737526 ( .a(n_42379), .b(n_42587), .o(n_42634) );
in01f80 g769084 ( .a(n_11700), .o(n_11701) );
no02f80 g772326 ( .a(n_8511), .b(n_8574), .o(n_8587) );
in01f80 g764312 ( .a(n_16429), .o(n_16430) );
in01f80 g760550 ( .a(n_19963), .o(n_19964) );
in01f80 g748345 ( .a(n_31829), .o(n_31830) );
na02f80 g745374 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35388), .o(n_35799) );
no02f80 g780412 ( .a(n_788), .b(n_936), .o(n_832) );
oa12f80 g762908 ( .a(n_17991), .b(n_17990), .c(n_17989), .o(n_18689) );
na02f80 g745361 ( .a(n_34463), .b(n_34351), .o(n_34464) );
no02f80 g766042 ( .a(n_14648), .b(n_14663), .o(n_14770) );
in01f80 FE_OCP_RBC2471_n_34285 ( .a(n_34285), .o(FE_OCP_RBN2471_n_34285) );
ao12f80 g743710 ( .a(n_35570), .b(n_36247), .c(n_35615), .o(n_36325) );
no02f80 FE_RC_4059_0 ( .a(n_35616), .b(n_35617), .o(FE_RN_1766_0) );
na02f80 g738498 ( .a(FE_OCP_RBN2316_n_41420), .b(n_41332), .o(n_41690) );
in01f80 FE_OCP_RBC2274_n_2457 ( .a(n_2457), .o(FE_OCP_RBN2274_n_2457) );
no02f80 g738335 ( .a(n_41816), .b(n_41794), .o(n_41860) );
no02f80 g743047 ( .a(n_37043), .b(n_37108), .o(n_37330) );
ao12f80 g748838 ( .a(n_32444), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_11_), .o(n_32840) );
in01f80 g740801 ( .a(n_39489), .o(n_39490) );
oa12f80 g755375 ( .a(n_24711), .b(n_24834), .c(n_24775), .o(n_24897) );
no02f80 g751416 ( .a(n_29176), .b(n_29223), .o(n_29224) );
oa12f80 g767447 ( .a(n_12697), .b(n_13097), .c(n_12656), .o(n_13235) );
oa12f80 g757761 ( .a(n_44288), .b(n_22481), .c(n_22482), .o(n_22518) );
na02f80 g753099 ( .a(n_27144), .b(FE_OCP_RBN2782_n_25997), .o(n_27186) );
no02f80 g750183 ( .a(n_29790), .b(n_29789), .o(n_29791) );
in01f80 FE_OCP_RBC3583_n_9245 ( .a(n_9245), .o(FE_OCP_RBN3583_n_9245) );
in01f80 g744027 ( .a(n_35707), .o(n_35624) );
in01f80 g742033 ( .a(n_38349), .o(n_38350) );
in01f80 g740712 ( .a(n_39581), .o(n_39582) );
no02f80 g771077 ( .a(n_10029), .b(n_10028), .o(n_10067) );
in01f80 g779461 ( .a(n_2019), .o(n_2020) );
ao12f80 g747708 ( .a(n_33951), .b(n_33372), .c(n_33670), .o(n_34168) );
in01f80 newInst_3688 ( .a(newNet_3687), .o(newNet_3688) );
in01f80 g771788 ( .a(n_8848), .o(n_8891) );
in01f80 fopt783499 ( .a(FE_OFN751_n_45003), .o(n_45065) );
in01f80 g747625 ( .a(n_33997), .o(n_33480) );
ao12f80 g778010 ( .a(n_2992), .b(n_2991), .c(n_2990), .o(n_4575) );
no02f80 g777875 ( .a(n_3214), .b(n_2913), .o(n_3237) );
no02f80 g743866 ( .a(n_35815), .b(n_36011), .o(n_36045) );
oa12f80 g749745 ( .a(n_31393), .b(FE_OCP_RBN3010_n_31117), .c(n_31281), .o(n_31633) );
in01f80 g747530 ( .a(n_32519), .o(n_32469) );
in01f80 g751252 ( .a(n_29944), .o(n_29932) );
na02f80 g744542 ( .a(n_35387), .b(FE_OCP_RBN3649_n_35169), .o(n_35399) );
in01f80 newInst_836 ( .a(newNet_835), .o(newNet_836) );
no02f80 g760556 ( .a(n_20450), .b(n_19935), .o(n_20423) );
na02f80 FE_RC_903_0 ( .a(FE_RN_266_0), .b(n_30564), .o(n_46959) );
no02f80 g769068 ( .a(n_11502), .b(n_11497), .o(n_11530) );
na02f80 g745407 ( .a(n_36049), .b(n_36111), .o(n_36112) );
in01f80 g743910 ( .a(n_36978), .o(n_36979) );
oa22f80 g759824 ( .a(n_21714), .b(n_21105), .c(n_21691), .d(n_21134), .o(n_21878) );
na02f80 g765286 ( .a(n_15875), .b(n_16255), .o(n_15926) );
oa12f80 g764724 ( .a(n_16028), .b(n_16029), .c(n_16027), .o(n_16105) );
na02f80 g778576 ( .a(n_2303), .b(n_2302), .o(n_2304) );
in01f80 g758091 ( .a(n_22079), .o(n_22164) );
in01f80 fopt784008 ( .a(n_45740), .o(n_45739) );
oa12f80 g768703 ( .a(n_12019), .b(n_12173), .c(n_12091), .o(n_12260) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_16_ ( .ck(newNet_1533), .d(n_32173), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_) );
in01f80 FE_OCP_RBC3558_n_8687 ( .a(n_8687), .o(FE_OCP_RBN3558_n_8687) );
in01f80 newInst_1621 ( .a(newNet_1620), .o(newNet_1621) );
in01f80 newInst_694 ( .a(newNet_693), .o(newNet_694) );
in01f80 FE_OCPC3795_FE_RN_1789_0 ( .a(FE_OCPN3794_FE_RN_1789_0), .o(FE_OCPN3795_FE_RN_1789_0) );
no02f80 g762920 ( .a(n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .o(n_17655) );
in01f80 FE_RC_2228_0 ( .a(n_37175), .o(FE_RN_810_0) );
in01f80 g759078 ( .a(n_21227), .o(n_21228) );
oa22f80 g743252 ( .a(n_36789), .b(n_36787), .c(n_36798), .d(n_36788), .o(n_36866) );
in01f80 newInst_420 ( .a(newNet_126), .o(newNet_420) );
no02f80 g743307 ( .a(n_36676), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36711) );
na02f80 g775726 ( .a(n_5410), .b(n_5150), .o(n_5510) );
no02f80 g740813 ( .a(n_39439), .b(n_39464), .o(n_39900) );
in01f80 g768595 ( .a(n_12275), .o(n_12276) );
in01f80 g763686 ( .a(n_16827), .o(n_16855) );
in01f80 FE_OCP_DRV_C1546_n_18860 ( .a(FE_OCP_DRV_N1545_n_18860), .o(FE_OCP_DRV_N1546_n_18860) );
na02f80 g745623 ( .a(n_34369), .b(n_33581), .o(n_34506) );
in01f80 FE_RC_1915_0 ( .a(FE_RN_603_0), .o(n_19323) );
na02f80 g746310 ( .a(n_33491), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33527) );
no02f80 g746332 ( .a(n_33504), .b(n_33494), .o(n_33594) );
in01f80 g782640 ( .a(n_44034), .o(n_44035) );
no02f80 g748132 ( .a(n_32768), .b(n_32603), .o(n_32783) );
in01f80 g760163 ( .a(n_20461), .o(n_20462) );
na02f80 g760084 ( .a(n_21023), .b(n_21022), .o(n_21024) );
in01f80 FE_RC_3628_0 ( .a(FE_RN_1590_0), .o(n_21092) );
no02f80 g758246 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .o(n_22843) );
oa12f80 g750351 ( .a(n_29668), .b(n_29667), .c(n_29666), .o(n_31264) );
in01f80 FE_OCPC849_n_2306 ( .a(n_2306), .o(FE_OCPN849_n_2306) );
na02f80 g743950 ( .a(n_35650), .b(n_35596), .o(n_35651) );
in01f80 newInst_76 ( .a(newNet_1), .o(newNet_76) );
oa12f80 g777960 ( .a(n_2906), .b(n_3030), .c(n_2830), .o(n_3114) );
na02f80 g756245 ( .a(n_24098), .b(FE_OCPN1780_n_24097), .o(n_24341) );
na02f80 g744863 ( .a(n_34985), .b(n_34961), .o(n_35057) );
oa22f80 FE_RC_928_0 ( .a(n_25850), .b(n_25478), .c(n_25477), .d(n_25849), .o(n_25938) );
no02f80 g776728 ( .a(n_4277), .b(n_4400), .o(n_4278) );
no02f80 g740859 ( .a(n_39380), .b(n_38973), .o(n_39401) );
ao12f80 g751923 ( .a(n_28955), .b(n_28919), .c(n_28942), .o(n_29459) );
na02f80 g774919 ( .a(n_6237), .b(n_6140), .o(n_6303) );
no02f80 g778226 ( .a(n_2679), .b(FE_OCP_RBN2290_n_2438), .o(n_2680) );
in01f80 FE_OCP_RBC2445_n_29684 ( .a(n_29684), .o(FE_OCP_RBN2445_n_29684) );
na02f80 g757824 ( .a(n_22423), .b(n_22388), .o(n_22511) );
in01f80 g748212 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_), .o(n_32793) );
no02f80 g753300 ( .a(n_27120), .b(n_26116), .o(n_27308) );
in01f80 FE_OCPC1461_n_23759 ( .a(n_23759), .o(FE_OCPN1461_n_23759) );
in01f80 FE_OCP_RBC3443_n_37945 ( .a(n_37945), .o(FE_OCP_RBN3443_n_37945) );
in01f80 g740351 ( .a(n_40386), .o(n_40387) );
oa12f80 g765377 ( .a(n_15875), .b(n_15874), .c(n_15958), .o(n_16300) );
ao12f80 g779652 ( .a(n_1643), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .o(n_1771) );
na02f80 g749586 ( .a(n_30407), .b(n_30406), .o(n_30408) );
na02f80 g765535 ( .a(n_15014), .b(n_14986), .o(n_15076) );
in01f80 FE_OCP_RBC2519_n_8762 ( .a(FE_OCP_RBN2518_n_8762), .o(FE_OCP_RBN2519_n_8762) );
na02f80 g743877 ( .a(n_35793), .b(n_35792), .o(n_35794) );
no02f80 g755292 ( .a(n_25066), .b(n_24969), .o(n_25184) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_5_ ( .ck(newNet_488), .d(n_22712), .o(delay_xor_ln22_unr15_stage6_stallmux_q_5_) );
na02f80 g770478 ( .a(n_10501), .b(n_10475), .o(n_10607) );
in01f80 newInst_3695 ( .a(newNet_3449), .o(newNet_3695) );
na02f80 g778740 ( .a(FE_OCPN871_n_2737), .b(n_2738), .o(n_2758) );
in01f80 g771733 ( .a(n_8915), .o(n_10484) );
na02f80 g765883 ( .a(n_14799), .b(n_14817), .o(n_14901) );
no02f80 g736628 ( .a(n_43479), .b(n_43266), .o(n_43527) );
oa12f80 g736658 ( .a(n_317), .b(n_43073), .c(FE_OFN5_n_43918), .o(n_43154) );
in01f80 g772424 ( .a(n_8571), .o(n_8572) );
oa12f80 FE_RC_2368_0 ( .a(FE_RN_917_0), .b(n_45718), .c(FE_RN_918_0), .o(FE_RN_919_0) );
na02f80 g745254 ( .a(n_36222), .b(n_35560), .o(n_35681) );
na02f80 g750324 ( .a(n_29648), .b(n_29604), .o(n_29689) );
ao12f80 g771311 ( .a(n_9346), .b(n_9567), .c(n_9376), .o(n_9639) );
in01f80 g742543 ( .a(n_37595), .o(n_37620) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_5_ ( .ck(newNet_2709), .d(n_15603), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_) );
in01f80 FE_RC_3088_0 ( .a(n_31178), .o(FE_RN_1363_0) );
oa12f80 g780256 ( .a(n_1024), .b(n_1023), .c(FE_OFN50_n_1045), .o(n_1114) );
in01f80 g772377 ( .a(n_46990), .o(n_10374) );
oa22f80 g742823 ( .a(n_38173), .b(n_45891), .c(n_45899), .d(n_45895), .o(n_38525) );
na02f80 g739934 ( .a(n_40257), .b(n_40156), .o(n_40374) );
no02f80 g760734 ( .a(n_19629), .b(FE_OCP_RBN1348_n_19270), .o(n_19694) );
na02f80 g761157 ( .a(FE_OCP_RBN1351_n_19148), .b(FE_OCP_RBN1178_n_18981), .o(n_19262) );
na02f80 g754516 ( .a(n_25429), .b(n_25207), .o(n_25513) );
in01f80 g740982 ( .a(n_39161), .o(n_39162) );
no02f80 g775297 ( .a(n_5894), .b(n_4864), .o(n_5950) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_8_ ( .ck(newNet_204), .d(n_46168), .o(delay_xor_ln22_unr6_stage3_stallmux_q_8_) );
in01f80 newInst_1795 ( .a(newNet_1270), .o(newNet_1795) );
na02f80 g758303 ( .a(FE_OCP_RBN3223_n_22068), .b(n_22251), .o(n_22294) );
no02f80 g779740 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .o(n_1783) );
in01f80 g767914 ( .a(n_12873), .o(n_12999) );
no02f80 g753975 ( .a(n_26267), .b(n_26214), .o(n_26215) );
na02f80 g769851 ( .a(n_11161), .b(n_11133), .o(n_11278) );
in01f80 g754276 ( .a(n_27217), .o(n_25980) );
in01f80 g775788 ( .a(n_5084), .o(n_5128) );
na02f80 g769275 ( .a(n_11439), .b(FE_OCP_RBN3693_n_10852), .o(n_11459) );
ao12f80 g784686 ( .a(n_3496), .b(n_3475), .c(n_3248), .o(n_47016) );
no02f80 g741831 ( .a(n_38288), .b(n_38116), .o(n_38342) );
na02f80 g770582 ( .a(FE_OCP_RBN2794_n_10106), .b(FE_OCP_RBN2499_n_8835), .o(n_10324) );
na02f80 g779247 ( .a(n_1827), .b(n_1033), .o(n_1900) );
in01f80 fopt783209 ( .a(FE_OCP_RBN3308_n_44722), .o(n_44761) );
na02f80 g767671 ( .a(n_12967), .b(n_13000), .o(n_13001) );
no02f80 g742842 ( .a(n_37214), .b(n_37080), .o(n_37230) );
na02f80 g784592 ( .a(n_12823), .b(n_12892), .o(n_46415) );
no02f80 g737375 ( .a(n_42790), .b(n_42506), .o(n_42834) );
in01f80 g737323 ( .a(n_42844), .o(n_42845) );
no02f80 g778125 ( .a(n_2889), .b(n_2674), .o(n_2966) );
in01f80 FE_OFC765_n_15670 ( .a(FE_OFN762_n_15670), .o(FE_OFN765_n_15670) );
no02f80 FE_RC_2353_0 ( .a(FE_RN_905_0), .b(n_1958), .o(FE_RN_906_0) );
in01f80 newInst_3323 ( .a(newNet_3322), .o(newNet_3323) );
in01f80 g760729 ( .a(n_19695), .o(n_19696) );
no02f80 g760504 ( .a(n_19944), .b(n_19685), .o(n_20002) );
no02f80 g752122 ( .a(n_28011), .b(n_28012), .o(n_28013) );
ao12f80 g779067 ( .a(n_2010), .b(n_2009), .c(n_2008), .o(n_2288) );
in01f80 g739144 ( .a(n_40962), .o(n_40976) );
no02f80 g754463 ( .a(n_25601), .b(n_25295), .o(n_25602) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_11_ ( .ck(newNet_1877), .d(n_16593), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_) );
no02f80 g738061 ( .a(n_42090), .b(n_41902), .o(n_42119) );
in01f80 g739315 ( .a(n_40888), .o(n_40845) );
no02f80 g766399 ( .a(n_14231), .b(n_14183), .o(n_14359) );
oa22f80 FE_RC_3320_0 ( .a(n_27893), .b(n_44025), .c(n_27816), .d(n_27859), .o(n_28035) );
no02f80 g757453 ( .a(n_22803), .b(n_44061), .o(n_22870) );
in01f80 FE_OCP_RBC2333_n_38446 ( .a(n_38446), .o(FE_OCP_RBN2333_n_38446) );
na02f80 g778196 ( .a(n_3208), .b(n_3207), .o(n_3209) );
in01f80 newInst_3605 ( .a(newNet_3604), .o(newNet_3605) );
no02f80 g753204 ( .a(n_27204), .b(n_27117), .o(n_27345) );
in01f80 g749649 ( .a(n_30324), .o(n_30350) );
na02f80 g752948 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_), .o(n_27926) );
na02f80 g771144 ( .a(n_9885), .b(n_9921), .o(n_9886) );
in01f80 FE_OCP_RBC2449_n_14114 ( .a(FE_OCP_RBN2448_n_14114), .o(FE_OCP_RBN2449_n_14114) );
in01f80 g749048 ( .a(n_31073), .o(n_31127) );
in01f80 FE_OCP_RBC3609_n_14905 ( .a(n_14905), .o(FE_OCP_RBN3609_n_14905) );
in01f80 g746287 ( .a(n_33706), .o(n_33844) );
na02f80 g781048 ( .a(sin_out_9), .b(FE_OFN3_n_43918), .o(n_320) );
na02f80 g781139 ( .a(n_211), .b(n_210), .o(n_212) );
in01f80 g770157 ( .a(n_10927), .o(n_10982) );
na02f80 g778356 ( .a(n_2507), .b(n_2469), .o(n_2623) );
no02f80 g775220 ( .a(n_5959), .b(n_5784), .o(n_6015) );
in01f80 g774922 ( .a(n_6281), .o(n_6282) );
in01f80 FE_OCP_RBC3128_n_32266 ( .a(n_32266), .o(FE_OCP_RBN3128_n_32266) );
in01f80 newInst_3463 ( .a(newNet_3462), .o(newNet_3463) );
in01f80 FE_OCP_RBC3137_n_32380 ( .a(n_32380), .o(FE_OCP_RBN3137_n_32380) );
no02f80 g752741 ( .a(n_27909), .b(n_27907), .o(n_27908) );
ao22s80 FE_RC_1549_0 ( .a(n_23012), .b(n_23101), .c(n_23011), .d(n_23126), .o(n_23225) );
in01f80 newInst_2755 ( .a(newNet_467), .o(newNet_2755) );
no02f80 FE_RC_1829_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .b(FE_OCP_RBN3284_n_44365), .o(FE_RN_549_0) );
na02f80 FE_RC_1991_0 ( .a(n_18140), .b(n_19580), .o(FE_RN_650_0) );
in01f80 fopt783369 ( .a(n_40579), .o(n_44958) );
no02f80 g759978 ( .a(n_20215), .b(n_20163), .o(n_20229) );
in01f80 newInst_461 ( .a(newNet_460), .o(newNet_461) );
in01f80 newInst_2064 ( .a(newNet_98), .o(newNet_2064) );
in01f80 FE_RC_766_0 ( .a(n_33787), .o(FE_RN_238_0) );
na02f80 g742408 ( .a(n_37718), .b(n_37760), .o(n_37761) );
no02f80 g775081 ( .a(n_5947), .b(n_5963), .o(n_6014) );
in01f80 FE_OCP_RBC2939_n_26276 ( .a(n_26276), .o(FE_OCP_RBN2939_n_26276) );
oa12f80 g761679 ( .a(n_18561), .b(n_18795), .c(n_18560), .o(n_18861) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_20_ ( .ck(newNet_1996), .d(n_11490), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_) );
no02f80 g746712 ( .a(n_34233), .b(n_33991), .o(n_34276) );
na02f80 g776906 ( .a(n_3811), .b(n_3711), .o(n_3864) );
oa12f80 g751322 ( .a(n_29538), .b(n_29537), .c(n_29536), .o(n_29600) );
in01f80 newInst_127 ( .a(newNet_114), .o(newNet_127) );
ao12f80 g752840 ( .a(n_28018), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .o(n_28314) );
no02f80 g757813 ( .a(n_23009), .b(n_22693), .o(n_23092) );
in01f80 g762370 ( .a(n_18841), .o(n_18692) );
in01f80 g759410 ( .a(n_21062), .o(n_21063) );
no02f80 g756478 ( .a(n_23629), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n_23660) );
in01f80 newInst_3330 ( .a(newNet_3329), .o(newNet_3330) );
na02f80 g748910 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .o(n_32495) );
no02f80 g737670 ( .a(FE_OCPN887_n_42367), .b(n_42441), .o(n_42742) );
in01f80 newInst_1300 ( .a(newNet_1005), .o(newNet_1300) );
na02f80 g774786 ( .a(n_45474), .b(n_5693), .o(n_6340) );
in01f80 fopt783253 ( .a(n_44819), .o(n_44818) );
no02f80 g770761 ( .a(n_10252), .b(n_10342), .o(n_10471) );
na02f80 g755436 ( .a(n_24803), .b(n_24754), .o(n_24804) );
oa12f80 g738305 ( .a(n_41744), .b(n_41648), .c(n_41769), .o(n_41839) );
oa12f80 g770190 ( .a(n_9953), .b(n_10869), .c(n_10039), .o(n_10951) );
na02f80 g766913 ( .a(n_13583), .b(n_13570), .o(n_13628) );
in01f80 g774005 ( .a(n_6930), .o(n_6931) );
na02f80 g758113 ( .a(n_44268), .b(FE_OCP_RBN1724_n_21004), .o(n_22227) );
in01f80 FE_OCP_RBC2142_FE_OCPN861_n_45450 ( .a(FE_OCPN861_n_45450), .o(FE_OCP_RBN2142_FE_OCPN861_n_45450) );
na02f80 g739300 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_24_), .o(n_40831) );
na02f80 g770985 ( .a(n_9579), .b(n_9465), .o(n_9580) );
in01f80 g761868 ( .a(n_18784), .o(n_18785) );
in01f80 g749871 ( .a(n_31407), .o(n_31387) );
na02f80 g753514 ( .a(n_26804), .b(n_23564), .o(n_26872) );
no02f80 g779590 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .o(n_1972) );
ao12f80 g754527 ( .a(n_26541), .b(n_26708), .c(n_26643), .o(n_26644) );
na02f80 g736985 ( .a(n_43242), .b(n_43002), .o(n_43520) );
oa12f80 g772637 ( .a(n_8282), .b(n_8289), .c(n_8281), .o(n_9369) );
in01f80 g773032 ( .a(n_7662), .o(n_7686) );
no02f80 g770369 ( .a(n_10582), .b(n_44464), .o(n_10590) );
na02f80 g746275 ( .a(n_34944), .b(n_34550), .o(n_35072) );
ao12f80 g752157 ( .a(n_28226), .b(FE_OCP_RBN2126_n_44734), .c(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .o(n_28088) );
no02f80 g745022 ( .a(n_34795), .b(n_34363), .o(n_34796) );
in01f80 newInst_1379 ( .a(newNet_1378), .o(newNet_1379) );
na02f80 g768063 ( .a(n_13004), .b(n_12223), .o(n_12810) );
in01f80 g748027 ( .a(n_33336), .o(n_33027) );
no02f80 g774047 ( .a(n_7172), .b(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .o(n_7196) );
in01f80 g743318 ( .a(n_36796), .o(n_36797) );
na02f80 g758930 ( .a(n_21394), .b(n_45073), .o(n_21430) );
in01f80 g741102 ( .a(n_39247), .o(n_39248) );
in01f80 newInst_78 ( .a(newNet_77), .o(newNet_78) );
in01f80 g741865 ( .a(n_38368), .o(n_38285) );
in01f80 newInst_2529 ( .a(newNet_1536), .o(newNet_2529) );
in01f80 g737357 ( .a(n_42850), .o(n_42851) );
in01f80 FE_OCP_RBC2942_n_5454 ( .a(n_5454), .o(FE_OCP_RBN2942_n_5454) );
no02f80 g739364 ( .a(n_41052), .b(n_41023), .o(n_41094) );
oa12f80 g777023 ( .a(n_3431), .b(n_3557), .c(n_3556), .o(n_3558) );
na02f80 g740895 ( .a(n_39147), .b(n_39086), .o(n_39310) );
in01f80 g779332 ( .a(n_1658), .o(n_1659) );
in01f80 g776189 ( .a(n_4980), .o(n_4981) );
in01f80 g774190 ( .a(n_6612), .o(n_6613) );
na02f80 g751302 ( .a(n_29638), .b(n_29637), .o(n_29639) );
in01f80 g739928 ( .a(n_40092), .o(n_40123) );
in01f80 newInst_2104 ( .a(newNet_2103), .o(newNet_2104) );
in01f80 g752445 ( .a(n_27799), .o(n_27766) );
na02f80 g756359 ( .a(n_24417), .b(n_23980), .o(n_24453) );
in01f80 g763440 ( .a(n_17042), .o(n_16991) );
in01f80 g780044 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_), .o(n_1381) );
ao12f80 g767465 ( .a(n_13445), .b(n_13444), .c(n_13443), .o(n_13936) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_6_ ( .ck(newNet_880), .d(n_32374), .o(delay_xor_ln21_unr21_stage8_stallmux_q_6_) );
in01f80 newInst_456 ( .a(newNet_455), .o(newNet_456) );
ao22s80 FE_RC_634_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .b(n_6957), .c(n_6585), .d(n_6763), .o(n_6900) );
in01f80 newInst_1131 ( .a(newNet_1130), .o(newNet_1131) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_7_ ( .ck(newNet_3099), .d(n_40439), .o(delay_add_ln22_unr27_stage10_stallmux_q_7_) );
na02f80 g764258 ( .a(n_16722), .b(n_16263), .o(n_16824) );
na02f80 g758676 ( .a(n_21791), .b(FE_OCPN1532_n_21790), .o(n_21815) );
no02f80 FE_RC_34_0 ( .a(FE_RN_6_0), .b(FE_RN_7_0), .o(FE_RN_8_0) );
in01f80 g746173 ( .a(n_33849), .o(n_33826) );
no02f80 g771826 ( .a(n_9775), .b(n_9774), .o(n_9955) );
ao12f80 g749730 ( .a(n_31118), .b(n_31066), .c(n_179), .o(n_31147) );
ao12f80 g738431 ( .a(n_41692), .b(n_41566), .c(n_41564), .o(n_41693) );
oa22f80 FE_RC_1387_0 ( .a(FE_OFN802_n_46285), .b(n_12162), .c(FE_OFN771_n_46337), .d(n_12132), .o(n_46349) );
in01f80 newInst_546 ( .a(newNet_545), .o(newNet_546) );
na02f80 g777262 ( .a(n_3526), .b(n_3525), .o(n_3527) );
in01f80 newInst_3387 ( .a(newNet_3386), .o(newNet_3387) );
no02f80 g775177 ( .a(n_5800), .b(FE_OCPN1028_n_4182), .o(n_5925) );
na02f80 g770468 ( .a(n_10499), .b(n_10402), .o(n_10531) );
in01f80 newInst_388 ( .a(newNet_387), .o(newNet_388) );
oa12f80 g764651 ( .a(FE_OCP_RBN2738_n_15300), .b(n_15772), .c(n_15771), .o(n_15815) );
no02f80 g776439 ( .a(n_4177), .b(n_4203), .o(n_4293) );
in01f80 newInst_1950 ( .a(newNet_1507), .o(newNet_1950) );
no02f80 g753453 ( .a(n_26845), .b(n_25364), .o(n_27192) );
in01f80 g737028 ( .a(n_43033), .o(n_43034) );
na02f80 g773169 ( .a(n_7730), .b(n_7164), .o(n_7827) );
na02f80 g769665 ( .a(n_11273), .b(n_11295), .o(n_11356) );
na02f80 g771463 ( .a(n_9212), .b(n_9136), .o(n_9290) );
no02f80 g780567 ( .a(n_666), .b(FE_OCPN1408_n_672), .o(n_673) );
na02f80 g771212 ( .a(n_9090), .b(n_8362), .o(n_9143) );
in01f80 g764209 ( .a(n_16930), .o(n_16885) );
na02f80 g748882 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .o(n_32454) );
oa22f80 g753805 ( .a(n_27064), .b(n_26900), .c(n_27063), .d(n_26899), .o(n_27107) );
in01f80 g755767 ( .a(n_24484), .o(n_24485) );
in01f80 FE_RC_1039_0 ( .a(n_32855), .o(FE_RN_300_0) );
ao12f80 g777721 ( .a(n_2546), .b(n_3246), .c(n_2522), .o(n_3313) );
na02f80 g748931 ( .a(n_31153), .b(n_31071), .o(n_31180) );
ao22s80 FE_RC_815_0 ( .a(n_42178), .b(n_42176), .c(n_42175), .d(n_42177), .o(n_42194) );
in01f80 newInst_562 ( .a(newNet_159), .o(newNet_562) );
in01f80 newInst_333 ( .a(newNet_332), .o(newNet_333) );
in01f80 g778957 ( .a(n_2247), .o(n_2248) );
in01f80 FE_OCPC3170_n_23227 ( .a(FE_OCPN3169_n_23227), .o(FE_OCPN3170_n_23227) );
na02f80 g757675 ( .a(FE_OCP_RBN1193_n_22542), .b(n_22274), .o(n_22583) );
no02f80 g770893 ( .a(n_10128), .b(n_10163), .o(n_10430) );
in01f80 g761753 ( .a(n_19337), .o(n_19796) );
in01f80 g756052 ( .a(n_25306), .o(n_25284) );
na02f80 g751467 ( .a(n_28549), .b(n_28548), .o(n_28973) );
oa12f80 g752296 ( .a(n_27911), .b(n_45200), .c(FE_OCP_RBN3306_n_44722), .o(n_28036) );
oa12f80 FE_RC_1833_0 ( .a(FE_RN_551_0), .b(n_14190), .c(n_14201), .o(n_14283) );
oa22f80 g741256 ( .a(FE_OCP_RBN2550_n_44944), .b(n_38888), .c(FE_OCPN942_n_44925), .d(n_38469), .o(n_39267) );
no02f80 g738536 ( .a(n_41390), .b(n_41389), .o(n_41452) );
ao12f80 g762838 ( .a(n_17885), .b(n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .o(n_17888) );
oa12f80 g739836 ( .a(n_40253), .b(n_40432), .c(n_39968), .o(n_40446) );
in01f80 g746500 ( .a(n_33341), .o(n_33342) );
no02f80 g765798 ( .a(n_14925), .b(n_14930), .o(n_14975) );
no02f80 g748895 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_10_), .o(n_32411) );
na02f80 g743949 ( .a(n_36306), .b(n_36305), .o(n_36334) );
in01f80 newInst_1791 ( .a(newNet_1790), .o(newNet_1791) );
na02f80 g758768 ( .a(n_21558), .b(n_21557), .o(n_21658) );
in01f80 g768810 ( .a(n_11922), .o(n_11923) );
in01f80 newInst_1907 ( .a(newNet_1906), .o(newNet_1907) );
no02f80 FE_RC_972_0 ( .a(FE_RN_279_0), .b(FE_RN_280_0), .o(FE_RN_281_0) );
no02f80 g745794 ( .a(n_44102), .b(FE_OCP_RBN2323_n_33942), .o(n_34364) );
in01f80 g763864 ( .a(n_16665), .o(n_16666) );
in01f80 newInst_2085 ( .a(newNet_2084), .o(newNet_2085) );
in01f80 g772868 ( .a(n_7985), .o(n_8019) );
na02f80 g764492 ( .a(n_16074), .b(n_14524), .o(n_16202) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_29_ ( .ck(newNet_2731), .d(n_17723), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_) );
ao12f80 g780092 ( .a(n_746), .b(n_1153), .c(n_771), .o(n_1184) );
in01f80 g748650 ( .a(n_31422), .o(n_31423) );
na02f80 g744695 ( .a(n_36555), .b(n_35996), .o(n_36575) );
in01f80 newInst_1193 ( .a(newNet_1192), .o(newNet_1193) );
na02f80 g771446 ( .a(n_9185), .b(FE_OCP_RBN3572_n_44563), .o(n_9345) );
na02f80 g763474 ( .a(n_17541), .b(n_17302), .o(n_17543) );
na02f80 FE_RC_1865_0 ( .a(FE_RN_573_0), .b(n_28183), .o(n_28322) );
ao12f80 g741849 ( .a(n_38364), .b(n_38363), .c(n_38362), .o(n_38495) );
in01f80 g754174 ( .a(n_26020), .o(n_26048) );
na02f80 g766165 ( .a(n_14463), .b(FE_OCP_RBN2253_n_13017), .o(n_14605) );
in01f80 newInst_17 ( .a(newNet_16), .o(newNet_17) );
in01f80 g756283 ( .a(n_24056), .o(n_24057) );
oa12f80 g736271 ( .a(n_289), .b(n_43861), .c(FE_OFN3_n_43918), .o(n_43903) );
no02f80 g756541 ( .a(n_23843), .b(delay_add_ln22_unr14_stage6_stallmux_q_28_), .o(n_23970) );
no02f80 g777613 ( .a(n_3418), .b(n_2682), .o(n_3451) );
oa12f80 g770430 ( .a(n_9811), .b(n_10633), .c(n_9772), .o(n_10687) );
na02f80 g753286 ( .a(n_27110), .b(n_26464), .o(n_27393) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_21_ ( .ck(newNet_1847), .d(n_16925), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_) );
in01f80 g747109 ( .a(n_34019), .o(n_34020) );
in01f80 newInst_242 ( .a(newNet_172), .o(newNet_242) );
no02f80 g766504 ( .a(n_14004), .b(FE_OCPN1420_n_14003), .o(n_14028) );
in01f80 newInst_3670 ( .a(newNet_3669), .o(newNet_3670) );
na02f80 g743894 ( .a(n_36040), .b(n_36038), .o(n_36204) );
in01f80 g752430 ( .a(n_27893), .o(n_27816) );
oa22f80 g758826 ( .a(n_21648), .b(n_21632), .c(n_21705), .d(n_21633), .o(n_21732) );
no02f80 g756047 ( .a(n_25032), .b(n_24627), .o(n_25604) );
in01f80 g754718 ( .a(n_26571), .o(n_26640) );
in01f80 g755075 ( .a(n_25719), .o(n_25720) );
oa12f80 g772985 ( .a(n_7790), .b(n_7789), .c(n_7788), .o(n_7897) );
na02f80 g761186 ( .a(n_19005), .b(n_17815), .o(n_19046) );
na02f80 g770834 ( .a(n_10010), .b(n_9942), .o(n_10090) );
in01f80 FE_RC_1782_0 ( .a(n_28016), .o(FE_RN_520_0) );
na02f80 g755109 ( .a(n_25201), .b(n_25228), .o(n_25321) );
in01f80 g759176 ( .a(n_21348), .o(n_21386) );
in01f80 g748770 ( .a(n_32535), .o(n_32536) );
in01f80 newInst_821 ( .a(newNet_820), .o(newNet_821) );
oa22f80 FE_RC_3869_0 ( .a(n_19238), .b(n_19429), .c(n_19203), .d(n_19428), .o(n_19591) );
oa22f80 g780015 ( .a(n_1259), .b(n_982), .c(n_1264), .d(n_983), .o(n_1272) );
no02f80 g759291 ( .a(n_20804), .b(n_45010), .o(n_20830) );
oa22f80 g746572 ( .a(n_34810), .b(n_34645), .c(n_34666), .d(n_33685), .o(n_35016) );
in01f80 g776355 ( .a(n_4680), .o(n_4681) );
in01f80 g770674 ( .a(n_10310), .o(n_10311) );
in01f80 g767497 ( .a(n_13302), .o(n_13303) );
in01f80 g758152 ( .a(n_23150), .o(n_23151) );
oa22f80 g772392 ( .a(n_8497), .b(n_46418), .c(n_8496), .d(n_8367), .o(n_8597) );
no02f80 g760619 ( .a(n_19856), .b(FE_OCPN1436_n_19855), .o(n_19880) );
in01f80 g778386 ( .a(n_2840), .o(n_2841) );
in01f80 g737073 ( .a(n_43164), .o(n_43200) );
in01f80 g776307 ( .a(n_4830), .o(n_4831) );
in01f80 FE_OCP_RBC3095_n_11413 ( .a(n_11413), .o(FE_OCP_RBN3095_n_11413) );
na02f80 g769096 ( .a(n_11658), .b(n_11657), .o(n_11713) );
in01f80 g750910 ( .a(n_29113), .o(n_29083) );
oa12f80 g743904 ( .a(n_35579), .b(n_35578), .c(n_35577), .o(n_35626) );
in01f80 newInst_33 ( .a(newNet_32), .o(newNet_33) );
in01f80 FE_RC_1123_0 ( .a(n_23322), .o(FE_RN_340_0) );
no02f80 g754110 ( .a(n_26019), .b(n_23339), .o(n_26093) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_24_ ( .ck(newNet_809), .d(n_1336), .o(delay_xor_ln21_unr3_stage2_stallmux_q_24_) );
in01f80 g736802 ( .a(n_43425), .o(n_43426) );
na02f80 g776782 ( .a(n_3740), .b(n_3938), .o(n_3946) );
ao22s80 g736432 ( .a(n_43765), .b(n_43258), .c(n_43764), .d(n_43259), .o(n_43815) );
na02f80 g772239 ( .a(n_8728), .b(FE_OCP_RBN2305_n_7817), .o(n_8799) );
no02f80 g744051 ( .a(n_44222), .b(n_35665), .o(n_35696) );
in01f80 FE_OCP_RBC1841_n_20505 ( .a(n_20505), .o(FE_OCP_RBN1841_n_20505) );
in01f80 newInst_1187 ( .a(newNet_1186), .o(newNet_1187) );
na02f80 g747881 ( .a(n_32142), .b(n_31932), .o(n_32188) );
in01f80 g744270 ( .a(n_35616), .o(n_35587) );
ao22s80 FE_RC_11_0 ( .a(n_1734), .b(n_1539), .c(n_1733), .d(n_1540), .o(n_1822) );
in01f80 g767750 ( .a(n_13238), .o(n_13124) );
in01f80 newInst_532 ( .a(newNet_75), .o(newNet_532) );
in01f80 FE_OCP_RBC2586_n_9009 ( .a(n_9009), .o(FE_OCP_RBN2586_n_9009) );
in01f80 newInst_2568 ( .a(newNet_2567), .o(newNet_2568) );
in01f80 g746725 ( .a(n_34233), .o(n_34234) );
no02f80 g750598 ( .a(n_29371), .b(n_29561), .o(n_29404) );
na02f80 g741588 ( .a(n_38640), .b(n_38635), .o(n_38665) );
in01f80 g759463 ( .a(n_20967), .o(n_20993) );
in01f80 FE_OCPC886_n_42367 ( .a(n_42367), .o(FE_OCPN886_n_42367) );
in01f80 FE_OCP_RBC2146_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2144_FE_OCPN861_n_45450), .o(FE_OCP_RBN2146_FE_OCPN861_n_45450) );
in01f80 g773170 ( .a(n_7839), .o(n_7840) );
in01f80 g752908 ( .a(n_27986), .o(n_27987) );
na02f80 g739462 ( .a(n_44775), .b(n_40761), .o(n_40837) );
ao12f80 g738967 ( .a(n_40978), .b(n_41207), .c(n_40718), .o(n_41270) );
na02f80 g763383 ( .a(FE_OCP_RBN3724_n_16975), .b(n_15901), .o(n_17182) );
in01f80 newInst_288 ( .a(newNet_287), .o(newNet_288) );
in01f80 g764648 ( .a(n_15911), .o(n_16842) );
oa12f80 g737853 ( .a(n_42384), .b(n_42547), .c(n_42350), .o(n_42691) );
in01f80 g744858 ( .a(n_35145), .o(n_35116) );
no02f80 g771176 ( .a(n_9358), .b(n_9416), .o(n_9514) );
in01f80 g748020 ( .a(n_31936), .o(n_31937) );
no02f80 g780831 ( .a(n_542), .b(n_531), .o(n_557) );
na02f80 g780626 ( .a(n_679), .b(n_693), .o(n_703) );
in01f80 g769887 ( .a(n_11081), .o(n_11082) );
oa12f80 g748853 ( .a(n_31196), .b(n_31177), .c(n_31151), .o(n_31353) );
no02f80 g747664 ( .a(n_47205), .b(n_32326), .o(n_32328) );
in01f80 g748507 ( .a(n_31702), .o(n_31716) );
no02f80 g739378 ( .a(n_40816), .b(n_40811), .o(n_41150) );
na02f80 g777749 ( .a(n_3294), .b(n_3322), .o(n_5178) );
na02f80 g757891 ( .a(n_22979), .b(n_22848), .o(n_23026) );
in01f80 FE_OCP_RBC2378_n_29480 ( .a(FE_OCP_RBN2377_n_29480), .o(FE_OCP_RBN2378_n_29480) );
no02f80 g777397 ( .a(n_3559), .b(n_3573), .o(n_3601) );
in01f80 g758242 ( .a(n_22734), .o(n_22652) );
no02f80 g760605 ( .a(n_19754), .b(n_19724), .o(n_19786) );
no02f80 g741787 ( .a(n_38451), .b(n_38450), .o(n_38452) );
oa22f80 g743271 ( .a(n_36738), .b(n_36696), .c(n_36737), .d(n_36677), .o(n_36782) );
in01f80 g766226 ( .a(n_14415), .o(n_14479) );
in01f80 g777013 ( .a(n_3764), .o(n_3765) );
in01f80 g741249 ( .a(n_38983), .o(n_39028) );
no02f80 g745094 ( .a(n_34848), .b(n_34847), .o(n_34849) );
in01f80 g781295 ( .a(n_82), .o(n_55) );
no02f80 g766365 ( .a(n_14124), .b(n_13130), .o(n_14193) );
in01f80 g754913 ( .a(n_25424), .o(n_25425) );
na02f80 g760537 ( .a(n_19936), .b(n_19968), .o(n_20032) );
oa22f80 g757820 ( .a(n_22359), .b(n_22801), .c(n_22317), .d(n_22580), .o(n_22424) );
in01f80 FE_OCP_RBC2178_n_33022 ( .a(n_33022), .o(FE_OCP_RBN2178_n_33022) );
in01f80 FE_OCP_RBC2441_n_8402 ( .a(FE_OCP_RBN2440_n_8402), .o(FE_OCP_RBN2441_n_8402) );
ao12f80 g766514 ( .a(n_13947), .b(n_14027), .c(FE_OCP_RBN2246_n_13017), .o(n_14102) );
ao12f80 g742620 ( .a(n_37526), .b(n_37525), .c(n_37524), .o(n_37619) );
in01f80 g776984 ( .a(n_4044), .o(n_4045) );
na02f80 g753121 ( .a(n_27256), .b(n_27218), .o(n_27300) );
in01f80 g749270 ( .a(n_30869), .o(n_30870) );
in01f80 g738384 ( .a(n_41549), .o(n_41550) );
no03m80 g742698 ( .a(n_37445), .b(n_37410), .c(n_37097), .o(n_37525) );
in01f80 g763307 ( .a(n_17188), .o(n_17189) );
in01f80 FE_RC_3824_0 ( .a(FE_RN_1667_0), .o(FE_RN_1668_0) );
in01f80 g749889 ( .a(n_31490), .o(n_29966) );
in01f80 FE_OCP_RBC2386_n_8342 ( .a(FE_OCP_RBN2384_n_8342), .o(FE_OCP_RBN2386_n_8342) );
na02f80 g745304 ( .a(n_36121), .b(n_36119), .o(n_36169) );
ao22s80 g751082 ( .a(n_28852), .b(n_28570), .c(n_28807), .d(n_28569), .o(n_28888) );
in01f80 newInst_3459 ( .a(newNet_3458), .o(newNet_3459) );
in01f80 g766531 ( .a(n_14026), .o(n_14062) );
in01f80 g762857 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_28_), .o(n_17696) );
in01f80 g745549 ( .a(n_34762), .o(n_34763) );
na02f80 g738136 ( .a(n_42031), .b(n_42023), .o(n_42024) );
in01f80 newInst_1366 ( .a(newNet_1062), .o(newNet_1366) );
na02f80 g759795 ( .a(n_20297), .b(n_20319), .o(n_20417) );
no02f80 g751159 ( .a(n_30097), .b(n_29335), .o(n_30290) );
in01f80 g757022 ( .a(n_24044), .o(n_24074) );
ao12f80 g755460 ( .a(n_25113), .b(n_25262), .c(n_25088), .o(n_25573) );
oa12f80 g764987 ( .a(n_15642), .b(n_15641), .c(n_15640), .o(n_15722) );
na02f80 g742244 ( .a(FE_OCP_RBN2240_n_44881), .b(n_37719), .o(n_38179) );
na02f80 g738193 ( .a(n_41983), .b(n_41982), .o(n_41984) );
oa12f80 g736350 ( .a(n_347), .b(n_43839), .c(n_43918), .o(n_43870) );
no02f80 g738205 ( .a(n_41971), .b(n_41828), .o(n_41989) );
na02f80 g762286 ( .a(n_18446), .b(n_18701), .o(n_18667) );
oa12f80 g782647 ( .a(n_44180), .b(FE_OCP_RBN2645_n_34980), .c(n_35774), .o(n_44040) );
ms00f80 delay_sub_ln23_unr13_stage5_stallmux_q_reg_1_ ( .ck(newNet_1057), .d(n_16887), .o(delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
in01f80 g742583 ( .a(n_37636), .o(n_38668) );
no02f80 g770809 ( .a(n_10135), .b(n_10053), .o(n_10216) );
no02f80 g739352 ( .a(n_40662), .b(n_40461), .o(n_40674) );
in01f80 g772475 ( .a(n_8380), .o(n_8388) );
in01f80 g763546 ( .a(n_16836), .o(n_16912) );
no03m80 FE_RC_628_0 ( .a(n_32704), .b(FE_RN_194_0), .c(n_32672), .o(n_32745) );
na02f80 g743755 ( .a(n_37285), .b(n_46219), .o(n_37328) );
in01f80 newInst_721 ( .a(newNet_720), .o(newNet_721) );
in01f80 g774517 ( .a(n_6765), .o(n_6722) );
in01f80 g738053 ( .a(n_42144), .o(n_42143) );
no02f80 g742214 ( .a(n_44887), .b(n_38273), .o(n_38274) );
no02f80 g742948 ( .a(n_37053), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37164) );
na02f80 g754131 ( .a(n_26053), .b(n_26025), .o(n_26176) );
in01f80 g750466 ( .a(n_30518), .o(n_30519) );
no02f80 g743954 ( .a(n_35669), .b(n_35703), .o(n_35704) );
ao12f80 g770337 ( .a(n_9775), .b(n_10689), .c(n_9870), .o(n_10752) );
in01f80 FE_OCP_RBC2227_n_7598 ( .a(n_7598), .o(FE_OCP_RBN2227_n_7598) );
na02f80 g775705 ( .a(n_5365), .b(n_3993), .o(n_5450) );
no02f80 g764667 ( .a(n_15807), .b(n_15293), .o(n_15906) );
oa12f80 g781262 ( .a(beta_31), .b(beta_16), .c(beta_15), .o(n_75) );
oa12f80 g758913 ( .a(n_21643), .b(n_21642), .c(n_21641), .o(n_21702) );
na02f80 g750087 ( .a(FE_OCP_RBN3561_n_29857), .b(FE_OCP_RBN1906_n_29080), .o(n_29956) );
na02f80 g748635 ( .a(n_31304), .b(FE_OCP_DRV_N3160_n_31303), .o(n_31382) );
na02f80 g755875 ( .a(n_25089), .b(n_25088), .o(n_25346) );
ao12f80 g774121 ( .a(n_7168), .b(n_7172), .c(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .o(n_7198) );
in01f80 g747765 ( .a(n_33758), .o(n_33759) );
no02f80 g781124 ( .a(n_216), .b(n_76), .o(n_223) );
ao12f80 g773393 ( .a(n_7552), .b(n_7551), .c(n_7550), .o(n_8062) );
in01f80 newInst_3433 ( .a(newNet_3432), .o(newNet_3433) );
in01f80 g776892 ( .a(n_5629), .o(n_3994) );
no02f80 g755096 ( .a(n_25180), .b(n_25179), .o(n_25233) );
na02f80 g739982 ( .a(n_39927), .b(n_39876), .o(n_39928) );
na02f80 g772936 ( .a(n_7938), .b(n_7844), .o(n_7845) );
no02f80 g770765 ( .a(FE_OCP_RBN3653_n_10100), .b(FE_OCP_RBN2523_n_8951), .o(n_10290) );
oa12f80 g743857 ( .a(n_35794), .b(n_35793), .c(n_35792), .o(n_35874) );
na02f80 g738422 ( .a(n_41546), .b(n_41545), .o(n_41547) );
in01f80 g780879 ( .a(n_441), .o(n_427) );
in01f80 g753712 ( .a(n_26504), .o(n_26562) );
na02f80 g770816 ( .a(n_9944), .b(FE_OFN755_n_44461), .o(n_10094) );
in01f80 g753490 ( .a(n_26913), .o(n_26914) );
na02f80 g738956 ( .a(n_41235), .b(n_41234), .o(n_41236) );
na02f80 g760000 ( .a(n_20668), .b(FE_OCP_RBN3663_n_20750), .o(n_20751) );
na02f80 g765843 ( .a(n_14906), .b(n_14875), .o(n_14907) );
in01f80 newInst_2021 ( .a(newNet_2020), .o(newNet_2021) );
na02f80 g778070 ( .a(n_3040), .b(n_3039), .o(n_3109) );
no02f80 g758800 ( .a(n_21586), .b(n_45081), .o(n_21615) );
na02f80 g761061 ( .a(n_19119), .b(n_19089), .o(n_19223) );
no02f80 g749482 ( .a(n_30470), .b(n_30471), .o(n_30472) );
na02f80 g744400 ( .a(n_35491), .b(n_35515), .o(n_35551) );
in01f80 newInst_3704 ( .a(newNet_3703), .o(newNet_3704) );
na02f80 g770842 ( .a(n_10052), .b(n_9893), .o(n_10136) );
na02f80 g742055 ( .a(n_37844), .b(FE_OCPN1762_n_37877), .o(n_37895) );
oa12f80 g776001 ( .a(n_5081), .b(n_5080), .c(n_5079), .o(n_5151) );
oa12f80 g764604 ( .a(n_16141), .b(n_16142), .c(n_16140), .o(n_16212) );
na02f80 g749409 ( .a(n_30603), .b(n_30295), .o(n_30624) );
na02f80 g750076 ( .a(n_29896), .b(n_30192), .o(n_30216) );
no03m80 g750521 ( .a(n_30001), .b(n_30442), .c(n_29877), .o(n_30549) );
na02f80 g778674 ( .a(n_2256), .b(n_2255), .o(n_2306) );
in01f80 g748428 ( .a(n_31681), .o(n_31703) );
no02f80 g743028 ( .a(n_36990), .b(n_36989), .o(n_37197) );
no02f80 g742207 ( .a(n_44867), .b(n_37882), .o(n_37883) );
na02f80 g768658 ( .a(n_12195), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_), .o(n_12294) );
oa22f80 FE_RC_1587_0 ( .a(FE_OFN802_n_46285), .b(n_12197), .c(FE_OFN771_n_46337), .d(n_12116), .o(n_46350) );
ao12f80 g754369 ( .a(n_25422), .b(FE_OCP_RBN2764_n_25732), .c(n_25760), .o(n_25785) );
in01f80 FE_OCP_RBC2823_n_10068 ( .a(n_10068), .o(FE_OCP_RBN2823_n_10068) );
no02f80 g763295 ( .a(n_17326), .b(n_17325), .o(n_17327) );
na02f80 g740730 ( .a(n_39357), .b(n_39259), .o(n_39446) );
no02f80 g764951 ( .a(n_15472), .b(n_14215), .o(n_15474) );
no02f80 g780863 ( .a(n_532), .b(n_526), .o(n_1045) );
na02f80 g757442 ( .a(FE_OCP_RBN2152_n_22822), .b(n_22931), .o(n_22988) );
na02f80 g779191 ( .a(n_1839), .b(n_1729), .o(n_1921) );
no02f80 g750371 ( .a(n_29687), .b(n_29669), .o(n_29670) );
in01f80 g741121 ( .a(n_39272), .o(n_39273) );
no02f80 FE_RC_2656_0 ( .a(FE_RN_1109_0), .b(n_12582), .o(n_12641) );
ao22s80 FE_RC_2806_0 ( .a(n_13211), .b(n_13709), .c(n_13212), .d(n_13695), .o(n_13818) );
in01f80 FE_RC_2715_0 ( .a(n_23186), .o(FE_RN_1145_0) );
na02f80 g739265 ( .a(n_40764), .b(n_44769), .o(n_40855) );
na02f80 g749546 ( .a(n_30354), .b(n_30176), .o(n_30409) );
in01f80 g741704 ( .a(n_39040), .o(n_38538) );
in01f80 newInst_2392 ( .a(newNet_2391), .o(newNet_2392) );
na02f80 g740137 ( .a(n_39770), .b(n_39785), .o(n_39802) );
in01f80 newInst_3441 ( .a(newNet_3440), .o(newNet_3441) );
no02f80 g767696 ( .a(n_13160), .b(n_13241), .o(n_13242) );
in01f80 g773492 ( .a(n_7498), .o(n_7499) );
no02f80 FE_RC_3128_0 ( .a(n_30703), .b(n_30944), .o(FE_RN_1386_0) );
no02f80 g742893 ( .a(n_37005), .b(n_37019), .o(n_37419) );
in01f80 g742808 ( .a(n_37258), .o(n_37272) );
na02f80 g768367 ( .a(n_12524), .b(n_11101), .o(n_12583) );
na02f80 g738169 ( .a(n_41999), .b(n_41998), .o(n_42000) );
na02f80 FE_RC_2797_0 ( .a(FE_RN_1195_0), .b(n_44104), .o(FE_RN_1196_0) );
oa12f80 g740986 ( .a(n_38876), .b(n_39107), .c(n_38957), .o(n_39137) );
in01f80 g774774 ( .a(n_6476), .o(n_6436) );
na02f80 g773060 ( .a(n_45826), .b(n_7647), .o(n_7745) );
in01f80 fopt782683 ( .a(FE_OCP_RBN3819_n_44061), .o(n_44084) );
ao12f80 g739930 ( .a(n_39928), .b(n_39959), .c(n_39873), .o(n_40050) );
no02f80 g756722 ( .a(n_24036), .b(n_24007), .o(n_24008) );
no02f80 g740572 ( .a(n_39614), .b(n_45840), .o(n_39647) );
no02f80 g746862 ( .a(n_34107), .b(n_34106), .o(n_34108) );
na02f80 g773914 ( .a(n_7063), .b(n_7062), .o(n_7138) );
na02f80 g762062 ( .a(n_18930), .b(n_18836), .o(n_18963) );
in01f80 g741845 ( .a(n_38469), .o(n_38888) );
in01f80 g744799 ( .a(n_35223), .o(n_35171) );
in01f80 FE_OCP_RBC2173_n_1813 ( .a(n_1813), .o(FE_OCP_RBN2173_n_1813) );
ao22s80 FE_RC_156_0 ( .a(FE_OCPN3773_n_15371), .b(n_15805), .c(n_15372), .d(n_15852), .o(n_16041) );
in01f80 FE_OCP_RBC1214_n_31847 ( .a(n_31847), .o(FE_OCP_RBN1214_n_31847) );
in01f80 FE_OCPC861_n_45450 ( .a(n_45450), .o(FE_OCPN861_n_45450) );
ao12f80 g774200 ( .a(n_7033), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .o(n_7119) );
in01f80 g759910 ( .a(n_21107), .o(n_21108) );
na02f80 g748148 ( .a(n_32138), .b(n_32072), .o(n_32161) );
ao22s80 FE_RC_1068_0 ( .a(n_37450), .b(n_37181), .c(n_37180), .d(n_37449), .o(n_37535) );
in01f80 newInst_2290 ( .a(newNet_2289), .o(newNet_2290) );
na02f80 g736962 ( .a(n_43242), .b(n_42969), .o(n_43456) );
in01f80 g744946 ( .a(n_35001), .o(n_35000) );
no02f80 g756915 ( .a(n_23347), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .o(n_23361) );
in01f80 g756069 ( .a(n_24979), .o(n_25304) );
no02f80 g780726 ( .a(n_619), .b(n_614), .o(n_615) );
na02f80 g766600 ( .a(n_14354), .b(n_14433), .o(n_14434) );
in01f80 newInst_3175 ( .a(newNet_3174), .o(newNet_3175) );
in01f80 g779734 ( .a(n_1407), .o(n_1408) );
na02f80 g742061 ( .a(FE_OCP_RBN3448_n_37945), .b(n_37912), .o(n_38281) );
no02f80 g743978 ( .a(n_36531), .b(n_35003), .o(n_36146) );
in01f80 newInst_1732 ( .a(newNet_1731), .o(newNet_1732) );
no02f80 g756390 ( .a(n_23946), .b(n_23774), .o(n_23973) );
na02f80 g754021 ( .a(FE_OCP_RBN1204_n_26121), .b(n_26178), .o(n_26206) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_27_ ( .ck(newNet_3511), .d(n_22903), .o(delay_add_ln22_unr14_stage6_stallmux_q_27_) );
no02f80 g742716 ( .a(n_37323), .b(n_37322), .o(n_37324) );
in01f80 g752264 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_8_), .o(n_27869) );
in01f80 g737617 ( .a(n_42400), .o(n_42401) );
na02f80 g738504 ( .a(FE_OCP_RBN2316_n_41420), .b(n_41543), .o(n_41638) );
no02f80 FE_RC_2540_0 ( .a(n_38953), .b(n_38901), .o(FE_RN_1037_0) );
ao12f80 FE_RC_3130_0 ( .a(FE_RN_1386_0), .b(FE_RN_1387_0), .c(n_30862), .o(n_31003) );
no02f80 g778060 ( .a(n_3041), .b(n_2784), .o(n_3042) );
oa12f80 g750665 ( .a(n_28789), .b(n_29237), .c(n_28787), .o(n_29343) );
na02f80 FE_RC_2503_0 ( .a(n_7827), .b(n_7805), .o(FE_RN_1016_0) );
ao12f80 g770261 ( .a(n_10463), .b(n_10740), .c(n_46420), .o(n_10779) );
oa12f80 g765175 ( .a(n_14927), .b(n_15023), .c(n_14877), .o(n_15124) );
in01f80 g751334 ( .a(n_29999), .o(n_29535) );
in01f80 FE_RC_3150_0 ( .a(n_20874), .o(FE_RN_1398_0) );
no02f80 g745812 ( .a(n_44102), .b(n_34143), .o(n_34522) );
in01f80 newInst_2826 ( .a(newNet_2825), .o(newNet_2826) );
in01f80 newInst_3018 ( .a(newNet_3017), .o(newNet_3018) );
na02f80 g778045 ( .a(n_3101), .b(n_3329), .o(n_3104) );
in01f80 newInst_60 ( .a(newNet_36), .o(newNet_60) );
na02f80 g762205 ( .a(n_18813), .b(n_18624), .o(n_19680) );
no02f80 g776491 ( .a(n_4487), .b(n_4350), .o(n_4488) );
in01f80 g751970 ( .a(n_29025), .o(n_29308) );
no02f80 g753790 ( .a(n_27097), .b(n_26642), .o(n_27135) );
in01f80 g744020 ( .a(n_36899), .o(n_36900) );
oa22f80 FE_RC_1237_0 ( .a(FE_OFN84_n_46137), .b(n_6618), .c(FE_OFN806_n_46196), .d(n_6648), .o(n_46188) );
no02f80 g736587 ( .a(n_43657), .b(n_43431), .o(n_43682) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_6_ ( .ck(newNet_1365), .d(n_36286), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_) );
na02f80 g737071 ( .a(n_43082), .b(n_46937), .o(n_43189) );
in01f80 g739877 ( .a(n_40380), .o(n_40432) );
in01f80 newInst_2884 ( .a(newNet_2883), .o(newNet_2884) );
in01f80 g779099 ( .a(n_2017), .o(n_2018) );
na02f80 FE_RC_3028_0 ( .a(FE_OCP_RBN2740_n_20565), .b(FE_RN_1326_0), .o(n_21149) );
no02f80 g739823 ( .a(n_40431), .b(n_40308), .o(n_40453) );
na02f80 g746620 ( .a(n_34473), .b(n_34523), .o(n_34638) );
in01f80 g758089 ( .a(n_22263), .o(n_22264) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_17_ ( .ck(newNet_1020), .d(n_17880), .o(delay_xor_ln21_unr12_stage5_stallmux_q_17_) );
in01f80 g771294 ( .a(n_9555), .o(n_9613) );
in01f80 g736931 ( .a(n_43062), .o(n_43085) );
ao22s80 FE_RC_1350_0 ( .a(n_4880), .b(n_4816), .c(n_4815), .d(n_4881), .o(n_5049) );
na02f80 g774509 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_27_), .o(n_6703) );
na02f80 g773466 ( .a(n_7534), .b(n_7523), .o(n_7524) );
in01f80 g736791 ( .a(n_43068), .o(n_43069) );
no02f80 g771966 ( .a(FE_OCP_RBN3647_n_44490), .b(n_9647), .o(n_9770) );
no02f80 g779091 ( .a(n_2051), .b(n_2050), .o(n_2052) );
oa12f80 g740698 ( .a(n_39079), .b(n_39414), .c(n_38987), .o(n_39475) );
na02f80 g767052 ( .a(FE_OCP_RBN2458_n_13765), .b(n_13875), .o(n_13898) );
no02f80 g770110 ( .a(n_10771), .b(n_10738), .o(n_10852) );
ao12f80 g746371 ( .a(n_33521), .b(n_33520), .c(n_33519), .o(n_33613) );
in01f80 g771561 ( .a(FE_OCP_RBN2544_n_9082), .o(n_10733) );
no02f80 g768053 ( .a(FE_OCPN860_n_12880), .b(n_12325), .o(n_13197) );
in01f80 g749241 ( .a(n_32116), .o(n_32154) );
no02f80 g737742 ( .a(n_42394), .b(n_42159), .o(n_42470) );
in01f80 FE_OCP_RBC3637_n_44490 ( .a(n_44490), .o(FE_OCP_RBN3637_n_44490) );
ao22s80 FE_RC_2977_0 ( .a(n_35139), .b(n_35332), .c(FE_OCP_RBN2682_n_35139), .d(n_35319), .o(n_35416) );
no02f80 g743885 ( .a(n_35914), .b(n_35698), .o(n_35955) );
in01f80 g766405 ( .a(n_14317), .o(n_14396) );
oa12f80 g770652 ( .a(n_9935), .b(n_9898), .c(n_9933), .o(n_10021) );
no02f80 g749750 ( .a(n_31091), .b(n_31090), .o(n_31092) );
no02f80 g761967 ( .a(n_18300), .b(n_18285), .o(n_18316) );
in01f80 newInst_2016 ( .a(newNet_2015), .o(newNet_2016) );
in01f80 newInst_1339 ( .a(newNet_1338), .o(newNet_1339) );
na02f80 g771883 ( .a(n_8838), .b(FE_OCPN917_n_46991), .o(n_8862) );
in01f80 g738740 ( .a(n_41527), .o(n_41528) );
in01f80 newInst_1145 ( .a(newNet_249), .o(newNet_1145) );
in01f80 newInst_520 ( .a(newNet_519), .o(newNet_520) );
no02f80 g763673 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .o(n_17575) );
in01f80 FE_OCP_RBC3551_n_44575 ( .a(FE_OCP_RBN3545_n_44575), .o(FE_OCP_RBN3551_n_44575) );
no02f80 g766881 ( .a(n_14303), .b(FE_OCP_RBN2506_n_13896), .o(n_14421) );
in01f80 g744951 ( .a(n_35046), .o(n_35047) );
na02f80 g781023 ( .a(cos_out_11), .b(FE_OFN2_n_43918), .o(n_303) );
no02f80 g766327 ( .a(n_14187), .b(n_14229), .o(n_14330) );
oa22f80 FE_RC_578_0 ( .a(n_42044), .b(n_41764), .c(n_42043), .d(n_41765), .o(n_42122) );
no02f80 g749134 ( .a(n_30910), .b(FE_OCPN1490_n_30823), .o(n_30911) );
in01f80 FE_OCP_RBC3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_ ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
in01f80 g759659 ( .a(n_20510), .o(n_20555) );
na02f80 FE_RC_3542_0 ( .a(FE_RN_1531_0), .b(FE_RN_1533_0), .o(FE_RN_1534_0) );
in01f80 FE_OCP_RBC3555_n_44575 ( .a(FE_OCP_RBN3553_n_44575), .o(FE_OCP_RBN3555_n_44575) );
in01f80 g773703 ( .a(n_7337), .o(n_7338) );
na02f80 g781060 ( .a(cos_out_10), .b(FE_OFN2_n_43918), .o(n_330) );
na02f80 g737924 ( .a(n_42270), .b(n_42500), .o(n_42580) );
na02f80 g762824 ( .a(n_17801), .b(n_17800), .o(n_17870) );
no02f80 g757496 ( .a(n_23357), .b(n_23356), .o(n_23358) );
no02f80 g777671 ( .a(n_3357), .b(n_3346), .o(n_3414) );
oa12f80 g743293 ( .a(n_37923), .b(n_37922), .c(n_46247), .o(n_38019) );
na02f80 g772852 ( .a(n_7967), .b(n_8752), .o(n_8008) );
oa22f80 FE_RC_3814_0 ( .a(n_12659), .b(n_13062), .c(n_12660), .d(n_13008), .o(n_13228) );
in01f80 g738799 ( .a(n_41491), .o(n_41537) );
na02f80 FE_RC_2616_0 ( .a(n_14587), .b(FE_RN_1089_0), .o(n_14673) );
no02f80 g759365 ( .a(n_21115), .b(n_21174), .o(n_21257) );
na02f80 FE_RC_3837_0 ( .a(n_44061), .b(FE_RN_1672_0), .o(n_22708) );
in01f80 g773301 ( .a(FE_OCP_RBN3475_n_7886), .o(n_9012) );
ao22s80 FE_RC_3919_0 ( .a(n_32134), .b(n_45754), .c(n_45755), .d(n_32135), .o(n_32395) );
na02f80 g774741 ( .a(n_6395), .b(n_6394), .o(n_6408) );
na02f80 g761085 ( .a(n_19990), .b(n_20041), .o(n_20042) );
na02f80 g756502 ( .a(n_23633), .b(n_23659), .o(n_23731) );
no02f80 g750449 ( .a(n_30518), .b(n_30066), .o(n_30551) );
in01f80 g765369 ( .a(n_16249), .o(n_16250) );
in01f80 g764711 ( .a(n_15861), .o(n_15901) );
in01f80 g754082 ( .a(n_26129), .o(n_26104) );
na02f80 g740515 ( .a(n_39746), .b(n_39745), .o(n_39774) );
in01f80 FE_OCP_RBC3606_n_8981 ( .a(FE_OCP_RBN3605_n_8981), .o(FE_OCP_RBN3606_n_8981) );
in01f80 FE_OFC826_n_1142 ( .a(n_1142), .o(FE_OFN826_n_1142) );
no02f80 g740943 ( .a(n_39282), .b(n_39162), .o(n_39335) );
na02f80 g758938 ( .a(n_21700), .b(n_21604), .o(n_21701) );
no02f80 g755999 ( .a(n_25160), .b(n_25109), .o(n_25521) );
in01f80 g779732 ( .a(n_1521), .o(n_1559) );
na02f80 g777360 ( .a(n_4759), .b(n_3471), .o(n_5330) );
in01f80 g754414 ( .a(n_25758), .o(n_25759) );
na02f80 FE_RC_4100_0 ( .a(FE_RN_1792_0), .b(FE_RN_1793_0), .o(FE_RN_1794_0) );
oa12f80 g770785 ( .a(n_10034), .b(n_10182), .c(n_9959), .o(n_10223) );
no02f80 g748561 ( .a(n_31386), .b(n_31202), .o(n_31449) );
na02f80 g757338 ( .a(n_23106), .b(n_44071), .o(n_23129) );
in01f80 newInst_347 ( .a(newNet_346), .o(newNet_347) );
na02f80 g740259 ( .a(n_39964), .b(n_39992), .o(n_39993) );
ao12f80 g778160 ( .a(n_2854), .b(n_2853), .c(n_2852), .o(n_4437) );
no02f80 g778457 ( .a(n_2415), .b(n_2401), .o(n_2511) );
in01f80 g767148 ( .a(n_14420), .o(n_14524) );
in01f80 g737629 ( .a(n_42644), .o(n_42645) );
in01f80 newInst_1831 ( .a(newNet_542), .o(newNet_1831) );
ao22s80 FE_RC_4021_0 ( .a(n_15349), .b(n_15309), .c(n_15313), .d(n_15308), .o(n_15610) );
in01f80 newInst_2646 ( .a(newNet_2645), .o(newNet_2646) );
ao22s80 g761386 ( .a(n_19787), .b(n_18886), .c(n_19980), .d(n_19913), .o(n_20114) );
in01f80 g771547 ( .a(n_9046), .o(n_9083) );
no02f80 g736764 ( .a(n_43272), .b(n_43271), .o(n_43321) );
na02f80 FE_RC_2785_0 ( .a(n_18230), .b(FE_OCP_RBN3510_n_19599), .o(FE_RN_1189_0) );
in01f80 g758878 ( .a(n_21442), .o(n_21443) );
oa22f80 g750041 ( .a(n_29869), .b(FE_OCP_RBN2376_n_29480), .c(n_29896), .d(n_29523), .o(n_30345) );
in01f80 g738901 ( .a(n_41299), .o(n_41590) );
na02f80 g776098 ( .a(n_4946), .b(n_4595), .o(n_5064) );
in01f80 FE_OCP_RBC3825_n_18951 ( .a(n_18951), .o(FE_OCP_RBN3825_n_18951) );
na02f80 g777180 ( .a(n_5330), .b(n_5297), .o(n_5380) );
na02f80 g744576 ( .a(n_35383), .b(n_35382), .o(n_35418) );
na02f80 g778660 ( .a(n_2386), .b(n_2385), .o(n_2425) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_14_ ( .ck(newNet_744), .d(n_46155), .o(delay_xor_ln21_unr6_stage3_stallmux_q_14_) );
no02f80 g740194 ( .a(FE_OCP_RBN3056_n_39913), .b(n_39822), .o(n_40217) );
no02f80 g756603 ( .a(n_23561), .b(n_23560), .o(n_23580) );
in01f80 newInst_435 ( .a(newNet_241), .o(newNet_435) );
na02f80 g775823 ( .a(n_5163), .b(n_4182), .o(n_5251) );
no02f80 g774375 ( .a(n_6658), .b(n_6592), .o(n_7229) );
in01f80 newInst_465 ( .a(newNet_464), .o(newNet_465) );
na02f80 g742053 ( .a(n_37945), .b(n_37495), .o(n_37975) );
oa22f80 FE_RC_3671_0 ( .a(n_27482), .b(n_27684), .c(n_27483), .d(n_27703), .o(n_27800) );
in01f80 newInst_2533 ( .a(newNet_2321), .o(newNet_2533) );
na02f80 g744886 ( .a(n_34934), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34961) );
no02f80 g746797 ( .a(n_32897), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n_32922) );
na02f80 g768343 ( .a(n_12469), .b(n_12468), .o(n_12522) );
na02f80 g767522 ( .a(n_13096), .b(n_13095), .o(n_13142) );
in01f80 g762744 ( .a(n_17872), .o(n_17873) );
in01f80 FE_OCP_RBC2311_n_41420 ( .a(n_41420), .o(FE_OCP_RBN2311_n_41420) );
na02f80 g773139 ( .a(n_7712), .b(n_7663), .o(n_7751) );
oa12f80 g761643 ( .a(n_19493), .b(n_19492), .c(n_19491), .o(n_19794) );
in01f80 g771442 ( .a(n_9406), .o(n_9407) );
no02f80 g737458 ( .a(n_42715), .b(n_42702), .o(n_42792) );
in01f80 g759387 ( .a(n_21064), .o(n_21065) );
oa12f80 g738310 ( .a(n_41834), .b(n_41833), .c(n_41832), .o(n_41916) );
in01f80 g770907 ( .a(n_9930), .o(n_9931) );
in01f80 FE_OCP_RBC3675_FE_RN_1581_0 ( .a(FE_RN_1581_0), .o(FE_OCP_RBN3675_FE_RN_1581_0) );
ao12f80 g779379 ( .a(n_1546), .b(n_1551), .c(n_1545), .o(n_2234) );
no02f80 g767762 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_), .o(n_13319) );
na02f80 g742132 ( .a(n_38297), .b(n_38277), .o(n_38409) );
in01f80 newInst_712 ( .a(newNet_711), .o(newNet_712) );
in01f80 g776493 ( .a(n_4476), .o(n_4477) );
in01f80 g740858 ( .a(n_39401), .o(n_39402) );
in01f80 g775964 ( .a(n_5149), .o(n_5177) );
ao12f80 g779511 ( .a(n_1971), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .o(n_1983) );
oa12f80 g776128 ( .a(n_4912), .b(n_4911), .c(n_4910), .o(n_4987) );
oa12f80 g763034 ( .a(n_17121), .b(n_17452), .c(n_17451), .o(n_17492) );
in01f80 FE_OCP_RBC3563_n_29857 ( .a(n_29857), .o(FE_OCP_RBN3563_n_29857) );
na02f80 g746583 ( .a(n_34810), .b(n_34802), .o(n_34938) );
no02f80 g747222 ( .a(n_32787), .b(n_32817), .o(n_32849) );
in01f80 g775262 ( .a(n_5972), .o(n_5937) );
ao12f80 g751625 ( .a(n_28370), .b(n_28391), .c(n_28369), .o(n_29573) );
na02f80 g780067 ( .a(n_1222), .b(n_769), .o(n_1225) );
na02f80 g763934 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .o(n_17152) );
in01f80 g761896 ( .a(n_18912), .o(n_18913) );
no02f80 g746024 ( .a(n_33942), .b(n_34037), .o(n_33961) );
in01f80 newInst_1569 ( .a(newNet_490), .o(newNet_1569) );
ao12f80 g764388 ( .a(n_15866), .b(n_16615), .c(n_15925), .o(n_16675) );
ao12f80 g781151 ( .a(n_57), .b(n_199), .c(n_101), .o(n_202) );
no02f80 g742389 ( .a(n_37771), .b(n_37770), .o(n_37808) );
in01f80 newInst_1117 ( .a(newNet_79), .o(newNet_1117) );
no02f80 g762654 ( .a(n_45528), .b(n_17607), .o(n_18294) );
in01f80 g769324 ( .a(n_11970), .o(n_11971) );
oa12f80 g776830 ( .a(n_2874), .b(n_3600), .c(n_2818), .o(n_3737) );
na02f80 g766278 ( .a(n_14332), .b(n_14370), .o(n_14407) );
in01f80 g762324 ( .a(n_18128), .o(n_18129) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_2_ ( .ck(newNet_2159), .d(n_1021), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_25_ ( .ck(newNet_1500), .d(n_32294), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_) );
no02f80 g740611 ( .a(FE_OCP_RBN2865_n_39640), .b(n_39638), .o(n_39735) );
no02f80 g760964 ( .a(n_19223), .b(n_19222), .o(n_19224) );
in01f80 g770353 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(n_12164) );
no02f80 g770102 ( .a(n_10702), .b(n_10674), .o(n_10797) );
no02f80 g756865 ( .a(n_24075), .b(n_24105), .o(n_24106) );
in01f80 g773191 ( .a(n_8036), .o(n_8037) );
oa12f80 g767251 ( .a(n_13542), .b(n_13541), .c(n_13540), .o(n_15337) );
in01f80 newInst_3340 ( .a(newNet_3339), .o(newNet_3340) );
na02f80 g774955 ( .a(n_6135), .b(FE_OCP_RBN2924_n_5130), .o(n_6197) );
in01f80 FE_RC_3749_0 ( .a(n_11983), .o(FE_RN_1645_0) );
na02f80 g758033 ( .a(n_22219), .b(n_22259), .o(n_22377) );
ao22s80 g737309 ( .a(n_42842), .b(n_42642), .c(n_42852), .d(n_42641), .o(n_43123) );
in01f80 g752323 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_8_), .o(n_27913) );
no02f80 g747196 ( .a(n_33890), .b(n_33889), .o(n_33891) );
in01f80 g742186 ( .a(n_38231), .o(n_38232) );
na02f80 g780766 ( .a(n_505), .b(n_408), .o(n_523) );
oa22f80 g759802 ( .a(n_21691), .b(n_21454), .c(n_21714), .d(n_20179), .o(n_21880) );
in01f80 g780154 ( .a(n_1164), .o(n_1157) );
na02f80 g772669 ( .a(n_8255), .b(n_8224), .o(n_8225) );
na02f80 g754015 ( .a(n_26140), .b(n_26103), .o(n_26180) );
in01f80 newInst_2975 ( .a(newNet_2974), .o(newNet_2975) );
na02f80 FE_RC_1730_0 ( .a(FE_RN_478_0), .b(FE_RN_480_0), .o(n_23579) );
in01f80 g747277 ( .a(n_33722), .o(n_33723) );
no02f80 g746416 ( .a(n_33429), .b(n_32935), .o(n_33458) );
in01f80 FE_RC_2884_0 ( .a(FE_OCP_RBN1159_n_18517), .o(FE_RN_1248_0) );
in01f80 g771838 ( .a(n_9813), .o(n_9814) );
ao12f80 g754945 ( .a(n_25647), .b(n_25552), .c(n_25551), .o(n_25668) );
in01f80 FE_OFC360_n_9391 ( .a(n_9391), .o(FE_OFN360_n_9391) );
in01f80 FE_RC_2707_0 ( .a(FE_RN_1139_0), .o(n_8440) );
in01f80 g737662 ( .a(n_42583), .o(n_42584) );
na02f80 g740178 ( .a(FE_OCP_RBN3715_n_39913), .b(n_39580), .o(n_40071) );
no02f80 g777017 ( .a(n_3846), .b(n_3742), .o(n_3853) );
oa22f80 g748697 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_), .c(n_32587), .d(n_32496), .o(n_32588) );
in01f80 newInst_2769 ( .a(newNet_2207), .o(newNet_2769) );
na02f80 g771944 ( .a(n_8803), .b(FE_OCP_RBN2304_n_7817), .o(n_8804) );
no02f80 g769110 ( .a(n_11620), .b(n_11584), .o(n_11749) );
na02f80 g747810 ( .a(n_33392), .b(n_33512), .o(n_33817) );
na02f80 g778698 ( .a(n_2235), .b(n_2766), .o(n_2233) );
oa22f80 g770545 ( .a(FE_OCP_RBN2794_n_10106), .b(n_10484), .c(FE_OCP_RBN3666_n_10106), .d(n_8937), .o(n_10363) );
in01f80 FE_RC_1927_0 ( .a(n_28764), .o(FE_RN_610_0) );
in01f80 fopt783276 ( .a(n_44849), .o(n_44850) );
in01f80 g747002 ( .a(n_33012), .o(n_33013) );
no02f80 g754926 ( .a(n_25542), .b(n_24959), .o(n_25672) );
in01f80 FE_OCP_RBC2980_n_5656 ( .a(n_5656), .o(FE_OCP_RBN2980_n_5656) );
ao22s80 g777039 ( .a(FE_OCP_RBN2583_n_3734), .b(FE_OCP_RBN3587_n_47016), .c(n_3700), .d(n_47016), .o(n_4014) );
na03f80 g737725 ( .a(n_42296), .b(n_42363), .c(n_42362), .o(n_42387) );
in01f80 g757503 ( .a(n_23029), .o(n_23030) );
in01f80 newInst_2346 ( .a(newNet_2345), .o(newNet_2346) );
in01f80 newInst_931 ( .a(newNet_930), .o(newNet_931) );
in01f80 g757833 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_15_), .o(n_23554) );
in01f80 newInst_393 ( .a(newNet_392), .o(newNet_393) );
ao12f80 g776403 ( .a(n_4589), .b(n_4710), .c(n_4492), .o(n_4827) );
in01f80 FE_RC_505_0 ( .a(n_45311), .o(FE_RN_154_0) );
in01f80 FE_OCP_RBC2923_n_5130 ( .a(FE_OCP_RBN3688_n_5130), .o(FE_OCP_RBN2923_n_5130) );
no02f80 g743198 ( .a(n_36908), .b(n_36906), .o(n_36907) );
no02f80 g740249 ( .a(n_39937), .b(n_39880), .o(n_39938) );
no02f80 g753967 ( .a(n_26240), .b(n_23564), .o(n_26281) );
no02f80 g778099 ( .a(n_2987), .b(n_2833), .o(n_2972) );
no02f80 g751554 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n_28566) );
in01f80 g736347 ( .a(n_43825), .o(n_43826) );
no02f80 g736530 ( .a(n_43686), .b(n_43276), .o(n_43699) );
no02f80 FE_RC_1637_0 ( .a(n_11992), .b(FE_RN_455_0), .o(n_12129) );
na02f80 g768457 ( .a(n_12350), .b(delay_add_ln22_unr8_stage4_stallmux_q_10_), .o(n_12391) );
in01f80 fopt783517 ( .a(n_18421), .o(n_45120) );
ao12f80 g754475 ( .a(n_25519), .b(n_25518), .c(n_25517), .o(n_25598) );
no02f80 g776249 ( .a(n_4792), .b(FE_OCP_RBN2578_n_47017), .o(n_4825) );
no02f80 g751487 ( .a(n_28505), .b(n_28451), .o(n_28832) );
no02f80 g760356 ( .a(n_20203), .b(n_20183), .o(n_20225) );
in01f80 g762647 ( .a(n_18039), .o(n_18040) );
no02f80 g755513 ( .a(n_24723), .b(n_24686), .o(n_24799) );
na02f80 g780448 ( .a(n_764), .b(n_46055), .o(n_935) );
no02f80 g775735 ( .a(n_5461), .b(n_4041), .o(n_5709) );
ao12f80 g751076 ( .a(n_29909), .b(n_30095), .c(n_29756), .o(n_30124) );
in01f80 FE_RC_2256_0 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(FE_RN_833_0) );
in01f80 g736758 ( .a(n_43220), .o(n_43221) );
oa12f80 g772775 ( .a(n_8054), .b(n_8057), .c(n_8006), .o(n_8197) );
in01f80 g767691 ( .a(n_12935), .o(n_12936) );
na02f80 g761769 ( .a(n_19229), .b(n_19228), .o(n_19230) );
no02f80 g751840 ( .a(n_29128), .b(n_29069), .o(n_29760) );
in01f80 g742023 ( .a(n_38034), .o(n_38035) );
na02f80 g754697 ( .a(FE_OCP_RBN2960_n_26231), .b(n_25547), .o(n_26865) );
in01f80 g737127 ( .a(FE_OCP_RBN3699_n_43015), .o(n_43038) );
no02f80 g757963 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n_23057) );
oa12f80 g746046 ( .a(n_34644), .b(n_35190), .c(n_35069), .o(n_35246) );
in01f80 newInst_2137 ( .a(newNet_2136), .o(newNet_2137) );
no02f80 g760060 ( .a(n_20316), .b(FE_OCP_RBN3846_FE_RN_1242_0), .o(n_20376) );
na02f80 FE_RC_4009_0 ( .a(FE_RN_1740_0), .b(n_20501), .o(n_20612) );
in01f80 g766665 ( .a(n_13815), .o(n_13866) );
oa12f80 g745085 ( .a(n_34791), .b(n_34790), .c(n_34789), .o(n_34870) );
no02f80 g761192 ( .a(n_19957), .b(n_20014), .o(n_20015) );
no02f80 g756913 ( .a(n_23384), .b(n_23391), .o(n_23385) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_18_ ( .ck(newNet_348), .d(n_1311), .o(delay_xor_ln22_unr3_stage2_stallmux_q_18_) );
no02f80 g765514 ( .a(n_15514), .b(n_15669), .o(n_15787) );
na02f80 g738294 ( .a(n_41865), .b(n_41864), .o(n_41866) );
in01f80 newInst_325 ( .a(newNet_262), .o(newNet_325) );
in01f80 newInst_3215 ( .a(newNet_3214), .o(newNet_3215) );
in01f80 g771387 ( .a(n_9152), .o(n_9266) );
na02f80 g770966 ( .a(n_9579), .b(n_9541), .o(n_9626) );
in01f80 g742177 ( .a(n_38303), .o(n_38304) );
no02f80 g742478 ( .a(n_37646), .b(n_37645), .o(n_37693) );
no02f80 g753600 ( .a(n_26666), .b(n_26665), .o(n_26748) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_1_ ( .ck(newNet_3146), .d(n_39786), .o(delay_add_ln22_unr27_stage10_stallmux_q_1_) );
no02f80 g740051 ( .a(n_40016), .b(n_40015), .o(n_40017) );
ao12f80 g777135 ( .a(n_4371), .b(n_4215), .c(n_4261), .o(n_4372) );
in01f80 g736316 ( .a(n_43874), .o(n_43875) );
no02f80 g755823 ( .a(FE_OCP_RBN2335_n_24359), .b(n_24289), .o(n_24462) );
oa12f80 g736401 ( .a(n_320), .b(n_43730), .c(FE_OFN3_n_43918), .o(n_43773) );
ao12f80 g746301 ( .a(n_34917), .b(n_34916), .c(n_34915), .o(n_35678) );
in01f80 newInst_2565 ( .a(newNet_1406), .o(newNet_2565) );
oa12f80 g745722 ( .a(n_33966), .b(n_34069), .c(n_34013), .o(n_34121) );
in01f80 g757092 ( .a(n_23264), .o(n_23265) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_19_ ( .ck(newNet_2860), .d(n_11453), .o(delay_add_ln22_unr8_stage4_stallmux_q_19_) );
no02f80 g743256 ( .a(n_37992), .b(n_37189), .o(n_38044) );
in01f80 g752129 ( .a(n_28071), .o(n_28042) );
no02f80 FE_RC_1892_0 ( .a(n_11879), .b(n_12121), .o(FE_RN_590_0) );
in01f80 g767991 ( .a(n_12688), .o(n_12689) );
na02f80 g777790 ( .a(n_3202), .b(n_3131), .o(n_3254) );
na02f80 g772727 ( .a(n_8180), .b(n_8197), .o(n_8181) );
oa22f80 g741559 ( .a(n_38690), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .c(n_38647), .d(n_38778), .o(n_38696) );
na02f80 g758127 ( .a(n_22298), .b(n_22149), .o(n_22299) );
in01f80 newInst_2273 ( .a(newNet_2084), .o(newNet_2273) );
na02f80 g775747 ( .a(n_5300), .b(n_4078), .o(n_5301) );
in01f80 g772007 ( .a(n_9281), .o(n_9282) );
in01f80 g742493 ( .a(n_37687), .o(n_37688) );
in01f80 g778734 ( .a(n_2612), .o(n_2613) );
no02f80 g760396 ( .a(n_20097), .b(n_20092), .o(n_20169) );
na02f80 g768969 ( .a(n_12085), .b(n_12084), .o(n_12086) );
na02f80 FE_RC_4085_0 ( .a(FE_RN_1785_0), .b(FE_OCP_RBN3728_FE_RN_1787_0), .o(FE_RN_1786_0) );
in01f80 FE_OCPC1533_n_29842 ( .a(n_29842), .o(FE_OCPN1533_n_29842) );
na02f80 g765251 ( .a(n_15025), .b(n_15058), .o(n_15204) );
oa22f80 FE_RC_1658_0 ( .a(FE_OCP_RBN2353_n_13858), .b(n_14034), .c(FE_OCP_RBN1173_n_13858), .d(n_14071), .o(n_14197) );
ao12f80 g737952 ( .a(n_42201), .b(n_42272), .c(n_42271), .o(n_42370) );
no02f80 g762089 ( .a(FE_OCP_RBN2205_n_18242), .b(n_17805), .o(n_18593) );
in01f80 newInst_1838 ( .a(newNet_1837), .o(newNet_1838) );
ao22s80 FE_RC_1295_0 ( .a(n_2913), .b(n_3645), .c(n_3029), .d(FE_OCP_RBN2536_n_3645), .o(n_3521) );
in01f80 g743765 ( .a(n_37294), .o(n_37295) );
in01f80 newInst_3199 ( .a(newNet_3198), .o(newNet_3199) );
oa12f80 g756180 ( .a(n_24817), .b(n_24816), .c(n_24815), .o(n_25285) );
no02f80 g748753 ( .a(n_31059), .b(n_30966), .o(n_31113) );
na02f80 g776772 ( .a(n_3955), .b(n_3954), .o(n_3956) );
no02f80 g758047 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_), .o(n_23053) );
no02f80 g773025 ( .a(n_8037), .b(n_8081), .o(n_8172) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_4_ ( .ck(newNet_2814), .d(n_10088), .o(delay_add_ln22_unr8_stage4_stallmux_q_4_) );
no02f80 g763081 ( .a(n_17414), .b(n_17234), .o(n_17415) );
in01f80 g751914 ( .a(n_29309), .o(n_29310) );
in01f80 g755256 ( .a(n_25114), .o(n_25115) );
oa12f80 g737849 ( .a(n_42362), .b(n_42547), .c(n_42309), .o(n_42622) );
in01f80 newInst_3397 ( .a(newNet_3396), .o(newNet_3397) );
oa22f80 g737652 ( .a(FE_OCPN887_n_42367), .b(n_42093), .c(n_42392), .d(n_42072), .o(n_42758) );
in01f80 FE_RC_3578_0 ( .a(n_14466), .o(FE_RN_1557_0) );
no02f80 g764820 ( .a(n_15688), .b(n_15727), .o(n_15728) );
na02f80 g749932 ( .a(n_30016), .b(n_29985), .o(n_30017) );
oa22f80 FE_RC_2917_0 ( .a(n_10089), .b(n_10315), .c(n_10090), .d(n_10314), .o(n_10477) );
in01f80 g740384 ( .a(n_39851), .o(n_40193) );
no02f80 g750163 ( .a(n_29738), .b(n_29740), .o(n_29816) );
na02f80 g777633 ( .a(n_3598), .b(FE_OCPN848_n_3597), .o(n_3701) );
in01f80 newInst_3002 ( .a(newNet_2194), .o(newNet_3002) );
na02f80 g779306 ( .a(n_1671), .b(n_1652), .o(n_1789) );
ao12f80 g775103 ( .a(n_5926), .b(n_5955), .c(n_5815), .o(n_6021) );
no02f80 g764128 ( .a(n_16563), .b(n_16475), .o(n_16585) );
oa12f80 g758002 ( .a(n_22725), .b(n_22734), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n_22736) );
in01f80 g754727 ( .a(n_26601), .o(n_26602) );
in01f80 FE_OCP_RBC2986_n_35539 ( .a(FE_OCP_RBN3697_n_35543), .o(FE_OCP_RBN2986_n_35539) );
no02f80 g740825 ( .a(n_39401), .b(n_39075), .o(n_39439) );
ao12f80 g770289 ( .a(n_10604), .b(n_10626), .c(n_10677), .o(n_10722) );
in01f80 g745242 ( .a(n_36025), .o(n_36026) );
na02f80 g751566 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_24_), .o(n_28631) );
in01f80 g764348 ( .a(n_16452), .o(n_16453) );
na02f80 FE_RC_3499_0 ( .a(FE_RN_1509_0), .b(n_31959), .o(n_32000) );
in01f80 FE_RC_4186_0 ( .a(n_24389), .o(FE_RN_1832_0) );
in01f80 FE_OCP_RBC1146_n_13098 ( .a(FE_OCP_RBN1145_n_13098), .o(FE_OCP_RBN1146_n_13098) );
in01f80 g744522 ( .a(n_35440), .o(n_35441) );
na02f80 g772283 ( .a(n_8684), .b(n_8120), .o(n_8733) );
in01f80 g768134 ( .a(n_12629), .o(n_12614) );
in01f80 g759953 ( .a(n_21599), .o(n_21104) );
oa12f80 g774396 ( .a(n_6849), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n_6965) );
na02f80 g751356 ( .a(n_29457), .b(n_29456), .o(n_29458) );
in01f80 FE_OCP_RBC3020_n_39942 ( .a(n_39942), .o(FE_OCP_RBN3020_n_39942) );
no02f80 g755984 ( .a(n_24265), .b(n_23788), .o(n_24309) );
in01f80 newInst_1516 ( .a(newNet_1323), .o(newNet_1516) );
no02f80 g779361 ( .a(n_1588), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .o(n_1644) );
in01f80 g751505 ( .a(n_28674), .o(n_28675) );
in01f80 g741685 ( .a(n_38591), .o(n_38605) );
no02f80 g744075 ( .a(n_44223), .b(n_34903), .o(n_36147) );
na02f80 g737501 ( .a(n_42541), .b(n_42289), .o(n_42554) );
ao12f80 g761218 ( .a(n_20050), .b(n_20011), .c(n_19980), .o(n_21137) );
na02f80 g750416 ( .a(n_29568), .b(FE_OCPN1464_n_29630), .o(n_29615) );
in01f80 g764558 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .o(n_16591) );
in01f80 FE_OCP_RBC3649_n_35169 ( .a(n_35169), .o(FE_OCP_RBN3649_n_35169) );
in01f80 FE_OCP_RBC2188_n_37686 ( .a(FE_OCP_RBN2187_n_37686), .o(FE_OCP_RBN2188_n_37686) );
in01f80 FE_OCP_RBC2132_n_40629 ( .a(n_40629), .o(FE_OCP_RBN2132_n_40629) );
na02f80 g765977 ( .a(n_13577), .b(n_14770), .o(n_14845) );
no02f80 g759221 ( .a(n_21154), .b(n_21181), .o(n_21271) );
in01f80 g775413 ( .a(n_5558), .o(n_5601) );
in01f80 g748685 ( .a(n_31208), .o(n_31300) );
no02f80 g767440 ( .a(n_13331), .b(n_13330), .o(n_13358) );
na02f80 g758090 ( .a(n_44268), .b(FE_OCP_RBN3854_n_20848), .o(n_22263) );
in01f80 FE_RC_1675_0 ( .a(FE_RN_467_0), .o(n_28368) );
na02f80 g773821 ( .a(FE_RN_955_0), .b(n_7165), .o(n_7469) );
no02f80 g776570 ( .a(n_4283), .b(FE_OCP_RBN2692_FE_OCPN843_n_3912), .o(n_4350) );
no02f80 g740968 ( .a(n_39235), .b(FE_OCP_RBN3626_n_38870), .o(n_39282) );
no02f80 FE_RC_2225_0 ( .a(FE_RN_804_0), .b(FE_RN_807_0), .o(n_33331) );
oa22f80 g779978 ( .a(n_1268), .b(n_999), .c(n_1267), .d(n_1000), .o(n_1274) );
no02f80 g775985 ( .a(n_5253), .b(n_47019), .o(n_5288) );
na02f80 g766928 ( .a(n_14041), .b(n_14040), .o(n_14076) );
no02f80 g755722 ( .a(n_24346), .b(n_24014), .o(n_24375) );
na02f80 g760949 ( .a(n_19356), .b(n_19348), .o(n_19514) );
oa12f80 g756444 ( .a(n_23599), .b(n_23738), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n_23856) );
oa12f80 g749535 ( .a(n_30495), .b(n_30494), .c(n_30493), .o(n_31871) );
in01f80 FE_OCP_RBC3472_n_7886 ( .a(FE_OCP_RBN3470_n_7886), .o(FE_OCP_RBN3472_n_7886) );
oa12f80 g784676 ( .a(n_4664), .b(n_4661), .c(n_4267), .o(n_47006) );
na02f80 g768423 ( .a(n_12453), .b(n_12452), .o(n_12507) );
oa12f80 g761230 ( .a(n_19072), .b(n_19186), .c(n_19130), .o(n_19200) );
na02f80 g738408 ( .a(n_41411), .b(n_41414), .o(n_41798) );
oa12f80 g761363 ( .a(n_19981), .b(n_20086), .c(n_19927), .o(n_20700) );
no02f80 g761053 ( .a(n_19180), .b(n_19209), .o(n_19355) );
in01f80 FE_OCP_RBC2836_FE_RN_745_0 ( .a(FE_RN_745_0), .o(FE_OCP_RBN2836_FE_RN_745_0) );
ao12f80 g737279 ( .a(n_42591), .b(n_42889), .c(n_42592), .o(n_42902) );
na02f80 g755459 ( .a(n_24800), .b(n_24644), .o(n_24870) );
na02f80 g767605 ( .a(n_13422), .b(n_13421), .o(n_13423) );
na02f80 g759569 ( .a(n_20794), .b(n_20795), .o(n_20878) );
no02f80 FE_RC_2424_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .b(FE_RN_960_0), .o(FE_RN_961_0) );
no02f80 g763910 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_), .o(n_17359) );
in01f80 FE_OCPC1751_n_29420 ( .a(n_29420), .o(FE_OCPN1751_n_29420) );
na02f80 g744985 ( .a(FE_OCP_RBN2640_n_34921), .b(n_30504), .o(n_34974) );
in01f80 FE_OCPC1435_n_19855 ( .a(n_19855), .o(FE_OCPN1435_n_19855) );
na02f80 g747189 ( .a(n_33931), .b(n_33930), .o(n_33932) );
no02f80 g778067 ( .a(n_3040), .b(n_3039), .o(n_3061) );
no02f80 g738941 ( .a(n_41154), .b(n_40862), .o(n_41197) );
na02f80 g769623 ( .a(n_11326), .b(n_11346), .o(n_11411) );
ao22s80 FE_RC_51_0 ( .a(n_5998), .b(n_6021), .c(n_5997), .d(n_6022), .o(n_6135) );
no02f80 g773230 ( .a(n_7572), .b(n_7571), .o(n_7573) );
in01f80 FE_OCPC3762_n_34222 ( .a(n_34222), .o(FE_OCPN3762_n_34222) );
no02f80 g751193 ( .a(n_29818), .b(n_29907), .o(n_30304) );
in01f80 g763174 ( .a(n_17475), .o(n_17550) );
na02f80 g762353 ( .a(n_18421), .b(n_18419), .o(n_18449) );
na02f80 g763067 ( .a(n_17588), .b(n_17553), .o(n_17554) );
in01f80 g782633 ( .a(n_44060), .o(n_509) );
ao12f80 g777382 ( .a(n_3218), .b(n_3416), .c(n_3179), .o(n_3417) );
in01f80 newInst_1812 ( .a(newNet_1219), .o(newNet_1812) );
na02f80 g753810 ( .a(n_26330), .b(n_26246), .o(n_26410) );
in01f80 FE_OCP_RBC2526_n_3421 ( .a(n_3421), .o(FE_OCP_RBN2526_n_3421) );
in01f80 g738768 ( .a(n_41355), .o(n_41367) );
na02f80 g766144 ( .a(n_14576), .b(n_14549), .o(n_14689) );
na02f80 g760243 ( .a(FE_OCP_RBN3617_n_20249), .b(n_20523), .o(n_20628) );
no02f80 g741807 ( .a(n_38394), .b(n_38393), .o(n_38395) );
in01f80 newInst_2014 ( .a(newNet_503), .o(newNet_2014) );
ao12f80 g769290 ( .a(n_11337), .b(n_11410), .c(n_11392), .o(n_11434) );
in01f80 g750312 ( .a(n_29788), .o(n_29763) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_12_ ( .ck(newNet_1875), .d(n_16592), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_12_) );
in01f80 g768582 ( .a(n_12268), .o(n_12269) );
oa22f80 g751088 ( .a(n_30303), .b(n_29535), .c(n_30156), .d(n_29999), .o(n_30589) );
na02f80 g778024 ( .a(n_3000), .b(n_2231), .o(n_3001) );
in01f80 g753380 ( .a(n_27098), .o(n_27110) );
in01f80 newInst_1394 ( .a(newNet_1393), .o(newNet_1394) );
oa22f80 FE_RC_1229_0 ( .a(n_17378), .b(n_17627), .c(n_17379), .d(n_17601), .o(n_17759) );
na02f80 g751311 ( .a(n_29598), .b(n_29332), .o(n_29654) );
no02f80 g744693 ( .a(FE_OCP_RBN2808_n_35285), .b(n_35265), .o(n_35323) );
na02f80 g745736 ( .a(n_34219), .b(n_34184), .o(n_34220) );
in01f80 g762722 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_25_), .o(n_18331) );
in01f80 g748580 ( .a(n_31424), .o(n_31425) );
in01f80 g755356 ( .a(n_24983), .o(n_24984) );
in01f80 newInst_2083 ( .a(newNet_1933), .o(newNet_2083) );
in01f80 g743570 ( .a(n_36549), .o(n_36534) );
in01f80 g747828 ( .a(n_33390), .o(n_33440) );
na02f80 g763169 ( .a(n_17402), .b(n_17284), .o(n_17403) );
ao22s80 g736478 ( .a(n_43715), .b(n_43588), .c(n_43714), .d(n_43587), .o(n_43749) );
no02f80 g772396 ( .a(n_8529), .b(n_8544), .o(n_8619) );
in01f80 g739111 ( .a(n_41072), .o(n_41108) );
oa22f80 g745568 ( .a(FE_OCPN1732_n_34369), .b(n_33545), .c(n_34286), .d(n_34347), .o(n_34847) );
no02f80 g740391 ( .a(FE_OCP_RBN3021_n_39942), .b(n_39488), .o(n_39934) );
in01f80 g747819 ( .a(n_33311), .o(n_33312) );
na02f80 g769652 ( .a(n_11301), .b(FE_OCPN3785_FE_OCP_RBN2831_n_10198), .o(n_11325) );
no02f80 g738481 ( .a(n_41393), .b(n_41392), .o(n_41410) );
in01f80 g777226 ( .a(n_3751), .o(n_3752) );
na02f80 g775771 ( .a(n_6131), .b(n_4182), .o(n_5089) );
in01f80 g775125 ( .a(n_5947), .o(n_5948) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_8_ ( .ck(newNet_3470), .d(n_21732), .o(delay_add_ln22_unr14_stage6_stallmux_q_8_) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_10_ ( .ck(newNet_893), .d(n_32353), .o(delay_xor_ln21_unr21_stage8_stallmux_q_10_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_30_ ( .ck(newNet_1582), .d(n_27676), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_) );
in01f80 newInst_3159 ( .a(newNet_262), .o(newNet_3159) );
in01f80 g761864 ( .a(n_18407), .o(n_18408) );
na02f80 g774967 ( .a(n_6102), .b(n_6065), .o(n_6103) );
na02f80 g758868 ( .a(n_21441), .b(n_21395), .o(n_21586) );
na02f80 g773639 ( .a(n_7358), .b(n_7124), .o(n_7381) );
no02f80 g761552 ( .a(n_18861), .b(FE_OCPN1456_n_18860), .o(n_18862) );
no02f80 g754576 ( .a(n_25432), .b(n_25431), .o(n_25433) );
in01f80 newInst_2473 ( .a(newNet_56), .o(newNet_2473) );
ao12f80 g762422 ( .a(n_17977), .b(FE_OCP_RBN2147_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_15_), .o(n_18023) );
in01f80 g774945 ( .a(n_6181), .o(n_6182) );
in01f80 FE_OCPC1229_n_46101 ( .a(FE_OCPN1228_n_46101), .o(FE_OCPN1229_n_46101) );
no02f80 g777107 ( .a(n_3666), .b(n_3698), .o(n_3846) );
no02f80 FE_RC_215_0 ( .a(FE_RN_69_0), .b(FE_RN_70_0), .o(FE_RN_71_0) );
in01f80 g767772 ( .a(n_13083), .o(n_13213) );
na02f80 g746719 ( .a(n_33022), .b(n_32978), .o(n_33083) );
in01f80 newInst_1315 ( .a(newNet_1011), .o(newNet_1315) );
in01f80 g736847 ( .a(n_43549), .o(n_43550) );
na02f80 g751838 ( .a(n_29150), .b(n_29070), .o(n_29151) );
na02f80 g753331 ( .a(n_27100), .b(n_27099), .o(n_27243) );
oa12f80 g774847 ( .a(n_6012), .b(n_6080), .c(n_6178), .o(n_6238) );
in01f80 g750494 ( .a(n_31256), .o(n_31211) );
in01f80 g768685 ( .a(n_12186), .o(n_12187) );
in01f80 g777795 ( .a(n_3405), .o(n_3373) );
na02f80 g776912 ( .a(n_3776), .b(n_3862), .o(n_3855) );
no02f80 g767964 ( .a(n_12737), .b(n_12982), .o(n_13354) );
in01f80 newInst_297 ( .a(newNet_296), .o(newNet_297) );
in01f80 g763268 ( .a(n_17274), .o(n_17449) );
na02f80 g748116 ( .a(n_32824), .b(n_32823), .o(n_32825) );
in01f80 g750044 ( .a(n_29897), .o(n_29965) );
na02f80 g762254 ( .a(n_18729), .b(n_18728), .o(n_18730) );
in01f80 fopt783570 ( .a(n_38660), .o(n_45192) );
na02f80 g741965 ( .a(n_37975), .b(n_37986), .o(n_38040) );
in01f80 g766578 ( .a(n_13927), .o(n_13932) );
in01f80 g760673 ( .a(n_19747), .o(n_19814) );
oa12f80 g752624 ( .a(n_27301), .b(n_27476), .c(n_27219), .o(n_27569) );
na02f80 g749256 ( .a(n_30744), .b(n_30743), .o(n_30766) );
in01f80 g775475 ( .a(n_5724), .o(n_5708) );
na02f80 g745536 ( .a(n_34509), .b(n_34537), .o(n_34562) );
in01f80 FE_RC_4053_0 ( .a(FE_RN_1763_0), .o(n_16563) );
na02f80 g780132 ( .a(n_1181), .b(n_1180), .o(n_1182) );
na02f80 g755577 ( .a(FE_OCP_RBN2420_n_24505), .b(n_22393), .o(n_24573) );
in01f80 FE_OCPC1773_n_30210 ( .a(n_30210), .o(FE_OCPN1773_n_30210) );
in01f80 FE_RC_2084_0 ( .a(FE_RN_714_0), .o(n_30843) );
in01f80 g737165 ( .a(n_43103), .o(n_43097) );
no02f80 g778254 ( .a(n_2704), .b(n_2650), .o(n_2871) );
na02f80 g765189 ( .a(n_15198), .b(n_14210), .o(n_15311) );
oa12f80 g758696 ( .a(n_21501), .b(FE_OCP_RBN1705_n_21658), .c(n_21711), .o(n_21745) );
na02f80 g775585 ( .a(n_5728), .b(n_5727), .o(n_5729) );
no02f80 g741290 ( .a(n_44955), .b(n_38908), .o(n_38940) );
in01f80 newInst_2498 ( .a(newNet_2497), .o(newNet_2498) );
no02f80 g779578 ( .a(n_1374), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1399) );
ao12f80 g741800 ( .a(n_38392), .b(n_38391), .c(n_38390), .o(n_38493) );
in01f80 g765938 ( .a(n_14815), .o(n_14816) );
na02f80 g758064 ( .a(n_22646), .b(n_22699), .o(n_23319) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_1_ ( .ck(newNet_1998), .d(n_9878), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_) );
oa22f80 g765407 ( .a(n_15874), .b(n_16246), .c(n_16245), .d(n_14433), .o(n_16349) );
oa22f80 FE_RC_2976_0 ( .a(n_10692), .b(n_10722), .c(n_10693), .d(FE_OCP_RBN2947_n_10722), .o(n_10828) );
na02f80 g771346 ( .a(n_9344), .b(n_9294), .o(n_9535) );
na02f80 g741815 ( .a(n_38441), .b(n_38440), .o(n_38442) );
na02f80 g769749 ( .a(n_11197), .b(n_11174), .o(n_11297) );
ao12f80 g754596 ( .a(n_26385), .b(FE_OCP_RBN2960_n_26231), .c(n_26310), .o(n_26951) );
oa12f80 g780115 ( .a(n_1182), .b(n_1181), .c(n_1180), .o(n_1206) );
no02f80 g775616 ( .a(n_4556), .b(FE_OCP_RBN2932_n_5307), .o(n_5388) );
in01f80 newInst_1999 ( .a(newNet_1553), .o(newNet_1999) );
in01f80 newInst_1269 ( .a(newNet_1268), .o(newNet_1269) );
na02f80 g755050 ( .a(n_25413), .b(n_25412), .o(n_25414) );
in01f80 FE_RC_1361_0 ( .a(n_5310), .o(FE_RN_405_0) );
in01f80 newInst_3466 ( .a(newNet_375), .o(newNet_3466) );
ao12f80 g781274 ( .a(n_93), .b(n_46055), .c(beta_22), .o(n_254) );
na02f80 g739728 ( .a(n_40538), .b(n_40170), .o(n_40542) );
no02f80 g746924 ( .a(n_32860), .b(n_32464), .o(n_32963) );
oa12f80 g776122 ( .a(n_4892), .b(n_4891), .c(n_4890), .o(n_4997) );
na02f80 g745167 ( .a(n_36230), .b(n_36229), .o(n_36231) );
in01f80 g775540 ( .a(n_5486), .o(n_5419) );
in01f80 g767453 ( .a(n_13301), .o(n_13329) );
ao12f80 g780848 ( .a(n_452), .b(n_521), .c(n_447), .o(n_611) );
in01f80 newInst_1607 ( .a(newNet_1466), .o(newNet_1607) );
no02f80 g778540 ( .a(n_2299), .b(n_2766), .o(n_2310) );
na02f80 FE_RC_360_0 ( .a(FE_RN_105_0), .b(FE_RN_106_0), .o(FE_RN_107_0) );
in01f80 newInst_2806 ( .a(newNet_2805), .o(newNet_2806) );
oa12f80 g761250 ( .a(n_19765), .b(n_19764), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21052) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_15_ ( .ck(newNet_2016), .d(n_11278), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_) );
in01f80 g754148 ( .a(n_26057), .o(n_26058) );
in01f80 g749924 ( .a(n_30320), .o(n_30321) );
in01f80 g751792 ( .a(n_28316), .o(n_28317) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_1_ ( .ck(newNet_863), .d(n_40599), .o(delay_xor_ln21_unr28_stage10_stallmux_q_1_) );
na02f80 g758075 ( .a(n_22150), .b(n_20688), .o(n_22200) );
na02f80 g763120 ( .a(n_17146), .b(n_16880), .o(n_17200) );
oa22f80 FE_RC_3147_0 ( .a(n_14881), .b(n_14901), .c(n_14882), .d(n_14902), .o(n_15001) );
no02f80 g777243 ( .a(n_3508), .b(n_3514), .o(n_5447) );
no02f80 g778656 ( .a(n_2387), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .o(n_2437) );
na02f80 g776316 ( .a(n_4429), .b(FE_OCP_RBN2731_n_4219), .o(n_4507) );
in01f80 g748712 ( .a(n_31244), .o(n_31245) );
oa12f80 g766096 ( .a(n_14379), .b(n_14484), .c(n_14479), .o(n_14485) );
no02f80 g769727 ( .a(n_11293), .b(n_11292), .o(n_11394) );
in01f80 g766159 ( .a(n_14550), .o(n_14551) );
ao12f80 g760671 ( .a(n_19594), .b(n_19656), .c(n_19719), .o(n_19809) );
na02f80 g771302 ( .a(n_9152), .b(n_9355), .o(n_9356) );
oa12f80 g750486 ( .a(n_29444), .b(n_29542), .c(n_29498), .o(n_29606) );
oa22f80 FE_RC_58_0 ( .a(n_18262), .b(n_18412), .c(n_18261), .d(n_18438), .o(n_18600) );
in01f80 newInst_2361 ( .a(newNet_2360), .o(newNet_2361) );
in01f80 newInst_2073 ( .a(newNet_2072), .o(newNet_2073) );
in01f80 FE_OCP_RBC1339_n_32653 ( .a(n_32653), .o(FE_OCP_RBN1339_n_32653) );
no02f80 g745018 ( .a(n_34927), .b(n_34747), .o(n_34971) );
no02f80 g762098 ( .a(n_18265), .b(n_18264), .o(n_18276) );
oa22f80 g780260 ( .a(n_45816), .b(n_1122), .c(n_863), .d(n_1208), .o(n_1010) );
oa12f80 g761102 ( .a(n_19144), .b(n_19143), .c(n_19142), .o(n_21058) );
na02f80 g746166 ( .a(n_33715), .b(n_33714), .o(n_33777) );
no02f80 g741015 ( .a(n_39008), .b(n_38986), .o(n_39141) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_14_ ( .ck(newNet_2488), .d(n_32234), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_) );
na02f80 g736573 ( .a(n_43682), .b(n_43563), .o(n_43681) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_3_ ( .ck(newNet_378), .d(n_40587), .o(delay_xor_ln22_unr28_stage10_stallmux_q_3_) );
in01f80 newInst_1071 ( .a(newNet_1070), .o(newNet_1071) );
in01f80 g774078 ( .a(n_6775), .o(n_6776) );
in01f80 g764275 ( .a(n_47340), .o(n_16484) );
na02f80 g750325 ( .a(n_29664), .b(n_29631), .o(n_29718) );
in01f80 newInst_636 ( .a(newNet_635), .o(newNet_636) );
no02f80 g774329 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .o(n_6880) );
in01f80 g774584 ( .a(n_6563), .o(n_6556) );
in01f80 g742114 ( .a(n_38160), .o(n_38161) );
in01f80 g747398 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .o(n_32401) );
ao12f80 g777756 ( .a(n_3043), .b(n_3293), .c(n_3329), .o(n_3340) );
na02f80 g757547 ( .a(n_23320), .b(n_23319), .o(n_23321) );
in01f80 FE_RC_1945_0 ( .a(FE_RN_622_0), .o(n_13957) );
in01f80 FE_OCPC1735_n_37877 ( .a(n_37877), .o(FE_OCPN1735_n_37877) );
no02f80 g778535 ( .a(n_2762), .b(n_2838), .o(n_2839) );
no02f80 g759117 ( .a(n_21461), .b(n_45080), .o(n_21490) );
oa12f80 g775753 ( .a(n_4917), .b(n_4907), .c(n_4825), .o(n_5031) );
no02f80 g756387 ( .a(n_24330), .b(n_23958), .o(n_24380) );
na02f80 g784773 ( .a(n_9410), .b(FE_OCPN997_n_44460), .o(n_47259) );
in01f80 g776790 ( .a(n_4331), .o(n_4332) );
in01f80 g739327 ( .a(n_40738), .o(n_40698) );
na02f80 g776228 ( .a(n_4814), .b(n_4447), .o(n_4845) );
na02f80 g775135 ( .a(n_5788), .b(n_5801), .o(n_5910) );
na02f80 g750847 ( .a(n_29039), .b(n_29036), .o(n_29037) );
na02f80 FE_RC_1734_0 ( .a(n_36886), .b(FE_RN_482_0), .o(n_36921) );
no02f80 g750516 ( .a(n_29473), .b(n_29430), .o(n_29503) );
in01f80 newInst_3294 ( .a(newNet_2089), .o(newNet_3294) );
na02f80 g742921 ( .a(n_36956), .b(n_37068), .o(n_37116) );
oa12f80 g776659 ( .a(n_3997), .b(n_4297), .c(n_4108), .o(n_4432) );
na02f80 g758742 ( .a(n_22246), .b(n_21723), .o(n_22363) );
ao12f80 g738101 ( .a(n_42055), .b(n_42070), .c(n_42054), .o(n_42102) );
in01f80 g747211 ( .a(n_32697), .o(n_32736) );
ao12f80 g773042 ( .a(FE_OCP_RBN3453_FE_OCPN1240_n_7721), .b(n_7824), .c(n_7908), .o(n_7965) );
na02f80 g766591 ( .a(n_13924), .b(n_13277), .o(n_13925) );
no02f80 g743432 ( .a(n_36588), .b(n_36750), .o(n_36614) );
no02f80 g766488 ( .a(n_13998), .b(n_13262), .o(n_14093) );
no02f80 g779767 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_), .o(n_1603) );
no02f80 g739296 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_41038) );
no02f80 g776372 ( .a(n_4689), .b(n_4765), .o(n_5058) );
no02f80 g765337 ( .a(FE_OCP_RBN2707_n_15135), .b(n_15518), .o(n_15519) );
na02f80 g775500 ( .a(n_5456), .b(FE_OCP_RBN2734_n_4219), .o(n_5524) );
na02f80 g776215 ( .a(n_4667), .b(n_4017), .o(n_4740) );
na02f80 g736821 ( .a(n_43133), .b(n_43129), .o(n_43142) );
no02f80 g767677 ( .a(n_13356), .b(n_13377), .o(n_13375) );
in01f80 newInst_2577 ( .a(newNet_1637), .o(newNet_2577) );
in01f80 g771002 ( .a(n_9891), .o(n_9985) );
na02f80 g773820 ( .a(n_7153), .b(n_6925), .o(n_7188) );
no02f80 g763107 ( .a(n_17507), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_4_), .o(n_17548) );
in01f80 g753155 ( .a(n_27523), .o(n_27524) );
na03f80 g751850 ( .a(n_28991), .b(n_28926), .c(n_28925), .o(n_28992) );
in01f80 newInst_3458 ( .a(newNet_3457), .o(newNet_3458) );
no02f80 g755488 ( .a(n_24623), .b(FE_OCPN1474_n_24624), .o(n_24704) );
no02f80 g740022 ( .a(n_40010), .b(FE_OCP_RBN3715_n_39913), .o(n_40120) );
na02f80 g774817 ( .a(n_6228), .b(n_5640), .o(n_6395) );
na02f80 g754505 ( .a(n_26933), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_26934) );
no02f80 g743520 ( .a(n_36559), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36580) );
in01f80 g748125 ( .a(n_31968), .o(n_31969) );
ao12f80 g768892 ( .a(n_11888), .b(FE_OCP_RBN2124_n_45224), .c(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .o(n_11945) );
na02f80 g762432 ( .a(n_18021), .b(n_17873), .o(n_18090) );
in01f80 FE_OCP_RBC2007_n_45209 ( .a(n_45209), .o(FE_OCP_RBN2007_n_45209) );
in01f80 g768404 ( .a(n_12459), .o(n_12460) );
no02f80 g746272 ( .a(n_33583), .b(n_33541), .o(n_33617) );
in01f80 g753440 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n_27575) );
no02f80 g766973 ( .a(n_13668), .b(n_13682), .o(n_15609) );
no02f80 g740354 ( .a(n_39729), .b(n_39687), .o(n_39742) );
ao12f80 g766761 ( .a(n_13214), .b(n_13711), .c(n_13174), .o(n_13732) );
in01f80 g741560 ( .a(n_38712), .o(n_39679) );
in01f80 newInst_1014 ( .a(newNet_267), .o(newNet_1014) );
in01f80 g752939 ( .a(n_27878), .o(n_27879) );
ao12f80 g764765 ( .a(n_15461), .b(n_45137), .c(n_15410), .o(n_15704) );
in01f80 newInst_1468 ( .a(newNet_494), .o(newNet_1468) );
no02f80 g768796 ( .a(n_12062), .b(n_12061), .o(n_12092) );
in01f80 g742747 ( .a(n_37348), .o(n_37349) );
na02f80 g768246 ( .a(n_12571), .b(n_12570), .o(n_12572) );
in01f80 g777330 ( .a(n_4426), .o(n_4503) );
in01f80 g737204 ( .a(n_42983), .o(n_42984) );
na02f80 g773630 ( .a(n_7370), .b(n_7359), .o(n_7425) );
in01f80 g756551 ( .a(n_23853), .o(n_23820) );
no02f80 g746384 ( .a(n_33518), .b(n_33201), .o(n_33558) );
oa12f80 g758636 ( .a(n_21670), .b(n_22396), .c(n_21600), .o(n_22487) );
in01f80 g752609 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_16_), .o(n_27710) );
na02f80 g776963 ( .a(n_3985), .b(n_3984), .o(n_3986) );
no02f80 g778465 ( .a(n_2629), .b(n_2126), .o(n_2684) );
in01f80 g773619 ( .a(n_7349), .o(n_7350) );
no02f80 g780386 ( .a(n_1079), .b(n_919), .o(n_874) );
ao22s80 g736550 ( .a(n_43567), .b(n_43592), .c(n_43568), .d(n_43591), .o(n_43662) );
in01f80 newInst_907 ( .a(newNet_906), .o(newNet_907) );
na02f80 g773632 ( .a(n_7358), .b(n_7178), .o(n_7359) );
oa22f80 FE_RC_1257_0 ( .a(n_34533), .b(n_34900), .c(n_34534), .d(n_34874), .o(n_35001) );
ao22s80 g736397 ( .a(n_43783), .b(n_43425), .c(n_43792), .d(n_43426), .o(n_43847) );
no02f80 g741311 ( .a(n_38830), .b(n_38829), .o(n_38993) );
na02f80 g742404 ( .a(n_37722), .b(n_37708), .o(n_37838) );
no02f80 g750725 ( .a(n_29193), .b(n_28767), .o(n_29220) );
na02f80 g772920 ( .a(n_7902), .b(n_7870), .o(n_7871) );
na02f80 g757034 ( .a(n_23743), .b(n_23903), .o(n_23986) );
in01f80 g758419 ( .a(FE_OCPN1514_FE_OFN738_n_22641), .o(n_23398) );
in01f80 g747805 ( .a(n_33740), .o(n_33741) );
na02f80 g739441 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_22_), .o(n_40882) );
in01f80 newInst_863 ( .a(newNet_862), .o(newNet_863) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_17_ ( .ck(newNet_1860), .d(n_16815), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_) );
in01f80 g758847 ( .a(n_21506), .o(n_21550) );
no02f80 g778595 ( .a(n_2366), .b(n_44344), .o(n_2477) );
na02f80 g749976 ( .a(n_30245), .b(n_30215), .o(n_30275) );
no02f80 g763810 ( .a(n_17104), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .o(n_17105) );
ao22s80 g738886 ( .a(n_41163), .b(n_41079), .c(n_41164), .d(n_41080), .o(n_41263) );
in01f80 fopt783509 ( .a(FE_OCP_RBN3410_n_45120), .o(n_45002) );
in01f80 newInst_802 ( .a(newNet_801), .o(newNet_802) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_18_ ( .ck(newNet_833), .d(n_1333), .o(delay_xor_ln21_unr3_stage2_stallmux_q_18_) );
in01f80 FE_OCPC3184_n_22294 ( .a(FE_OCPN3183_n_22294), .o(FE_OCPN3184_n_22294) );
in01f80 g755602 ( .a(n_24719), .o(n_24681) );
in01f80 newInst_356 ( .a(newNet_355), .o(newNet_356) );
no02f80 g760432 ( .a(n_20070), .b(n_18793), .o(n_20125) );
in01f80 g767905 ( .a(n_12743), .o(n_12744) );
in01f80 g750749 ( .a(n_29233), .o(n_29265) );
oa22f80 g784428 ( .a(n_36637), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46204), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .o(n_46240) );
no02f80 g737533 ( .a(n_42510), .b(n_42447), .o(n_42550) );
no02f80 g749195 ( .a(n_30737), .b(FE_OCPN1490_n_30823), .o(n_30809) );
in01f80 newInst_1756 ( .a(newNet_1038), .o(newNet_1756) );
na02f80 g739472 ( .a(n_40715), .b(n_40714), .o(n_40848) );
in01f80 FE_RC_2521_0 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_), .o(FE_RN_1026_0) );
ao22s80 g768949 ( .a(n_11775), .b(n_11680), .c(n_11665), .d(n_11681), .o(n_12692) );
oa22f80 g765957 ( .a(FE_OCP_RBN3618_n_14841), .b(n_14738), .c(n_14841), .d(n_14706), .o(n_15032) );
in01f80 g737423 ( .a(n_46942), .o(n_42774) );
na02f80 g739318 ( .a(n_45153), .b(n_40590), .o(n_40890) );
na02f80 g758923 ( .a(n_21240), .b(n_21288), .o(n_21330) );
in01f80 g763710 ( .a(n_16810), .o(n_16781) );
na02f80 g746340 ( .a(n_33558), .b(n_33198), .o(n_33635) );
no02f80 g763469 ( .a(FE_OCP_RBN3210_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_3_), .o(n_17084) );
no02f80 g771782 ( .a(n_9099), .b(n_9051), .o(n_9177) );
oa22f80 FE_RC_3289_0 ( .a(n_30766), .b(n_30864), .c(n_30767), .d(n_30863), .o(n_31013) );
in01f80 g773539 ( .a(n_7480), .o(n_7493) );
in01f80 g772599 ( .a(n_8482), .o(n_8483) );
no02f80 g765191 ( .a(n_16020), .b(n_16016), .o(n_16065) );
in01f80 g768234 ( .a(n_12677), .o(n_12721) );
in01f80 FE_OCP_RBC3710_n_46337 ( .a(FE_OCP_RBN3039_n_46337), .o(FE_OCP_RBN3710_n_46337) );
na02f80 g774528 ( .a(n_6397), .b(n_45474), .o(n_6463) );
in01f80 g759061 ( .a(n_21322), .o(n_21323) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_5_ ( .ck(newNet_3370), .d(n_26731), .o(delay_add_ln22_unr17_stage7_stallmux_q_5_) );
oa12f80 g736494 ( .a(n_43519), .b(n_43665), .c(n_43108), .o(n_43689) );
na02f80 g737732 ( .a(n_42285), .b(n_42073), .o(n_42503) );
oa22f80 g777841 ( .a(n_2913), .b(n_4022), .c(n_3301), .d(n_2759), .o(n_3347) );
in01f80 FE_RC_3243_0 ( .a(FE_RN_1434_0), .o(FE_OFN756_n_44461) );
na02f80 FE_RC_4101_0 ( .a(FE_RN_1794_0), .b(n_31685), .o(FE_RN_1795_0) );
in01f80 newInst_2765 ( .a(newNet_1310), .o(newNet_2765) );
na02f80 g765315 ( .a(n_15021), .b(FE_OCP_RBN2362_n_13785), .o(n_15157) );
na02f80 g766990 ( .a(n_13513), .b(n_12955), .o(n_13519) );
in01f80 g759269 ( .a(n_20949), .o(n_20979) );
ao12f80 g754814 ( .a(n_25281), .b(n_25280), .c(n_25279), .o(n_25363) );
no02f80 g756564 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_23_), .o(n_23823) );
oa22f80 g769741 ( .a(n_11213), .b(n_10248), .c(n_11214), .d(n_10249), .o(n_11286) );
in01f80 newInst_1531 ( .a(newNet_1530), .o(newNet_1531) );
na02f80 g736702 ( .a(n_43274), .b(n_43222), .o(n_43328) );
no02f80 g777690 ( .a(n_3437), .b(FE_OCP_RBN2465_n_4336), .o(n_3462) );
oa12f80 g766856 ( .a(n_13686), .b(n_13685), .c(n_13684), .o(n_13742) );
no02f80 g742443 ( .a(n_37733), .b(n_37716), .o(n_37774) );
no02f80 g768110 ( .a(n_12589), .b(n_12631), .o(n_12632) );
in01f80 g749580 ( .a(n_30527), .o(n_30506) );
no02f80 g761493 ( .a(n_19980), .b(n_19733), .o(n_20069) );
in01f80 g742688 ( .a(n_37377), .o(n_37420) );
in01f80 g767241 ( .a(n_13529), .o(n_13554) );
in01f80 g759683 ( .a(n_20597), .o(n_20598) );
in01f80 newInst_3251 ( .a(newNet_3250), .o(newNet_3251) );
oa12f80 g775939 ( .a(n_5132), .b(n_5144), .c(n_5131), .o(n_5211) );
ao12f80 g741406 ( .a(n_38677), .b(n_38770), .c(n_38708), .o(n_38785) );
na02f80 g780611 ( .a(n_779), .b(n_839), .o(n_868) );
in01f80 g739738 ( .a(n_40540), .o(n_40541) );
na02f80 g764269 ( .a(n_16392), .b(n_16433), .o(n_16485) );
in01f80 newInst_1120 ( .a(newNet_1119), .o(newNet_1120) );
in01f80 g761876 ( .a(n_18546), .o(n_18547) );
in01f80 g742533 ( .a(n_37578), .o(n_37598) );
in01f80 g771692 ( .a(n_9355), .o(n_9328) );
oa12f80 g751400 ( .a(n_29288), .b(n_29287), .c(n_29286), .o(n_29907) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_16_ ( .ck(newNet_3435), .d(n_27580), .o(delay_add_ln22_unr17_stage7_stallmux_q_16_) );
in01f80 g741173 ( .a(n_38951), .o(n_38952) );
oa12f80 g766668 ( .a(n_13707), .b(n_13813), .c(n_13781), .o(n_13814) );
na02f80 g749551 ( .a(n_30355), .b(n_30197), .o(n_30387) );
na02f80 g767782 ( .a(n_12823), .b(n_13086), .o(n_13122) );
in01f80 g769875 ( .a(n_11129), .o(n_11162) );
in01f80 g749843 ( .a(n_31143), .o(n_31144) );
oa12f80 g740323 ( .a(n_39762), .b(n_39761), .c(n_39760), .o(n_39779) );
in01f80 g744280 ( .a(n_35732), .o(n_35821) );
no02f80 g738492 ( .a(FE_OCP_RBN2316_n_41420), .b(n_41628), .o(n_41671) );
no02f80 g741623 ( .a(n_38594), .b(n_38778), .o(n_38648) );
in01f80 g755328 ( .a(n_24969), .o(n_25008) );
in01f80 g745821 ( .a(n_34177), .o(n_34178) );
no02f80 g777299 ( .a(n_4675), .b(n_5168), .o(n_5186) );
in01f80 g761117 ( .a(n_20430), .o(n_19340) );
na02f80 g758725 ( .a(n_21897), .b(n_21896), .o(n_21947) );
in01f80 FE_OCPC1440_n_23339 ( .a(FE_OCPN1439_n_23339), .o(FE_OCPN1440_n_23339) );
oa12f80 g737634 ( .a(n_42446), .b(n_42392), .c(n_42391), .o(n_42764) );
no02f80 g739425 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n_40777) );
ao12f80 g765373 ( .a(n_15876), .b(n_15874), .c(n_15779), .o(n_16572) );
na02f80 g748348 ( .a(n_31682), .b(n_31722), .o(n_31796) );
na02f80 FE_RC_2184_0 ( .a(n_22553), .b(FE_RN_780_0), .o(n_22591) );
na02f80 g746806 ( .a(n_33199), .b(n_33198), .o(n_33215) );
oa22f80 g784347 ( .a(FE_OFN775_n_46137), .b(n_5676), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5748), .o(n_46153) );
na02f80 g755047 ( .a(n_25352), .b(n_25350), .o(n_25382) );
no02f80 g766817 ( .a(n_14342), .b(n_14425), .o(n_14526) );
na02f80 g748969 ( .a(n_30919), .b(n_30744), .o(n_30949) );
no02f80 g746137 ( .a(n_35127), .b(n_35126), .o(n_35128) );
no02f80 g755143 ( .a(n_25050), .b(n_25024), .o(n_25151) );
no02f80 g749447 ( .a(n_30511), .b(n_30790), .o(n_30561) );
in01f80 g756826 ( .a(n_23838), .o(n_23911) );
no02f80 g753135 ( .a(n_27188), .b(n_27391), .o(n_27496) );
ao12f80 g772036 ( .a(n_8822), .b(n_8821), .c(n_8820), .o(n_10079) );
no02f80 g764155 ( .a(n_16561), .b(n_16516), .o(n_16562) );
in01f80 g761098 ( .a(n_19243), .o(n_19244) );
na02f80 g770140 ( .a(n_10902), .b(FE_OCP_RBN2704_n_9411), .o(n_10983) );
ao12f80 g757997 ( .a(n_22849), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n_23618) );
in01f80 FE_OCPC3178_n_21901 ( .a(FE_OCPN3177_n_21901), .o(FE_OCPN3178_n_21901) );
in01f80 g748005 ( .a(n_33029), .o(n_33030) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_2_ ( .ck(newNet_160), .d(n_46382), .o(delay_xor_ln22_unr9_stage4_stallmux_q_2_) );
na02f80 FE_RC_1971_0 ( .a(FE_RN_638_0), .b(n_25321), .o(n_25355) );
na02f80 g762778 ( .a(n_18123), .b(n_17502), .o(n_18157) );
na02f80 g755297 ( .a(n_24967), .b(n_24774), .o(n_24985) );
in01f80 g777459 ( .a(n_3564), .o(n_3604) );
no02f80 g776623 ( .a(n_3982), .b(n_4093), .o(n_4094) );
na02f80 g768927 ( .a(n_11600), .b(n_11664), .o(n_11821) );
na02f80 g767020 ( .a(FE_OCP_RBN2457_n_13765), .b(n_13787), .o(n_13863) );
in01f80 g774873 ( .a(n_6247), .o(n_6236) );
na02f80 g761431 ( .a(n_18869), .b(FE_OCPN1384_n_18345), .o(n_18924) );
in01f80 g759264 ( .a(n_20984), .o(n_20985) );
ao12f80 g768986 ( .a(n_11860), .b(FE_OCP_RBN2119_n_45224), .c(delay_xor_ln22_unr9_stage4_stallmux_q_9_), .o(n_11900) );
na02f80 g746590 ( .a(n_34666), .b(n_34228), .o(n_34775) );
no02f80 g778339 ( .a(n_2506), .b(n_2573), .o(n_2667) );
na02f80 g753359 ( .a(n_27012), .b(n_27027), .o(n_27070) );
in01f80 g753076 ( .a(n_27190), .o(n_27191) );
no02f80 FE_RC_3121_0 ( .a(FE_OCP_RBN1715_n_20734), .b(n_20862), .o(FE_RN_1383_0) );
in01f80 g765529 ( .a(n_15873), .o(n_15821) );
in01f80 FE_RC_2185_0 ( .a(n_22793), .o(FE_RN_781_0) );
ao12f80 g773907 ( .a(n_6884), .b(n_6883), .c(n_6882), .o(n_6952) );
na02f80 g776365 ( .a(n_47007), .b(n_4662), .o(n_4727) );
in01f80 FE_OCP_RBC2276_n_24077 ( .a(n_24077), .o(FE_OCP_RBN2276_n_24077) );
na02f80 g745422 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35653), .o(n_35723) );
in01f80 newInst_2999 ( .a(newNet_2998), .o(newNet_2999) );
no02f80 g764453 ( .a(n_16218), .b(FE_OCP_RBN2591_n_14460), .o(n_16272) );
no02f80 g739377 ( .a(n_40724), .b(n_40721), .o(n_41234) );
no02f80 g759755 ( .a(n_21450), .b(n_20871), .o(n_21449) );
no02f80 g746265 ( .a(n_33529), .b(n_33080), .o(n_33550) );
no02f80 g753263 ( .a(n_27287), .b(n_27170), .o(n_27332) );
in01f80 fopt782903 ( .a(n_32966), .o(n_44347) );
na02f80 g763111 ( .a(n_17482), .b(n_17407), .o(n_17553) );
na02f80 g778140 ( .a(n_2930), .b(n_2929), .o(n_2999) );
no02f80 g748247 ( .a(FE_OCP_RBN3734_n_31819), .b(FE_OCP_RBN1297_n_30451), .o(n_32056) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_31_ ( .ck(newNet_2720), .d(n_17687), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_) );
no02f80 FE_RC_2545_0 ( .a(FE_RN_1040_0), .b(FE_RN_1041_0), .o(FE_RN_1042_0) );
no02f80 g769640 ( .a(n_11301), .b(FE_OCPN3182_FE_OCP_RBN2831_n_10198), .o(n_11351) );
in01f80 g767367 ( .a(n_13468), .o(n_13540) );
no02f80 g758274 ( .a(FE_OCPN992_n_22249), .b(FE_OCP_RBN1717_n_20734), .o(n_22411) );
no02f80 g762221 ( .a(n_18698), .b(n_18536), .o(n_18731) );
in01f80 FE_RC_2191_0 ( .a(n_14951), .o(FE_RN_785_0) );
na02f80 g748518 ( .a(n_32676), .b(n_32497), .o(n_32726) );
no02f80 g742735 ( .a(n_37320), .b(n_37319), .o(n_37321) );
oa22f80 g784551 ( .a(FE_OFN801_n_46285), .b(n_11252), .c(FE_OCP_RBN3044_n_46337), .d(n_11220), .o(n_46372) );
no02f80 g763919 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n_17297) );
in01f80 FE_OCPUNCOC1804_n_18111 ( .a(FE_OCPUNCON1803_n_18111), .o(FE_OCPUNCON1804_n_18111) );
na02f80 g751289 ( .a(n_29721), .b(n_29202), .o(n_29744) );
na02f80 g756712 ( .a(n_23502), .b(delay_add_ln22_unr14_stage6_stallmux_q_14_), .o(n_23517) );
na02f80 g741875 ( .a(n_38205), .b(n_38122), .o(n_38363) );
in01f80 g759988 ( .a(n_20582), .o(n_20583) );
in01f80 newInst_427 ( .a(newNet_426), .o(newNet_427) );
no02f80 g775454 ( .a(n_5812), .b(n_5891), .o(n_5822) );
in01f80 newInst_3584 ( .a(newNet_3062), .o(newNet_3584) );
na02f80 g753325 ( .a(n_26970), .b(n_26755), .o(n_26991) );
in01f80 g749438 ( .a(n_30692), .o(n_30693) );
in01f80 g742564 ( .a(n_37575), .o(n_38032) );
no02f80 g763692 ( .a(n_16739), .b(FE_OCP_RBN2787_n_15079), .o(n_16760) );
na02f80 g755416 ( .a(n_24783), .b(n_24806), .o(n_24868) );
in01f80 g741215 ( .a(n_39228), .o(n_39229) );
no02f80 g742002 ( .a(n_38332), .b(n_38282), .o(n_38396) );
in01f80 newInst_87 ( .a(newNet_86), .o(newNet_87) );
in01f80 g764090 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17255) );
oa12f80 g777043 ( .a(n_3904), .b(n_3903), .c(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n_4031) );
na02f80 g766317 ( .a(n_14272), .b(n_13515), .o(n_14368) );
no02f80 g737680 ( .a(n_42285), .b(n_42053), .o(n_42505) );
no02f80 g757979 ( .a(n_22345), .b(n_22344), .o(n_22346) );
no02f80 g755706 ( .a(n_24520), .b(n_24519), .o(n_24547) );
in01f80 g737580 ( .a(n_42425), .o(n_42426) );
in01f80 newInst_3260 ( .a(newNet_3259), .o(newNet_3260) );
in01f80 g780797 ( .a(n_412), .o(n_422) );
ao12f80 g743068 ( .a(n_37092), .b(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .o(n_37479) );
ao22s80 g773847 ( .a(n_7028), .b(n_6927), .c(n_7015), .d(n_6926), .o(n_7090) );
in01f80 g747995 ( .a(n_32081), .o(n_32109) );
na02f80 g773097 ( .a(n_7627), .b(n_7611), .o(n_7685) );
ao12f80 g752312 ( .a(n_27830), .b(n_27829), .c(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n_29109) );
no02f80 g759717 ( .a(n_20677), .b(n_18974), .o(n_20716) );
oa12f80 g756346 ( .a(n_24030), .b(n_24453), .c(n_24026), .o(n_24478) );
in01f80 FE_OCP_RBC2943_n_5454 ( .a(n_5454), .o(FE_OCP_RBN2943_n_5454) );
ao12f80 g746853 ( .a(n_32995), .b(n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n_33017) );
no02f80 g737051 ( .a(n_43171), .b(n_43102), .o(n_43204) );
in01f80 g764146 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_), .o(n_18152) );
in01f80 newInst_559 ( .a(newNet_558), .o(newNet_559) );
in01f80 g754904 ( .a(n_25275), .o(n_25358) );
in01f80 g748797 ( .a(n_32425), .o(n_32426) );
na02f80 g738591 ( .a(n_41561), .b(n_41662), .o(n_42032) );
in01f80 newInst_1429 ( .a(newNet_1428), .o(newNet_1429) );
no02f80 g743429 ( .a(n_36669), .b(n_36750), .o(n_36670) );
in01f80 newInst_2520 ( .a(newNet_2519), .o(newNet_2520) );
in01f80 g767895 ( .a(n_13040), .o(n_13041) );
in01f80 FE_OCP_RBC2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01f80 FE_OCPC1255_n_8499 ( .a(FE_OCPN1254_n_8499), .o(FE_OCPN1255_n_8499) );
na02f80 g743257 ( .a(n_35466), .b(delay_sub_ln21_unr24_stage9_stallmux_q_2_), .o(n_36884) );
na02f80 g741785 ( .a(n_38526), .b(n_39230), .o(n_38527) );
in01f80 g759996 ( .a(n_20710), .o(n_20711) );
na02f80 g742888 ( .a(n_37007), .b(n_46254), .o(n_37128) );
in01f80 newInst_1198 ( .a(newNet_1197), .o(newNet_1198) );
no02f80 g759943 ( .a(n_21374), .b(n_21514), .o(n_21600) );
in01f80 g751020 ( .a(n_30034), .o(n_30035) );
na02f80 g779050 ( .a(n_2105), .b(n_2088), .o(n_2089) );
in01f80 g771768 ( .a(n_9127), .o(n_9128) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_16_ ( .ck(newNet_838), .d(n_1304), .o(delay_xor_ln21_unr3_stage2_stallmux_q_16_) );
in01f80 g738307 ( .a(n_41796), .o(n_41797) );
in01f80 g761308 ( .a(n_19005), .o(n_19006) );
no02f80 FE_RC_2742_0 ( .a(n_37662), .b(n_37661), .o(FE_RN_1164_0) );
in01f80 g780493 ( .a(n_1057), .o(n_1058) );
in01f80 g752544 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_), .o(n_27623) );
na02f80 g748298 ( .a(n_31681), .b(n_31682), .o(n_31706) );
no02f80 g757055 ( .a(n_23646), .b(n_23645), .o(n_23704) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_26_ ( .ck(newNet_2838), .d(n_12158), .o(delay_add_ln22_unr8_stage4_stallmux_q_26_) );
in01f80 FE_OCP_RBC2393_n_8288 ( .a(n_8288), .o(FE_OCP_RBN2393_n_8288) );
in01f80 g777817 ( .a(n_3375), .o(n_3370) );
no02f80 g778528 ( .a(n_2318), .b(n_2317), .o(n_2319) );
oa12f80 g750714 ( .a(n_29189), .b(n_29299), .c(n_29190), .o(n_29322) );
na02f80 g739155 ( .a(n_40895), .b(n_41009), .o(n_41012) );
oa12f80 g754760 ( .a(n_25306), .b(n_26106), .c(n_25191), .o(n_26132) );
in01f80 g752854 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_9_), .o(n_28305) );
oa22f80 g748089 ( .a(n_31550), .b(n_31525), .c(n_31551), .d(n_31524), .o(n_31670) );
no02f80 g760115 ( .a(n_20289), .b(n_47257), .o(n_20337) );
no02f80 g754754 ( .a(n_25336), .b(n_25335), .o(n_25337) );
ms00f80 cos_out_reg_11_ ( .ck(newNet_3751), .d(n_43797), .o(cos_out_11) );
in01f80 FE_OCP_RBC3030_n_39942 ( .a(FE_OCP_RBN3027_n_39942), .o(FE_OCP_RBN3030_n_39942) );
in01f80 g747685 ( .a(n_32324), .o(n_32343) );
in01f80 g745805 ( .a(n_34146), .o(n_34414) );
na02f80 g780467 ( .a(n_708), .b(n_707), .o(n_709) );
no02f80 g769056 ( .a(FE_OCP_RBN2119_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_8_), .o(n_11756) );
na02f80 g765112 ( .a(n_15277), .b(n_15310), .o(n_15463) );
no02f80 g761756 ( .a(n_18518), .b(n_18215), .o(n_18647) );
ao22s80 FE_RC_1275_0 ( .a(n_2810), .b(n_3635), .c(n_2809), .d(n_3579), .o(n_3718) );
oa12f80 g756334 ( .a(n_24003), .b(n_24002), .c(n_24001), .o(n_24054) );
in01f80 newInst_2488 ( .a(newNet_375), .o(newNet_2488) );
no02f80 g744463 ( .a(n_35470), .b(n_35469), .o(n_35502) );
na02f80 g744254 ( .a(n_44174), .b(n_36091), .o(n_35571) );
no02f80 g775626 ( .a(n_5661), .b(n_5626), .o(n_5701) );
in01f80 g772506 ( .a(n_8448), .o(n_8449) );
na02f80 g752529 ( .a(n_27621), .b(n_27609), .o(n_27693) );
in01f80 g771601 ( .a(n_9396), .o(n_9470) );
in01f80 FE_OCP_RBC3656_n_25997 ( .a(n_25997), .o(FE_OCP_RBN3656_n_25997) );
ao12f80 g748073 ( .a(n_32866), .b(n_32865), .c(n_32864), .o(n_33441) );
no02f80 g780633 ( .a(n_662), .b(n_413), .o(n_659) );
na02f80 g745371 ( .a(FE_OCP_RBN2987_n_35539), .b(n_35371), .o(n_35890) );
in01f80 newInst_750 ( .a(newNet_77), .o(newNet_750) );
na02f80 g773795 ( .a(n_7182), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .o(n_7233) );
ao22s80 g757522 ( .a(n_22686), .b(n_22343), .c(n_22720), .d(n_22306), .o(n_22755) );
no02f80 g749033 ( .a(n_30918), .b(n_30917), .o(n_30947) );
oa22f80 g779895 ( .a(n_44652), .b(n_1019), .c(n_44623), .d(n_947), .o(n_1320) );
in01f80 g775016 ( .a(n_6184), .o(n_6185) );
no03m80 FE_RC_609_0 ( .a(n_40828), .b(n_40909), .c(n_40908), .o(n_40910) );
no02f80 g756142 ( .a(n_24818), .b(n_24193), .o(n_24906) );
na02f80 g775516 ( .a(n_5272), .b(n_5022), .o(n_5348) );
in01f80 g765183 ( .a(n_15235), .o(n_15236) );
in01f80 FE_RC_811_0 ( .a(n_28701), .o(FE_RN_243_0) );
in01f80 g746413 ( .a(n_33409), .o(n_33410) );
na02f80 g765169 ( .a(n_15579), .b(FE_OCP_RBN3622_n_15135), .o(n_15639) );
no02f80 g760291 ( .a(n_20173), .b(n_20193), .o(n_20245) );
no03m80 g737562 ( .a(n_42468), .b(n_42419), .c(n_42467), .o(n_42492) );
no02f80 g768091 ( .a(n_12914), .b(n_12909), .o(n_13150) );
na02f80 g751776 ( .a(n_29008), .b(n_28945), .o(n_29047) );
no02f80 FE_RC_1988_0 ( .a(FE_RN_648_0), .b(n_13732), .o(n_13774) );
no02f80 g775806 ( .a(n_5407), .b(n_5435), .o(n_5549) );
oa12f80 g753611 ( .a(n_26495), .b(n_26623), .c(n_26559), .o(n_26701) );
no02f80 g769222 ( .a(n_11585), .b(n_45300), .o(n_11589) );
na02f80 g742798 ( .a(n_37258), .b(n_37127), .o(n_37514) );
in01f80 newInst_960 ( .a(newNet_959), .o(newNet_960) );
in01f80 FE_OCP_RBC1376_n_20889 ( .a(n_20889), .o(FE_OCP_RBN1376_n_20889) );
in01f80 g755963 ( .a(n_29630), .o(n_25859) );
na02f80 g753738 ( .a(n_26379), .b(n_26447), .o(n_26524) );
in01f80 newInst_3186 ( .a(newNet_2022), .o(newNet_3186) );
in01f80 newInst_935 ( .a(newNet_934), .o(newNet_935) );
na02f80 g784411 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_), .o(n_46223) );
no02f80 g767804 ( .a(n_13064), .b(n_13210), .o(n_13202) );
na02f80 g759169 ( .a(n_20951), .b(n_45013), .o(n_21016) );
no02f80 g778446 ( .a(FE_OCP_RBN2285_n_2433), .b(n_2341), .o(n_2538) );
in01f80 g760897 ( .a(n_20265), .o(n_20266) );
no02f80 g767889 ( .a(n_12677), .b(n_13889), .o(n_12865) );
na02f80 g778290 ( .a(n_2548), .b(n_2647), .o(n_2725) );
na02f80 g744630 ( .a(n_35273), .b(n_35266), .o(n_35328) );
in01f80 g772013 ( .a(n_9433), .o(n_9505) );
no02f80 g738724 ( .a(n_41386), .b(n_41385), .o(n_41399) );
in01f80 newInst_2584 ( .a(newNet_1188), .o(newNet_2584) );
na03f80 g752638 ( .a(n_28204), .b(n_28205), .c(n_27926), .o(n_28239) );
in01f80 g778292 ( .a(n_2674), .o(n_3378) );
in01f80 FE_OCP_DRV_C3150_n_12773 ( .a(FE_OCP_DRV_N3149_n_12773), .o(FE_OCP_DRV_N3150_n_12773) );
in01f80 newInst_893 ( .a(newNet_420), .o(newNet_893) );
no02f80 g773669 ( .a(n_7320), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .o(n_7341) );
in01f80 newInst_877 ( .a(newNet_876), .o(newNet_877) );
ao12f80 g743053 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_37017) );
na02f80 g776606 ( .a(n_4389), .b(n_4122), .o(n_4430) );
in01f80 g772343 ( .a(n_8629), .o(n_8630) );
no02f80 g752150 ( .a(n_28065), .b(n_28064), .o(n_28090) );
in01f80 newInst_3042 ( .a(newNet_90), .o(newNet_3042) );
in01f80 newInst_2603 ( .a(newNet_1095), .o(newNet_2603) );
no02f80 g778279 ( .a(n_2623), .b(n_2622), .o(n_2669) );
no02f80 g761691 ( .a(n_18791), .b(n_18746), .o(n_18856) );
in01f80 g742962 ( .a(n_37054), .o(n_37055) );
no02f80 g740654 ( .a(n_39583), .b(n_45840), .o(n_39610) );
in01f80 g779566 ( .a(n_1599), .o(n_1600) );
in01f80 g778304 ( .a(n_44059), .o(n_2579) );
no02f80 g768026 ( .a(n_12914), .b(n_12964), .o(n_12992) );
in01f80 g758720 ( .a(n_21687), .o(n_21738) );
in01f80 newInst_166 ( .a(newNet_9), .o(newNet_166) );
in01f80 g756190 ( .a(n_24147), .o(n_24145) );
na02f80 g772818 ( .a(n_8122), .b(n_8053), .o(n_8180) );
in01f80 g749724 ( .a(n_31431), .o(n_31432) );
ao22s80 g756949 ( .a(n_23803), .b(n_23869), .c(n_24059), .d(n_23812), .o(n_24170) );
in01f80 g761815 ( .a(n_18554), .o(n_18555) );
no02f80 g743843 ( .a(n_36043), .b(n_35909), .o(n_36072) );
no02f80 g771978 ( .a(n_44575), .b(FE_OCP_RBN2540_n_8781), .o(n_9019) );
ao22s80 FE_RC_245_0 ( .a(n_19061), .b(n_18638), .c(n_19060), .d(n_18637), .o(n_19177) );
in01f80 g743811 ( .a(n_37246), .o(n_37247) );
ao12f80 g761829 ( .a(n_18786), .b(n_18672), .c(n_18355), .o(n_18787) );
in01f80 FE_RC_3007_0 ( .a(FE_RN_1317_0), .o(n_30935) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_11_ ( .ck(newNet_195), .d(n_46369), .o(delay_xor_ln22_unr9_stage4_stallmux_q_11_) );
in01f80 g750366 ( .a(n_30687), .o(n_30688) );
na02f80 FE_RC_1747_0 ( .a(n_12317), .b(FE_RN_491_0), .o(FE_RN_492_0) );
in01f80 FE_OCP_RBC1190_n_14911 ( .a(n_14911), .o(FE_OCP_RBN1190_n_14911) );
na02f80 g780906 ( .a(n_403), .b(n_417), .o(n_432) );
in01f80 FE_OCPC3187_n_11012 ( .a(n_11012), .o(FE_OCPN3187_n_11012) );
in01f80 FE_RC_478_0 ( .a(n_23165), .o(FE_RN_142_0) );
no02f80 g746453 ( .a(n_33381), .b(n_33190), .o(n_33468) );
in01f80 g760624 ( .a(n_19835), .o(n_19836) );
ao12f80 g770523 ( .a(n_10265), .b(FE_OCP_RBN2876_n_10354), .c(n_10313), .o(n_10499) );
no02f80 g745316 ( .a(n_35605), .b(n_35562), .o(n_35656) );
na03f80 g743149 ( .a(n_37201), .b(n_45896), .c(n_37224), .o(n_38221) );
oa12f80 g780715 ( .a(n_625), .b(n_626), .c(n_624), .o(n_748) );
no02f80 g765360 ( .a(n_15038), .b(n_15108), .o(n_15126) );
in01f80 newInst_569 ( .a(newNet_319), .o(newNet_569) );
in01f80 g738714 ( .a(n_41419), .o(n_41440) );
in01f80 g754231 ( .a(n_26014), .o(n_26015) );
na02f80 g761908 ( .a(n_18704), .b(n_17749), .o(n_18915) );
in01f80 g766737 ( .a(n_13774), .o(n_13806) );
in01f80 g773280 ( .a(n_7617), .o(n_7712) );
no02f80 g755841 ( .a(n_24271), .b(n_24294), .o(n_24366) );
no02f80 g748747 ( .a(n_32461), .b(n_32489), .o(n_32505) );
in01f80 g754933 ( .a(n_25239), .o(n_25397) );
in01f80 g738731 ( .a(n_41532), .o(n_41557) );
no02f80 g767320 ( .a(n_13622), .b(n_13346), .o(n_13696) );
no02f80 g760999 ( .a(n_19216), .b(n_19252), .o(n_19360) );
no02f80 g771060 ( .a(n_9359), .b(n_8232), .o(n_9461) );
in01f80 g745340 ( .a(n_36211), .o(n_36212) );
in01f80 g779496 ( .a(n_2046), .o(n_2047) );
na02f80 g760659 ( .a(n_19802), .b(FE_OCPUNCON1806_n_19801), .o(n_19882) );
no02f80 g777085 ( .a(n_3755), .b(n_3637), .o(n_3795) );
in01f80 g772207 ( .a(n_8782), .o(n_8783) );
na02f80 g776096 ( .a(n_4981), .b(n_5052), .o(n_5290) );
in01f80 FE_RC_3201_0 ( .a(n_7579), .o(FE_RN_1422_0) );
no02f80 g771656 ( .a(n_8850), .b(n_8637), .o(n_8912) );
na02f80 g736412 ( .a(n_43790), .b(n_43682), .o(n_43819) );
oa12f80 g754488 ( .a(n_25277), .b(n_25433), .c(n_25243), .o(n_25545) );
no02f80 g778999 ( .a(n_2172), .b(n_2164), .o(n_2165) );
in01f80 g758890 ( .a(n_21507), .o(n_21501) );
no02f80 g738116 ( .a(n_42046), .b(n_42500), .o(n_42045) );
na02f80 g771841 ( .a(n_9826), .b(n_9873), .o(n_10816) );
in01f80 g739042 ( .a(n_41494), .o(n_41123) );
in01f80 FE_OCP_RBC1138_n_11779 ( .a(n_11779), .o(FE_OCP_RBN1138_n_11779) );
na02f80 g745811 ( .a(n_44100), .b(n_33517), .o(n_34144) );
in01f80 newInst_2036 ( .a(newNet_2035), .o(newNet_2036) );
in01f80 FE_OCP_RBC3837_n_19513 ( .a(n_19513), .o(FE_OCP_RBN3837_n_19513) );
in01f80 FE_RC_2036_0 ( .a(n_26666), .o(FE_RN_680_0) );
no02f80 g762642 ( .a(n_17932), .b(n_17931), .o(n_17952) );
na02f80 g752332 ( .a(n_27893), .b(n_27885), .o(n_27970) );
ao22s80 FE_RC_98_0 ( .a(n_18240), .b(n_18563), .c(n_18241), .d(n_18562), .o(n_18713) );
in01f80 g743674 ( .a(n_36427), .o(n_36428) );
na02f80 g764568 ( .a(n_15816), .b(n_14650), .o(n_15918) );
ao22s80 g779509 ( .a(n_1368), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(n_1358), .d(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .o(n_1446) );
in01f80 g740704 ( .a(n_40005), .o(n_39599) );
ao12f80 g760598 ( .a(n_19750), .b(n_19701), .c(n_19809), .o(n_19817) );
no02f80 g760543 ( .a(n_19894), .b(n_19893), .o(n_19921) );
in01f80 g781393 ( .a(beta_6), .o(n_67) );
na02f80 g772832 ( .a(n_8008), .b(n_8033), .o(n_8136) );
no02f80 FE_RC_2392_0 ( .a(FE_RN_938_0), .b(n_42738), .o(FE_RN_939_0) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_21_ ( .ck(newNet_1995), .d(n_11655), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_) );
in01f80 g759254 ( .a(n_21216), .o(n_22134) );
in01f80 g778889 ( .a(n_2289), .o(n_2365) );
ao22s80 FE_RC_1588_0 ( .a(n_11958), .b(n_11755), .c(n_11754), .d(n_11874), .o(n_12037) );
na02f80 g779206 ( .a(n_1847), .b(n_1730), .o(n_1839) );
in01f80 FE_RC_910_0 ( .a(FE_RN_269_0), .o(n_12022) );
oa22f80 FE_RC_1449_0 ( .a(n_32566), .b(n_32340), .c(n_28336), .d(n_32309), .o(n_32374) );
no02f80 FE_RC_2280_0 ( .a(FE_RN_851_0), .b(n_28176), .o(FE_RN_852_0) );
na02f80 g742871 ( .a(n_37184), .b(n_37210), .o(n_37445) );
oa12f80 g741459 ( .a(n_38744), .b(n_38780), .c(n_38760), .o(n_38801) );
no02f80 g760155 ( .a(n_20537), .b(FE_OCP_RBN2419_n_19601), .o(n_20662) );
oa12f80 g740871 ( .a(n_39236), .b(n_44312), .c(n_39192), .o(n_39440) );
in01f80 g744667 ( .a(n_35340), .o(n_35341) );
na02f80 g767271 ( .a(n_13409), .b(n_12847), .o(n_13432) );
na03f80 FE_RC_1_0 ( .a(beta_31), .b(beta_11), .c(n_206), .o(n_207) );
na02f80 g750477 ( .a(n_29572), .b(n_29571), .o(n_29587) );
in01f80 g741537 ( .a(n_38703), .o(n_38717) );
no02f80 g780764 ( .a(n_506), .b(n_410), .o(n_547) );
in01f80 g749452 ( .a(n_30537), .o(n_30559) );
no02f80 g751171 ( .a(n_29932), .b(n_30063), .o(n_30092) );
in01f80 FE_RC_1204_0 ( .a(n_17489), .o(FE_RN_364_0) );
na02f80 g771834 ( .a(n_9386), .b(n_9475), .o(n_9815) );
na02f80 g757030 ( .a(n_23700), .b(n_23645), .o(n_23832) );
na02f80 g760696 ( .a(FE_OCP_RBN2418_n_19601), .b(n_18140), .o(n_19669) );
in01f80 FE_OCPC1036_n_28288 ( .a(FE_OCPN1035_n_28288), .o(FE_OCPN1036_n_28288) );
in01f80 g768080 ( .a(n_12982), .o(n_12916) );
in01f80 g760992 ( .a(n_19414), .o(n_19454) );
na02f80 FE_RC_4225_0 ( .a(FE_RN_1853_0), .b(n_29929), .o(FE_RN_1854_0) );
oa22f80 FE_RC_259_0 ( .a(n_14907), .b(n_14965), .c(n_14964), .d(n_14924), .o(n_15083) );
in01f80 g737240 ( .a(FE_OCP_RBN3000_n_42959), .o(n_42967) );
na02f80 g752616 ( .a(FE_OCP_RBN3736_n_27535), .b(n_27430), .o(n_27571) );
in01f80 g775189 ( .a(n_6066), .o(n_6087) );
na02f80 g745267 ( .a(n_35852), .b(FE_OCP_RBN2992_n_35539), .o(n_35939) );
oa22f80 g764137 ( .a(n_16819), .b(n_16250), .c(n_16818), .d(n_16249), .o(n_16926) );
ao12f80 g761389 ( .a(n_19576), .b(n_19613), .c(n_19575), .o(n_19678) );
no02f80 g779752 ( .a(n_1379), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_16_), .o(n_1508) );
no02f80 g746802 ( .a(n_33061), .b(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(n_33062) );
oa22f80 g781279 ( .a(n_18), .b(n_46055), .c(n_7), .d(beta_20), .o(n_246) );
na02f80 g764571 ( .a(n_15910), .b(n_14452), .o(n_16005) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_9_ ( .ck(newNet_941), .d(n_22815), .o(delay_xor_ln21_unr15_stage6_stallmux_q_9_) );
na02f80 FE_RC_1893_0 ( .a(n_11879), .b(n_12121), .o(FE_RN_591_0) );
in01f80 newInst_2278 ( .a(newNet_2277), .o(newNet_2278) );
in01f80 newInst_2513 ( .a(newNet_2512), .o(newNet_2513) );
na02f80 g750615 ( .a(n_29516), .b(n_29467), .o(n_29559) );
in01f80 g781243 ( .a(n_149), .o(n_150) );
no02f80 g772526 ( .a(n_8454), .b(n_8453), .o(n_8487) );
na02f80 g764447 ( .a(n_16220), .b(n_14730), .o(n_16221) );
no02f80 g780622 ( .a(n_713), .b(n_734), .o(n_781) );
in01f80 g777878 ( .a(n_3212), .o(n_3228) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_7_ ( .ck(newNet_2047), .d(n_5363), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_) );
in01f80 g771138 ( .a(n_9663), .o(n_9741) );
in01f80 FE_RC_4047_0 ( .a(n_35591), .o(FE_RN_1758_0) );
in01f80 g766001 ( .a(n_14798), .o(n_14764) );
in01f80 newInst_2004 ( .a(newNet_2003), .o(newNet_2004) );
in01f80 newInst_1446 ( .a(newNet_508), .o(newNet_1446) );
in01f80 g779055 ( .a(n_2163), .o(n_2147) );
no02f80 FE_RC_2972_0 ( .a(FE_OCP_DRV_N1598_n_35644), .b(n_34707), .o(FE_RN_1300_0) );
oa22f80 g739843 ( .a(n_40232), .b(n_40294), .c(n_40233), .d(n_40293), .o(n_40403) );
na02f80 g771379 ( .a(n_9247), .b(FE_OCP_RBN3543_n_44575), .o(n_9294) );
no02f80 g742256 ( .a(n_44866), .b(n_37901), .o(n_37902) );
in01f80 newInst_923 ( .a(newNet_446), .o(newNet_923) );
ao12f80 g775883 ( .a(n_5002), .b(n_5140), .c(n_4979), .o(n_5233) );
no02f80 g759893 ( .a(n_21141), .b(n_21140), .o(n_21142) );
in01f80 newInst_1899 ( .a(newNet_768), .o(newNet_1899) );
oa22f80 FE_RC_1655_0 ( .a(n_24350), .b(n_27781), .c(n_27796), .d(n_27752), .o(n_27838) );
na02f80 g776339 ( .a(n_4560), .b(n_4548), .o(n_4667) );
no02f80 FE_RC_1803_0 ( .a(FE_OCP_RBN2595_n_25181), .b(FE_RN_533_0), .o(n_25401) );
in01f80 newInst_1553 ( .a(newNet_616), .o(newNet_1553) );
in01f80 g762767 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .o(n_17824) );
no02f80 g754965 ( .a(n_25803), .b(n_25802), .o(n_25804) );
na02f80 g745392 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35842), .o(n_35841) );
in01f80 g745356 ( .a(n_36209), .o(n_36210) );
na02f80 g767623 ( .a(n_12803), .b(n_12849), .o(n_12888) );
na02f80 g766034 ( .a(n_14615), .b(n_14472), .o(n_14750) );
na02f80 g744307 ( .a(n_44180), .b(n_35113), .o(n_36058) );
oa12f80 g745208 ( .a(n_36227), .b(n_36226), .c(n_36225), .o(n_36282) );
na02f80 g768465 ( .a(n_12419), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .o(n_12474) );
in01f80 g739414 ( .a(n_40726), .o(n_40727) );
na02f80 g765785 ( .a(n_14950), .b(n_14210), .o(n_15008) );
no02f80 g739950 ( .a(n_40228), .b(n_40083), .o(n_40257) );
ao12f80 g750291 ( .a(n_29707), .b(n_29720), .c(n_29706), .o(n_31327) );
in01f80 newInst_2128 ( .a(newNet_2127), .o(newNet_2128) );
na02f80 g738361 ( .a(n_41551), .b(n_41520), .o(n_41521) );
no02f80 g766079 ( .a(n_14585), .b(n_13329), .o(n_14611) );
na02f80 g771257 ( .a(n_9348), .b(n_9289), .o(n_9453) );
na02f80 g737058 ( .a(FE_OCP_RBN3729_n_43230), .b(n_42878), .o(n_43515) );
ao22s80 g756535 ( .a(n_23821), .b(n_22873), .c(n_23783), .d(delay_sub_ln21_0_unr14_stage6_stallmux_q_31_), .o(n_23962) );
ao12f80 g751725 ( .a(n_29247), .b(n_29246), .c(n_29245), .o(n_30038) );
oa12f80 g738095 ( .a(n_41731), .b(n_42070), .c(n_41670), .o(n_42087) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_2_ ( .ck(newNet_2361), .d(n_35419), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_) );
na02f80 g773193 ( .a(n_7650), .b(n_8444), .o(n_7672) );
in01f80 g757304 ( .a(n_23167), .o(n_23168) );
in01f80 FE_OCPC1013_n_41478 ( .a(FE_OCPN1012_n_41478), .o(FE_OCPN1013_n_41478) );
in01f80 newInst_3287 ( .a(newNet_3286), .o(newNet_3287) );
na02f80 g766247 ( .a(n_14374), .b(n_14409), .o(n_14547) );
na02f80 g736727 ( .a(n_43087), .b(n_43092), .o(n_43234) );
no02f80 g746534 ( .a(n_34808), .b(n_34692), .o(n_35355) );
in01f80 newInst_843 ( .a(newNet_398), .o(newNet_843) );
na02f80 g773875 ( .a(n_7107), .b(n_7106), .o(n_7283) );
na02f80 g771779 ( .a(n_9124), .b(FE_OCP_RBN3546_n_44575), .o(n_9228) );
na02f80 g741914 ( .a(n_38170), .b(n_38317), .o(n_38319) );
no02f80 g765293 ( .a(n_15961), .b(n_15874), .o(n_16099) );
in01f80 g736482 ( .a(n_43739), .o(n_43740) );
in01f80 g742619 ( .a(n_37619), .o(n_37589) );
oa12f80 g755916 ( .a(n_25253), .b(n_25160), .c(n_25135), .o(n_25708) );
in01f80 g773253 ( .a(n_7599), .o(n_7615) );
no02f80 FE_RC_3122_0 ( .a(FE_RN_1383_0), .b(FE_OCP_RBN3221_n_22068), .o(n_22304) );
na02f80 g770681 ( .a(n_10145), .b(n_10186), .o(n_10263) );
in01f80 g750882 ( .a(n_29136), .o(n_29137) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_16_ ( .ck(newNet_1243), .d(n_5753), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_) );
in01f80 g761183 ( .a(n_19797), .o(n_19798) );
no02f80 g741579 ( .a(n_38669), .b(n_38668), .o(n_38670) );
in01f80 g745122 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .o(n_36355) );
in01f80 newInst_2726 ( .a(newNet_2725), .o(newNet_2726) );
oa22f80 g748512 ( .a(n_31402), .b(n_31385), .c(n_31401), .d(n_31426), .o(n_31470) );
no02f80 g754744 ( .a(FE_OCP_RBN2957_n_26231), .b(n_25746), .o(n_26484) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_19_ ( .ck(newNet_830), .d(n_1334), .o(delay_xor_ln21_unr3_stage2_stallmux_q_19_) );
in01f80 g759633 ( .a(n_20756), .o(n_20757) );
no02f80 g758701 ( .a(n_21688), .b(n_21689), .o(n_21744) );
oa22f80 g756956 ( .a(n_23803), .b(n_24111), .c(n_24059), .d(n_23807), .o(n_24237) );
in01f80 g754405 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .o(n_27988) );
in01f80 fopt783141 ( .a(n_44672), .o(n_44637) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_31_ ( .ck(newNet_1477), .d(n_32293), .o(delay_sub_ln23_unr25_stage8_stallmux_q_3_) );
ao22s80 g768998 ( .a(FE_OCP_RBN3268_n_45224), .b(n_11595), .c(FE_OCP_RBN2113_n_45224), .d(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n_11767) );
na02f80 g778079 ( .a(n_2939), .b(n_2949), .o(n_4642) );
in01f80 g768077 ( .a(n_12854), .o(n_12813) );
in01f80 g736999 ( .a(n_43339), .o(n_43390) );
oa22f80 FE_RC_1054_0 ( .a(n_36739), .b(n_36760), .c(n_36740), .d(n_36759), .o(n_36792) );
no02f80 g747409 ( .a(n_32595), .b(n_32522), .o(n_32523) );
in01f80 g742463 ( .a(n_37690), .o(n_37754) );
na02f80 g745718 ( .a(n_34218), .b(n_44102), .o(n_34260) );
ao12f80 g749617 ( .a(n_30446), .b(FE_OCP_RBN1357_n_30298), .c(n_30444), .o(n_30526) );
no02f80 g756769 ( .a(n_23476), .b(n_23475), .o(n_23496) );
in01f80 g776326 ( .a(n_4823), .o(n_4824) );
oa22f80 g774389 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .c(FE_OCPN895_n_6521), .d(n_5104), .o(n_7110) );
oa12f80 g739107 ( .a(n_41056), .b(n_41055), .c(n_41054), .o(n_41392) );
no02f80 g757239 ( .a(n_23469), .b(n_22845), .o(n_23470) );
na02f80 g753131 ( .a(n_27326), .b(n_27393), .o(n_27394) );
in01f80 FE_RC_3575_0 ( .a(FE_RN_1555_0), .o(n_35869) );
oa22f80 FE_RC_3211_0 ( .a(n_1205), .b(n_44659), .c(n_1200), .d(n_44637), .o(n_1354) );
no02f80 g762608 ( .a(n_18039), .b(n_17950), .o(n_18069) );
in01f80 newInst_1854 ( .a(newNet_772), .o(newNet_1854) );
in01f80 g743632 ( .a(n_37538), .o(n_37539) );
no02f80 g744114 ( .a(n_35620), .b(n_35619), .o(n_35640) );
no02f80 FE_RC_2729_0 ( .a(FE_OCP_RBN3827_n_18951), .b(FE_RN_1155_0), .o(n_19088) );
na02f80 g756088 ( .a(n_24306), .b(n_24283), .o(n_24284) );
in01f80 g748337 ( .a(n_31916), .o(n_31917) );
in01f80 newInst_2697 ( .a(newNet_2696), .o(newNet_2697) );
in01f80 g743228 ( .a(n_38128), .o(n_38129) );
in01f80 newInst_1918 ( .a(newNet_1917), .o(newNet_1918) );
na02f80 g767431 ( .a(n_13339), .b(n_13360), .o(n_13397) );
no02f80 g759173 ( .a(n_21218), .b(FE_OCPN1524_n_45072), .o(n_21275) );
no02f80 g777170 ( .a(n_4504), .b(n_4503), .o(n_5131) );
ao12f80 g745276 ( .a(n_34387), .b(n_34386), .c(n_34385), .o(n_35504) );
na02f80 g757256 ( .a(n_23004), .b(n_44071), .o(n_23111) );
na02f80 g766652 ( .a(n_13756), .b(FE_OCPN860_n_12880), .o(n_13783) );
no02f80 g747297 ( .a(n_32731), .b(n_32754), .o(n_32752) );
in01f80 g747270 ( .a(n_32617), .o(n_32643) );
in01f80 g762397 ( .a(n_18499), .o(n_18446) );
in01f80 newInst_1746 ( .a(newNet_1745), .o(newNet_1746) );
ao12f80 g768272 ( .a(n_12552), .b(n_12553), .c(n_12551), .o(n_12585) );
in01f80 FE_RC_2135_0 ( .a(FE_RN_747_0), .o(n_26727) );
ao22s80 FE_RC_3334_0 ( .a(n_18670), .b(n_19477), .c(n_18669), .d(n_19476), .o(n_19599) );
na02f80 FE_RC_1736_0 ( .a(n_37131), .b(FE_RN_483_0), .o(FE_RN_484_0) );
na02f80 FE_RC_2390_0 ( .a(n_42434), .b(FE_RN_936_0), .o(FE_RN_937_0) );
in01f80 g775713 ( .a(n_5459), .o(n_5460) );
in01f80 g749817 ( .a(n_31615), .o(n_31616) );
na02f80 g771400 ( .a(n_9116), .b(n_9201), .o(n_9205) );
no02f80 g743995 ( .a(n_35910), .b(n_36293), .o(n_36363) );
na02f80 g770332 ( .a(n_10405), .b(n_10324), .o(n_10485) );
na02f80 g773956 ( .a(n_7239), .b(n_7276), .o(n_7476) );
na02f80 g744554 ( .a(n_35365), .b(n_35214), .o(n_35366) );
no02f80 g780551 ( .a(FE_OCPN852_n_694), .b(n_420), .o(n_936) );
na02f80 g744244 ( .a(n_46206), .b(n_36810), .o(n_36868) );
in01f80 g757226 ( .a(n_23521), .o(n_23522) );
in01f80 g758590 ( .a(n_21903), .o(n_21904) );
na02f80 g752393 ( .a(n_44420), .b(FE_OCP_RBN3306_n_44722), .o(n_27885) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_1_ ( .ck(newNet_175), .d(n_46387), .o(n_45622) );
in01f80 g744105 ( .a(n_36915), .o(n_36916) );
in01f80 fopt784020 ( .a(n_32280), .o(n_45755) );
no02f80 g778087 ( .a(n_2897), .b(n_2943), .o(n_3597) );
no02f80 g750704 ( .a(n_29364), .b(n_29157), .o(n_29390) );
in01f80 g773345 ( .a(FE_OCP_RBN3468_n_7886), .o(n_8104) );
na02f80 g773084 ( .a(n_7665), .b(n_7668), .o(n_7761) );
na02f80 g762081 ( .a(FE_OCP_RBN2203_n_18242), .b(delay_add_ln22_unr11_stage5_stallmux_q_23_), .o(n_18393) );
oa12f80 g743145 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_37104) );
in01f80 newInst_2235 ( .a(newNet_510), .o(newNet_2235) );
in01f80 g768675 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n_12209) );
in01f80 g760444 ( .a(n_20167), .o(n_20141) );
na02f80 g779234 ( .a(n_1866), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .o(n_1952) );
in01f80 g772964 ( .a(n_8009), .o(n_7953) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_10_ ( .ck(newNet_2129), .d(n_5618), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_) );
oa22f80 FE_RC_3785_0 ( .a(n_36778), .b(n_36754), .c(n_36753), .d(n_36779), .o(n_36830) );
ao12f80 g757726 ( .a(n_23159), .b(n_23158), .c(n_23157), .o(n_23807) );
na02f80 g770185 ( .a(n_10914), .b(n_10979), .o(n_11013) );
in01f80 newInst_792 ( .a(newNet_791), .o(newNet_792) );
na02f80 g755700 ( .a(n_24550), .b(n_24549), .o(n_24551) );
in01f80 g751802 ( .a(n_44045), .o(n_28961) );
na02f80 g749166 ( .a(n_30851), .b(n_30874), .o(n_30991) );
no02f80 g755634 ( .a(n_24566), .b(n_24560), .o(n_24561) );
na02f80 g740234 ( .a(n_39771), .b(n_39752), .o(n_39782) );
na02f80 g742418 ( .a(n_37694), .b(n_37055), .o(n_37708) );
in01f80 FE_OCPC989_n_28353 ( .a(FE_OCPN988_n_28353), .o(FE_OCPN989_n_28353) );
no02f80 g755595 ( .a(n_24568), .b(n_24567), .o(n_24569) );
in01f80 newInst_2856 ( .a(newNet_2855), .o(newNet_2856) );
in01f80 FE_OCP_RBC3361_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3361_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
no02f80 g738763 ( .a(n_41372), .b(n_41337), .o(n_41360) );
in01f80 g771282 ( .a(n_9615), .o(n_9616) );
ao12f80 g757892 ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(n_22854), .c(n_22658), .o(n_22855) );
in01f80 g751824 ( .a(n_28254), .o(n_28291) );
na02f80 g776794 ( .a(n_4169), .b(n_2584), .o(n_4329) );
no02f80 g775578 ( .a(n_5512), .b(n_5476), .o(n_5513) );
na02f80 g757861 ( .a(n_23008), .b(n_22840), .o(n_23060) );
no02f80 g768550 ( .a(FE_OCP_RBN2162_n_12312), .b(n_11888), .o(n_12365) );
ao12f80 g757368 ( .a(n_23229), .b(n_44066), .c(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .o(n_23038) );
na02f80 g771208 ( .a(n_9058), .b(FE_OCP_RBN3476_n_7886), .o(n_9161) );
ms00f80 delay_sub_ln23_0_unr25_stage9_stallmux_q_reg ( .ck(newNet_1456), .d(n_33571), .o(delay_sub_ln23_0_unr25_stage9_stallmux_q) );
in01f80 newInst_2354 ( .a(newNet_2353), .o(newNet_2354) );
na02f80 g776466 ( .a(n_4443), .b(n_4511), .o(n_4671) );
na02f80 g759783 ( .a(n_21670), .b(n_21560), .o(n_21695) );
in01f80 g757575 ( .a(n_22902), .o(n_22862) );
na02f80 g773714 ( .a(n_7321), .b(n_7286), .o(n_7311) );
in01f80 g740373 ( .a(n_39854), .o(n_39940) );
na02f80 g744238 ( .a(n_46223), .b(n_36822), .o(n_36870) );
na02f80 g773784 ( .a(n_7207), .b(n_7166), .o(n_7523) );
no02f80 g751615 ( .a(n_28467), .b(n_27713), .o(n_28510) );
in01f80 FE_OCP_RBC1130_n_24179 ( .a(FE_OCP_RBN1129_n_24179), .o(FE_OCP_RBN1130_n_24179) );
na02f80 g768412 ( .a(n_12401), .b(n_12207), .o(n_12383) );
na02f80 g740203 ( .a(n_39812), .b(n_39461), .o(n_39925) );
oa22f80 g752773 ( .a(n_27089), .b(n_26984), .c(n_27088), .d(n_26983), .o(n_27160) );
oa12f80 g738127 ( .a(n_42022), .b(n_42021), .c(n_42020), .o(n_42072) );
oa12f80 g738449 ( .a(n_41513), .b(FE_OCPN952_n_41540), .c(n_41473), .o(n_41930) );
no02f80 g749774 ( .a(n_31342), .b(n_31219), .o(n_31343) );
ao22s80 g736451 ( .a(n_43690), .b(n_43537), .c(n_43689), .d(n_43536), .o(n_43730) );
no02f80 g770454 ( .a(n_10399), .b(FE_OCP_RBN3600_FE_OCPN1243_n_44460), .o(n_10449) );
oa22f80 g769621 ( .a(n_11342), .b(n_10343), .c(n_11333), .d(n_10344), .o(n_11402) );
in01f80 g749373 ( .a(n_32008), .o(n_32035) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_6_ ( .ck(newNet_2437), .d(n_31514), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_) );
in01f80 g769155 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_6_), .o(n_11595) );
in01f80 g738478 ( .a(n_41642), .o(n_41592) );
ao12f80 g780070 ( .a(n_1016), .b(n_1215), .c(n_1051), .o(n_1228) );
in01f80 g772740 ( .a(n_8235), .o(n_8236) );
oa22f80 g765413 ( .a(FE_OCP_RBN2717_n_14982), .b(FE_OCP_RBN2356_n_13858), .c(FE_OCP_RBN2715_n_14982), .d(n_13950), .o(n_15187) );
in01f80 g747719 ( .a(n_32150), .o(n_32145) );
in01f80 g749113 ( .a(n_32232), .o(n_32233) );
no02f80 g767534 ( .a(n_13006), .b(n_13012), .o(n_13154) );
in01f80 g739709 ( .a(n_40517), .o(n_40518) );
no02f80 g755588 ( .a(n_24683), .b(n_24682), .o(n_24775) );
in01f80 FE_OCPC1732_n_34369 ( .a(FE_OCPN1731_n_34369), .o(FE_OCPN1732_n_34369) );
in01f80 FE_OCP_RBC1369_n_20763 ( .a(FE_OCP_RBN1368_n_20763), .o(FE_OCP_RBN1369_n_20763) );
in01f80 FE_OCP_RBC2711_n_35075 ( .a(FE_OCP_RBN2710_n_35075), .o(FE_OCP_RBN2711_n_35075) );
no02f80 FE_RC_3203_0 ( .a(FE_RN_1423_0), .b(n_7580), .o(n_8676) );
in01f80 newInst_3596 ( .a(newNet_2405), .o(newNet_3596) );
na02f80 g738916 ( .a(n_41202), .b(n_41201), .o(n_41203) );
oa12f80 g751210 ( .a(n_29761), .b(n_29771), .c(n_29760), .o(n_30033) );
no02f80 g756593 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n_23874) );
na02f80 g741968 ( .a(n_38039), .b(n_38033), .o(n_38116) );
in01f80 g749145 ( .a(n_32230), .o(n_32231) );
oa22f80 FE_RC_2674_0 ( .a(n_11786), .b(n_11817), .c(n_11704), .d(n_11818), .o(n_12005) );
na02f80 g764216 ( .a(n_16488), .b(n_16511), .o(n_16602) );
in01f80 FE_OCPC960_n_3951 ( .a(FE_OCPN958_n_3951), .o(FE_OCPN960_n_3951) );
oa22f80 FE_RC_1357_0 ( .a(FE_OCP_RBN3050_n_11329), .b(n_11324), .c(n_11323), .d(n_11329), .o(n_11403) );
oa22f80 g779882 ( .a(n_44652), .b(n_1168), .c(n_44637), .d(n_1150), .o(n_1333) );
na02f80 g754866 ( .a(n_25277), .b(n_25242), .o(n_25517) );
na02f80 g749676 ( .a(n_30152), .b(n_30151), .o(n_30153) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_3_ ( .ck(newNet_3004), .d(n_966), .o(delay_add_ln22_unr2_stage2_stallmux_q_3_) );
na02f80 g751715 ( .a(n_28359), .b(n_28127), .o(n_28383) );
oa22f80 g765265 ( .a(FE_OCP_RBN3622_n_15135), .b(FE_OCP_RBN2450_n_14114), .c(FE_OCP_RBN2709_n_15135), .d(n_14274), .o(n_15523) );
in01f80 FE_RC_1282_0 ( .a(n_3031), .o(FE_RN_379_0) );
in01f80 newInst_1414 ( .a(newNet_1413), .o(newNet_1414) );
in01f80 g763364 ( .a(n_17039), .o(n_17083) );
no02f80 FE_RC_4160_0 ( .a(FE_RN_1811_0), .b(n_33034), .o(FE_RN_1812_0) );
in01f80 FE_OCP_RBC1374_n_35275 ( .a(n_35275), .o(FE_OCP_RBN1374_n_35275) );
na02f80 g769262 ( .a(n_11627), .b(FE_OCPN3188_n_11012), .o(n_11621) );
in01f80 g748094 ( .a(n_31876), .o(n_31877) );
na02f80 g742229 ( .a(n_44887), .b(n_38269), .o(n_38291) );
no02f80 g741905 ( .a(n_38075), .b(n_37979), .o(n_38338) );
in01f80 newInst_141 ( .a(newNet_140), .o(newNet_141) );
oa12f80 g750343 ( .a(n_29943), .b(n_30663), .c(n_30380), .o(n_30721) );
no02f80 g750178 ( .a(n_29793), .b(n_29792), .o(n_29794) );
in01f80 g779062 ( .a(n_2111), .o(n_2112) );
ao22s80 FE_RC_690_0 ( .a(n_39177), .b(n_39469), .c(n_39176), .d(n_39441), .o(n_39553) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_21_ ( .ck(newNet_2281), .d(n_40507), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_) );
in01f80 newInst_3269 ( .a(newNet_3268), .o(newNet_3269) );
na02f80 g755583 ( .a(n_24450), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24477) );
in01f80 FE_OCPC1389_n_9220 ( .a(n_9220), .o(FE_OCPN1389_n_9220) );
oa12f80 g754601 ( .a(n_25234), .b(n_25365), .c(n_25175), .o(n_25429) );
na02f80 g755288 ( .a(n_24971), .b(n_24915), .o(n_24986) );
in01f80 g736464 ( .a(n_43768), .o(n_43762) );
in01f80 FE_OCP_RBC1683_n_33491 ( .a(FE_OCP_RBN1682_n_33491), .o(FE_OCP_RBN1683_n_33491) );
ao22s80 g779198 ( .a(n_44811), .b(n_1809), .c(n_44812), .d(n_1810), .o(n_1887) );
in01f80 newInst_99 ( .a(newNet_61), .o(newNet_99) );
no02f80 FE_RC_2421_0 ( .a(FE_RN_957_0), .b(n_6836), .o(FE_RN_958_0) );
no02f80 g748957 ( .a(n_31155), .b(n_31133), .o(n_31265) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_1_ ( .ck(newNet_2478), .d(n_31176), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_0_ ( .ck(newNet_2888), .d(n_9474), .o(delay_add_ln22_unr8_stage4_stallmux_q_0_) );
ao12f80 g777831 ( .a(n_2922), .b(n_3236), .c(n_2977), .o(n_3255) );
no02f80 g775282 ( .a(n_5810), .b(n_4759), .o(n_5836) );
na02f80 g766648 ( .a(FE_OCP_RBN2357_n_13818), .b(FE_OCP_RBN2246_n_13017), .o(n_13862) );
in01f80 g766074 ( .a(n_14719), .o(n_14661) );
na02f80 g738082 ( .a(n_42042), .b(n_41904), .o(n_42074) );
in01f80 newInst_977 ( .a(newNet_976), .o(newNet_977) );
no02f80 g780025 ( .a(n_1256), .b(n_985), .o(n_1262) );
no02f80 g773518 ( .a(n_7468), .b(n_7467), .o(n_8303) );
na02f80 g777344 ( .a(n_3562), .b(n_3012), .o(n_3590) );
no02f80 g754693 ( .a(FE_OCP_RBN2961_n_26231), .b(n_26507), .o(n_26861) );
oa12f80 g767505 ( .a(n_12774), .b(n_13382), .c(n_12982), .o(n_13426) );
in01f80 g760752 ( .a(n_19688), .o(n_19689) );
in01f80 g739017 ( .a(n_41141), .o(n_41526) );
no02f80 g774456 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_18_), .o(n_6749) );
na02f80 g765892 ( .a(n_15092), .b(n_14968), .o(n_14970) );
oa12f80 g759137 ( .a(n_20674), .b(n_20983), .c(n_20575), .o(n_21088) );
na02f80 g745965 ( .a(n_34059), .b(n_34058), .o(n_34076) );
na02f80 g739058 ( .a(n_41131), .b(n_41130), .o(n_41132) );
no02f80 g784781 ( .a(n_44222), .b(FE_OCP_RBN2563_n_34905), .o(n_47267) );
ao12f80 g768763 ( .a(n_12096), .b(n_12095), .c(n_12094), .o(n_12223) );
in01f80 newInst_2002 ( .a(newNet_1153), .o(newNet_2002) );
oa22f80 FE_RC_1462_0 ( .a(n_27523), .b(n_27695), .c(n_27524), .d(n_27673), .o(n_27783) );
na02f80 g737766 ( .a(n_42193), .b(n_42209), .o(n_42210) );
na02f80 FE_RC_2383_0 ( .a(FE_RN_930_0), .b(n_12623), .o(FE_RN_931_0) );
oa12f80 g764855 ( .a(n_15685), .b(n_15684), .c(n_15683), .o(n_15757) );
no02f80 g743748 ( .a(n_36110), .b(n_35692), .o(n_36247) );
in01f80 g756377 ( .a(n_23948), .o(n_23889) );
no02f80 g767413 ( .a(n_13367), .b(FE_OCPN1854_n_13366), .o(n_13417) );
na02f80 g780162 ( .a(n_1170), .b(n_1148), .o(n_1149) );
no02f80 g766311 ( .a(n_14201), .b(n_14120), .o(n_14165) );
no02f80 g768533 ( .a(n_12269), .b(n_12193), .o(n_12357) );
no02f80 g763598 ( .a(n_17607), .b(n_17604), .o(n_17608) );
na02f80 FE_RC_1733_0 ( .a(n_36887), .b(n_36910), .o(FE_RN_482_0) );
na02f80 g775539 ( .a(n_5484), .b(FE_OCP_RBN2733_n_4219), .o(n_5650) );
in01f80 g769129 ( .a(n_11741), .o(n_11742) );
no02f80 g775449 ( .a(n_5531), .b(n_4759), .o(n_5544) );
in01f80 g766831 ( .a(n_14423), .o(n_14424) );
in01f80 g758013 ( .a(n_22336), .o(n_22337) );
in01f80 g770950 ( .a(n_10165), .o(n_10166) );
in01f80 g752005 ( .a(n_29098), .o(n_29099) );
na02f80 g754710 ( .a(FE_OCP_RBN2960_n_26231), .b(n_26451), .o(n_26863) );
in01f80 g761847 ( .a(n_18515), .o(n_18551) );
oa22f80 FE_RC_2192_0 ( .a(FE_RN_784_0), .b(n_14951), .c(FE_RN_785_0), .d(n_15009), .o(n_15208) );
no02f80 g741619 ( .a(n_38614), .b(n_38602), .o(n_38690) );
no02f80 g738693 ( .a(n_41537), .b(n_41255), .o(n_41560) );
in01f80 newInst_1294 ( .a(newNet_1162), .o(newNet_1294) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_2_ ( .ck(newNet_917), .d(n_27737), .o(delay_xor_ln21_unr18_stage7_stallmux_q_2_) );
in01f80 newInst_2713 ( .a(newNet_2712), .o(newNet_2713) );
in01f80 g737691 ( .a(n_42334), .o(n_42364) );
na02f80 FE_RC_2999_0 ( .a(FE_RN_1309_0), .b(FE_RN_1312_0), .o(n_6720) );
no02f80 g737067 ( .a(n_43082), .b(n_43123), .o(n_43215) );
no02f80 g738026 ( .a(n_42147), .b(n_42196), .o(n_42166) );
na02f80 g744395 ( .a(n_35501), .b(FE_OCP_DRV_N1582_n_35500), .o(n_35517) );
oa12f80 g773121 ( .a(n_7910), .b(n_8362), .c(n_7356), .o(n_8638) );
na02f80 g776210 ( .a(n_4740), .b(n_4795), .o(n_5048) );
na02f80 g745647 ( .a(n_34452), .b(n_34427), .o(n_34453) );
ao12f80 g762050 ( .a(n_47248), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_21_), .o(n_18456) );
in01f80 g774978 ( .a(n_6100), .o(n_6101) );
na02f80 g779340 ( .a(n_1657), .b(n_1656), .o(n_1698) );
na02f80 g766951 ( .a(n_14758), .b(n_14257), .o(n_14297) );
no02f80 g767288 ( .a(n_13547), .b(n_13569), .o(n_13606) );
in01f80 newInst_487 ( .a(newNet_363), .o(newNet_487) );
in01f80 g745559 ( .a(n_34558), .o(n_34559) );
in01f80 FE_OCP_RBC2875_n_5082 ( .a(n_5082), .o(FE_OCP_RBN2875_n_5082) );
in01f80 g744214 ( .a(n_36093), .o(n_36094) );
no02f80 g744269 ( .a(n_44180), .b(n_34871), .o(n_35690) );
in01f80 g772212 ( .a(n_8637), .o(n_8612) );
in01f80 g779633 ( .a(n_1504), .o(n_1505) );
in01f80 g777575 ( .a(n_3788), .o(n_3938) );
in01f80 g767381 ( .a(n_13270), .o(n_13298) );
in01f80 g761473 ( .a(n_19953), .o(n_19926) );
ao22s80 g781145 ( .a(n_206), .b(n_147), .c(n_208), .d(n_148), .o(n_387) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_4_ ( .ck(newNet_1371), .d(n_36285), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_) );
no02f80 g739208 ( .a(n_40862), .b(n_40861), .o(n_40911) );
na02f80 g770504 ( .a(n_10274), .b(n_44464), .o(n_10325) );
no02f80 g753766 ( .a(n_26519), .b(n_26219), .o(n_26520) );
in01f80 g748879 ( .a(n_32376), .o(n_32377) );
in01f80 g757515 ( .a(n_22806), .o(n_22776) );
in01f80 g746888 ( .a(n_33097), .o(n_33180) );
in01f80 g736754 ( .a(n_43274), .o(n_43275) );
ao12f80 g765223 ( .a(FE_OFN765_n_15670), .b(n_15837), .c(n_14779), .o(n_15878) );
in01f80 g764663 ( .a(n_15992), .o(n_16191) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_5_ ( .ck(newNet_883), .d(n_32334), .o(delay_xor_ln21_unr21_stage8_stallmux_q_5_) );
oa22f80 g784366 ( .a(FE_OFN775_n_46137), .b(n_5210), .c(FE_OFN805_n_46196), .d(n_5244), .o(n_46172) );
ao22s80 g773963 ( .a(n_6822), .b(n_6660), .c(FE_OCP_RBN3375_n_6822), .d(n_6661), .o(n_6934) );
no02f80 g770273 ( .a(n_10601), .b(n_10696), .o(n_10736) );
in01f80 g759525 ( .a(n_20849), .o(n_20999) );
in01f80 g746465 ( .a(n_34964), .o(n_34965) );
na02f80 g761655 ( .a(n_19492), .b(n_19491), .o(n_19493) );
in01f80 g738961 ( .a(n_41215), .o(n_41216) );
oa12f80 g772451 ( .a(n_8406), .b(n_8354), .c(n_45212), .o(n_8407) );
na02f80 g769591 ( .a(n_11375), .b(n_11374), .o(n_11376) );
in01f80 FE_RC_2874_0 ( .a(n_18716), .o(FE_RN_1241_0) );
no02f80 g746578 ( .a(n_33407), .b(n_33327), .o(n_33450) );
na02f80 g762440 ( .a(n_18049), .b(n_18048), .o(n_18109) );
ao12f80 g759742 ( .a(n_21778), .b(n_21694), .c(n_21714), .o(n_21863) );
no02f80 g760452 ( .a(n_20049), .b(n_19888), .o(n_20064) );
no02f80 g752184 ( .a(n_27939), .b(delay_add_ln22_unr17_stage7_stallmux_q_2_), .o(n_28067) );
in01f80 g777152 ( .a(n_4819), .o(n_4779) );
in01f80 g740033 ( .a(n_39984), .o(n_39985) );
in01f80 g769302 ( .a(n_11510), .o(n_11915) );
in01f80 g749854 ( .a(n_31321), .o(n_31280) );
in01f80 g737065 ( .a(n_43292), .o(n_43293) );
in01f80 g746894 ( .a(n_33199), .o(n_33153) );
in01f80 newInst_2115 ( .a(newNet_959), .o(newNet_2115) );
in01f80 g738217 ( .a(n_42065), .o(n_41988) );
in01f80 g747758 ( .a(n_32143), .o(n_32144) );
in01f80 newInst_277 ( .a(newNet_276), .o(newNet_277) );
no02f80 g761279 ( .a(n_19073), .b(n_19130), .o(n_19187) );
in01f80 FE_OCP_RBC2743_n_15319 ( .a(n_15319), .o(FE_OCP_RBN2743_n_15319) );
na02f80 g739171 ( .a(n_40869), .b(n_40795), .o(n_40914) );
no02f80 g737555 ( .a(n_42521), .b(n_42505), .o(n_42590) );
oa12f80 g744664 ( .a(n_35270), .b(n_35269), .c(n_35268), .o(n_35309) );
in01f80 g760607 ( .a(n_19816), .o(n_19839) );
oa12f80 g743780 ( .a(n_37264), .b(n_37283), .c(n_46234), .o(n_37305) );
na02f80 g777647 ( .a(n_3490), .b(n_3489), .o(n_3491) );
in01f80 g775121 ( .a(n_5968), .o(n_5969) );
no02f80 g769453 ( .a(n_11387), .b(n_11410), .o(n_11480) );
na02f80 g740832 ( .a(n_39264), .b(n_39057), .o(n_39265) );
na02f80 g756801 ( .a(n_23455), .b(n_23419), .o(n_23473) );
in01f80 g741289 ( .a(n_38940), .o(n_38976) );
in01f80 g769587 ( .a(n_11405), .o(n_11424) );
na02f80 g774014 ( .a(n_6903), .b(n_47210), .o(n_6994) );
in01f80 g763761 ( .a(n_17704), .o(n_17705) );
na02f80 g755478 ( .a(n_24649), .b(n_22393), .o(n_24803) );
na02f80 g737785 ( .a(n_42624), .b(n_42557), .o(n_42641) );
no02f80 g740925 ( .a(n_39261), .b(n_39281), .o(n_39368) );
na02f80 g746938 ( .a(n_32862), .b(n_32861), .o(n_32919) );
in01f80 g780988 ( .a(n_374), .o(n_377) );
in01f80 g776265 ( .a(n_4454), .o(n_4505) );
in01f80 g767024 ( .a(n_14347), .o(n_14294) );
in01f80 FE_OCP_RBC3530_n_13765 ( .a(FE_OCP_RBN3527_n_13765), .o(FE_OCP_RBN3530_n_13765) );
in01f80 g776994 ( .a(n_3909), .o(n_3910) );
no02f80 g770623 ( .a(n_10063), .b(n_10020), .o(n_10149) );
no02f80 g758881 ( .a(n_21330), .b(n_21365), .o(n_21366) );
in01f80 g748309 ( .a(n_31768), .o(n_31769) );
in01f80 newInst_2607 ( .a(newNet_841), .o(newNet_2607) );
in01f80 newInst_919 ( .a(newNet_918), .o(newNet_919) );
ao12f80 g762957 ( .a(n_17985), .b(n_17984), .c(n_17983), .o(n_18487) );
na02f80 FE_RC_3702_0 ( .a(FE_RN_1628_0), .b(FE_RN_1629_0), .o(FE_RN_1630_0) );
in01f80 fopt783576 ( .a(n_45204), .o(n_45203) );
na02f80 g775715 ( .a(n_5255), .b(n_4556), .o(n_5345) );
in01f80 FE_OCP_RBC3510_n_19599 ( .a(n_19599), .o(FE_OCP_RBN3510_n_19599) );
in01f80 newInst_597 ( .a(newNet_596), .o(newNet_597) );
na02f80 g749796 ( .a(n_31311), .b(n_31416), .o(n_31511) );
no03m80 g784071 ( .a(n_45808), .b(n_970), .c(n_754), .o(n_45817) );
in01f80 g736857 ( .a(n_43543), .o(n_43544) );
na02f80 g761013 ( .a(n_19301), .b(n_18032), .o(n_19351) );
in01f80 g759565 ( .a(n_20730), .o(n_20731) );
in01f80 FE_RC_1869_0 ( .a(FE_OCP_RBN3368_n_32436), .o(FE_RN_576_0) );
no02f80 g742680 ( .a(n_37398), .b(n_37875), .o(n_37414) );
in01f80 g745037 ( .a(n_35567), .o(n_34926) );
no02f80 g768339 ( .a(n_12590), .b(n_12355), .o(n_12607) );
oa12f80 g777967 ( .a(n_2871), .b(n_3063), .c(n_2800), .o(n_3064) );
no02f80 g774162 ( .a(n_6654), .b(n_4373), .o(n_6669) );
no02f80 FE_RC_2579_0 ( .a(FE_RN_1061_0), .b(FE_RN_1062_0), .o(FE_RN_1063_0) );
no02f80 g739469 ( .a(n_44769), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .o(n_40802) );
na02f80 FE_RC_1104_0 ( .a(FE_RN_329_0), .b(n_45153), .o(n_40757) );
in01f80 g768473 ( .a(n_12418), .o(n_12373) );
no02f80 FE_RC_2824_0 ( .a(FE_RN_1209_0), .b(FE_RN_1212_0), .o(n_34820) );
in01f80 g764366 ( .a(n_16369), .o(n_16370) );
in01f80 newInst_3724 ( .a(newNet_3723), .o(newNet_3724) );
in01f80 g743393 ( .a(n_37826), .o(n_37827) );
no02f80 g741481 ( .a(n_38745), .b(n_38760), .o(n_38781) );
na02f80 g773564 ( .a(n_7454), .b(n_7093), .o(n_7507) );
na02f80 g767953 ( .a(n_12841), .b(n_12810), .o(n_12842) );
no02f80 g739310 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40902) );
oa12f80 g736357 ( .a(n_342), .b(n_43835), .c(n_43918), .o(n_43865) );
in01f80 g745251 ( .a(FE_OCP_DRV_N1592_n_34327), .o(n_35598) );
no02f80 FE_RC_1695_0 ( .a(n_26016), .b(n_25614), .o(FE_RN_469_0) );
in01f80 FE_OCP_RBC1159_n_18517 ( .a(FE_OCP_RBN1158_n_18517), .o(FE_OCP_RBN1159_n_18517) );
in01f80 g765920 ( .a(n_14802), .o(n_14803) );
no02f80 g765872 ( .a(n_15210), .b(n_15209), .o(n_15211) );
na02f80 g738515 ( .a(n_41420), .b(n_41316), .o(n_41677) );
na02f80 g743787 ( .a(n_37283), .b(n_46234), .o(n_37264) );
in01f80 g764353 ( .a(n_16371), .o(n_16392) );
no02f80 g745360 ( .a(n_34487), .b(n_34511), .o(n_34539) );
na02f80 g753637 ( .a(n_26657), .b(n_26656), .o(n_26754) );
in01f80 g759328 ( .a(n_21242), .o(n_21339) );
in01f80 g759105 ( .a(n_21421), .o(n_21422) );
no02f80 g769597 ( .a(n_11320), .b(FE_OCP_RBN2845_n_10326), .o(n_11337) );
in01f80 newInst_1657 ( .a(newNet_780), .o(newNet_1657) );
in01f80 g754515 ( .a(n_25513), .o(n_25544) );
in01f80 g752687 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_13_), .o(n_28449) );
no02f80 g765924 ( .a(n_15089), .b(n_14347), .o(n_15245) );
ao12f80 g746857 ( .a(n_33098), .b(n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n_33140) );
in01f80 newInst_3561 ( .a(newNet_3560), .o(newNet_3561) );
na02f80 g769021 ( .a(n_11519), .b(n_11440), .o(n_11600) );
no02f80 g766870 ( .a(n_13976), .b(n_13937), .o(n_13977) );
in01f80 g753924 ( .a(n_26322), .o(n_26405) );
in01f80 newInst_1802 ( .a(newNet_1344), .o(newNet_1802) );
na02f80 g749026 ( .a(n_31029), .b(n_27536), .o(n_31031) );
no02f80 g758680 ( .a(n_21791), .b(FE_OCPN1532_n_21790), .o(n_21812) );
in01f80 g737172 ( .a(n_43020), .o(n_43032) );
no02f80 g775339 ( .a(n_5814), .b(n_5000), .o(n_5894) );
in01f80 g768298 ( .a(n_12565), .o(n_12566) );
in01f80 g753827 ( .a(n_26462), .o(n_26463) );
in01f80 g745638 ( .a(n_34398), .o(n_34399) );
na02f80 g763401 ( .a(FE_OCP_RBN3724_n_16975), .b(FE_OCP_RBN2918_n_16084), .o(n_17180) );
na02f80 g740056 ( .a(n_39950), .b(n_39561), .o(n_39981) );
na02f80 g770762 ( .a(FE_OCP_RBN3654_n_10100), .b(n_9111), .o(n_10414) );
in01f80 FE_OFC86_n_46137 ( .a(FE_OFN773_n_46137), .o(FE_OFN86_n_46137) );
no02f80 g750356 ( .a(n_29658), .b(n_29663), .o(n_29686) );
na02f80 g773127 ( .a(FE_OCP_RBN2229_n_7598), .b(n_7707), .o(n_7741) );
oa22f80 FE_RC_1440_0 ( .a(n_32566), .b(n_32310), .c(n_28336), .d(n_32285), .o(n_32353) );
no02f80 g777400 ( .a(n_3478), .b(n_3559), .o(n_3570) );
in01f80 newInst_1897 ( .a(newNet_1896), .o(newNet_1897) );
in01f80 FE_OCP_RBC2244_n_13017 ( .a(FE_OCP_RBN2242_n_13017), .o(FE_OCP_RBN2244_n_13017) );
ao22s80 g773728 ( .a(n_7270), .b(n_6977), .c(n_7280), .d(n_6976), .o(n_7828) );
in01f80 g772611 ( .a(n_8186), .o(n_8206) );
in01f80 g748911 ( .a(n_32457), .o(n_32409) );
na02f80 g745874 ( .a(n_35338), .b(n_35337), .o(n_35339) );
in01f80 g755409 ( .a(n_24918), .o(n_24911) );
na02f80 g781054 ( .a(sin_out_8), .b(FE_OFN3_n_43918), .o(n_335) );
oa12f80 g761511 ( .a(n_19649), .b(n_19760), .c(n_19758), .o(n_19876) );
no02f80 g752242 ( .a(n_27938), .b(n_44735), .o(n_28004) );
in01f80 FE_OCP_RBC3818_n_44061 ( .a(n_44061), .o(FE_OCP_RBN3818_n_44061) );
na02f80 g769712 ( .a(n_11202), .b(n_11224), .o(n_11301) );
no02f80 g760485 ( .a(n_19978), .b(n_20004), .o(n_20103) );
na02f80 g754301 ( .a(n_25876), .b(n_25854), .o(n_25928) );
oa12f80 g745556 ( .a(n_34383), .b(n_34286), .c(n_34313), .o(n_34929) );
na02f80 g756998 ( .a(n_23265), .b(n_23290), .o(n_23457) );
no02f80 g771541 ( .a(n_9086), .b(FE_OCPN1251_n_8210), .o(n_9135) );
na02f80 g757847 ( .a(n_22318), .b(n_21970), .o(n_22358) );
in01f80 newInst_1277 ( .a(newNet_1276), .o(newNet_1277) );
na02f80 g759129 ( .a(n_21459), .b(FE_OCP_DRV_N1596_n_21458), .o(n_21569) );
oa22f80 g784352 ( .a(FE_OFN86_n_46137), .b(n_6071), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_6105), .o(n_46158) );
in01f80 g750642 ( .a(n_29349), .o(n_29350) );
na02f80 FE_RC_2669_0 ( .a(FE_RN_1115_0), .b(n_3690), .o(FE_RN_1116_0) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_8_ ( .ck(newNet_1162), .d(n_4987), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_) );
ao12f80 g745346 ( .a(n_36055), .b(n_35956), .c(n_35633), .o(n_36113) );
in01f80 FE_OCP_RBC2475_n_8664 ( .a(FE_OCP_RBN2473_n_8664), .o(FE_OCP_RBN2475_n_8664) );
oa12f80 g748780 ( .a(n_30857), .b(n_31061), .c(n_30943), .o(n_31062) );
no02f80 g747640 ( .a(n_32151), .b(n_31787), .o(n_32195) );
oa12f80 g777946 ( .a(n_3047), .b(n_3116), .c(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(n_3161) );
in01f80 g775621 ( .a(n_5377), .o(n_5378) );
na02f80 g775435 ( .a(n_5349), .b(n_5422), .o(n_5423) );
ao12f80 g774211 ( .a(n_6924), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .o(n_7024) );
in01f80 FE_OCP_RBC3085_n_31819 ( .a(FE_OCP_RBN3084_n_31819), .o(FE_OCP_RBN3085_n_31819) );
in01f80 FE_OCP_RBC2150_n_11763 ( .a(n_11763), .o(FE_OCP_RBN2150_n_11763) );
na02f80 g773207 ( .a(n_7817), .b(n_7828), .o(n_7891) );
no02f80 g748434 ( .a(FE_OCPN1052_n_31674), .b(FE_OCPN975_n_46956), .o(n_31758) );
in01f80 FE_OCPC1752_n_29420 ( .a(FE_OCPN1751_n_29420), .o(FE_OCPN1752_n_29420) );
in01f80 newInst_537 ( .a(newNet_536), .o(newNet_537) );
no02f80 g775668 ( .a(n_5545), .b(n_5213), .o(n_5570) );
in01f80 FE_OCPC3783_n_16463 ( .a(FE_OCPN3782_n_16463), .o(FE_OCPN3783_n_16463) );
in01f80 g767625 ( .a(n_12980), .o(n_13055) );
no02f80 g754331 ( .a(n_25820), .b(n_25647), .o(n_25895) );
in01f80 g757624 ( .a(n_22718), .o(n_22679) );
no02f80 g738877 ( .a(n_41304), .b(n_41303), .o(n_41305) );
na02f80 g738462 ( .a(n_41669), .b(n_41690), .o(n_41764) );
oa22f80 g779072 ( .a(n_1974), .b(n_1779), .c(n_1975), .d(n_1778), .o(n_2515) );
in01f80 newInst_390 ( .a(newNet_389), .o(newNet_390) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_16_ ( .ck(newNet_653), .d(n_46354), .o(delay_xor_ln21_unr9_stage4_stallmux_q_16_) );
in01f80 newInst_258 ( .a(newNet_257), .o(newNet_258) );
na02f80 FE_RC_2931_0 ( .a(FE_RN_1277_0), .b(n_39812), .o(n_39866) );
in01f80 FE_OCP_RBC1162_n_24701 ( .a(n_24701), .o(FE_OCP_RBN1162_n_24701) );
in01f80 g780224 ( .a(n_1102), .o(n_1064) );
in01f80 g771872 ( .a(n_9051), .o(n_9108) );
ao12f80 g768564 ( .a(n_12266), .b(n_12265), .c(n_12264), .o(n_12325) );
in01f80 g746058 ( .a(n_34427), .o(n_34026) );
in01f80 FE_OCP_RBC2888_n_46957 ( .a(n_46957), .o(FE_OCP_RBN2888_n_46957) );
in01f80 newInst_3172 ( .a(newNet_3171), .o(newNet_3172) );
in01f80 g771103 ( .a(n_9764), .o(n_9712) );
no02f80 g744298 ( .a(n_44180), .b(n_35090), .o(n_36095) );
no02f80 g757934 ( .a(n_22080), .b(n_21960), .o(n_22113) );
in01f80 FE_OCP_RBC2701_n_4041 ( .a(n_4041), .o(FE_OCP_RBN2701_n_4041) );
in01f80 g748376 ( .a(n_31477), .o(n_31559) );
na02f80 g741051 ( .a(n_39037), .b(n_38950), .o(n_39483) );
no02f80 g740087 ( .a(n_40107), .b(n_40206), .o(n_40253) );
in01f80 fopt783041 ( .a(n_44511), .o(n_44516) );
in01f80 g767840 ( .a(n_12997), .o(n_12998) );
no02f80 g760834 ( .a(n_19556), .b(n_19501), .o(n_19557) );
na02f80 g740146 ( .a(n_39816), .b(n_39864), .o(n_39843) );
ao12f80 g748840 ( .a(n_32442), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n_32747) );
in01f80 newInst_223 ( .a(newNet_222), .o(newNet_223) );
oa12f80 g762758 ( .a(n_17540), .b(n_18156), .c(n_17633), .o(n_18237) );
in01f80 g741195 ( .a(n_38986), .o(n_39035) );
in01f80 FE_OCP_RBC3335_n_44962 ( .a(n_44962), .o(FE_OCP_RBN3335_n_44962) );
na02f80 g775734 ( .a(n_5491), .b(n_3740), .o(n_5589) );
na02f80 g774050 ( .a(n_6746), .b(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_7224) );
na02f80 g751043 ( .a(n_29997), .b(n_29945), .o(n_30479) );
ao12f80 g773933 ( .a(n_6995), .b(n_6994), .c(n_7000), .o(n_7883) );
no02f80 g770968 ( .a(n_9847), .b(n_9928), .o(n_9929) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_26_ ( .ck(newNet_802), .d(n_1303), .o(delay_xor_ln21_unr3_stage2_stallmux_q_26_) );
oa12f80 g759721 ( .a(n_21107), .b(n_21172), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21877) );
in01f80 FE_OCP_RBC3368_n_32436 ( .a(n_32436), .o(FE_OCP_RBN3368_n_32436) );
no02f80 g756029 ( .a(n_24981), .b(n_24980), .o(n_25033) );
na02f80 g746878 ( .a(n_33108), .b(n_32354), .o(n_33376) );
in01f80 g742726 ( .a(n_38279), .o(n_37453) );
in01f80 g780195 ( .a(n_1137), .o(n_1121) );
ao12f80 g746839 ( .a(n_33233), .b(FE_OCP_RBN3384_n_33108), .c(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n_33250) );
in01f80 g738835 ( .a(n_41654), .o(n_41326) );
in01f80 newInst_2844 ( .a(newNet_418), .o(newNet_2844) );
ao12f80 g777707 ( .a(n_2803), .b(n_3367), .c(n_2745), .o(n_3490) );
in01f80 newInst_1827 ( .a(newNet_1826), .o(newNet_1827) );
in01f80 FE_OCPC1857_n_22207 ( .a(n_22207), .o(FE_OCPN1857_n_22207) );
in01f80 g753638 ( .a(n_26692), .o(n_26755) );
in01f80 FE_RC_69_0 ( .a(n_18515), .o(FE_RN_19_0) );
no02f80 g777239 ( .a(n_3748), .b(n_3797), .o(n_3989) );
in01f80 fopt783158 ( .a(n_40577), .o(n_44690) );
no02f80 g755793 ( .a(n_24958), .b(n_24929), .o(n_25006) );
oa12f80 g781088 ( .a(n_253), .b(n_252), .c(n_251), .o(n_476) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_13_ ( .ck(newNet_2490), .d(n_32252), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_) );
no02f80 g754014 ( .a(n_26136), .b(n_26122), .o(n_26181) );
no02f80 g740157 ( .a(FE_OCP_RBN3722_n_39913), .b(n_40183), .o(n_40218) );
na02f80 g755491 ( .a(n_24576), .b(n_23359), .o(n_24661) );
na03f80 FE_RC_40_0 ( .a(n_6393), .b(n_6404), .c(n_6463), .o(n_6535) );
in01f80 g774342 ( .a(n_7029), .o(n_7030) );
no02f80 g763242 ( .a(n_17335), .b(n_17232), .o(n_17438) );
in01f80 g780455 ( .a(n_840), .o(n_919) );
oa22f80 g778461 ( .a(n_2694), .b(n_2124), .c(n_2614), .d(n_2125), .o(n_2782) );
na02f80 g767348 ( .a(n_13636), .b(n_13256), .o(n_13678) );
no02f80 g737941 ( .a(n_42277), .b(n_42136), .o(n_42294) );
no02f80 g777353 ( .a(n_4759), .b(n_4970), .o(n_5090) );
ao12f80 g761390 ( .a(n_19574), .b(n_19573), .c(n_19572), .o(n_19931) );
in01f80 newInst_663 ( .a(newNet_662), .o(newNet_663) );
na02f80 g768129 ( .a(n_12597), .b(n_12596), .o(n_12598) );
oa12f80 g741868 ( .a(n_38014), .b(n_38190), .c(n_38016), .o(n_38366) );
na02f80 g756584 ( .a(n_23606), .b(n_23653), .o(n_23822) );
na02f80 g777367 ( .a(n_4182), .b(n_4136), .o(n_4193) );
in01f80 g748596 ( .a(n_33146), .o(n_32746) );
no02f80 g756483 ( .a(n_23629), .b(n_23630), .o(n_23718) );
in01f80 g746913 ( .a(n_33181), .o(n_33152) );
na02f80 g751285 ( .a(n_29693), .b(n_29692), .o(n_29694) );
in01f80 FE_OCP_RBC2750_n_9629 ( .a(n_9629), .o(FE_OCP_RBN2750_n_9629) );
na02f80 g780320 ( .a(n_941), .b(FE_OFN50_n_1045), .o(n_1113) );
ao22s80 g754610 ( .a(n_26856), .b(n_26855), .c(FE_OCP_RBN2960_n_26231), .d(n_26307), .o(n_26940) );
no02f80 FE_RC_3528_0 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_9_), .b(n_23266), .o(FE_RN_1525_0) );
in01f80 g773007 ( .a(n_8046), .o(n_8550) );
na02f80 g750695 ( .a(n_29369), .b(FE_OCP_RBN3436_n_29163), .o(n_29415) );
oa12f80 g737570 ( .a(n_42238), .b(n_42240), .c(n_42237), .o(n_43031) );
no02f80 g771084 ( .a(n_9704), .b(FE_OCP_RBN2394_n_8288), .o(n_9763) );
in01f80 FE_OCP_RBC3638_n_44490 ( .a(n_44490), .o(FE_OCP_RBN3638_n_44490) );
na02f80 g775394 ( .a(n_5874), .b(n_5873), .o(n_5875) );
no02f80 g763947 ( .a(n_16567), .b(n_16466), .o(n_16589) );
no02f80 g753728 ( .a(n_26529), .b(FE_OCPN1496_n_26528), .o(n_26557) );
na02f80 g777164 ( .a(n_4862), .b(n_4732), .o(n_5593) );
no02f80 g762273 ( .a(n_18693), .b(n_18528), .o(n_19547) );
no02f80 g778986 ( .a(n_2132), .b(n_2131), .o(n_2133) );
oa12f80 g740799 ( .a(n_39131), .b(n_39440), .c(n_38981), .o(n_39441) );
in01f80 newInst_553 ( .a(newNet_55), .o(newNet_553) );
no02f80 g780835 ( .a(n_645), .b(n_508), .o(n_643) );
in01f80 g748444 ( .a(n_31754), .o(n_31755) );
no02f80 g739195 ( .a(n_40681), .b(n_45153), .o(n_40748) );
ao22s80 FE_RC_1214_0 ( .a(n_7574), .b(n_8910), .c(n_7575), .d(n_8864), .o(n_9044) );
in01f80 g747430 ( .a(n_32472), .o(n_32473) );
oa12f80 g771254 ( .a(n_9689), .b(n_9688), .c(n_9687), .o(n_9760) );
oa12f80 g770707 ( .a(n_10018), .b(n_9910), .c(n_10059), .o(n_10095) );
na02f80 g736488 ( .a(n_43676), .b(n_43164), .o(n_43719) );
in01f80 FE_OCPC1399_n_8670 ( .a(n_8670), .o(FE_OCPN1399_n_8670) );
oa12f80 g748740 ( .a(n_32504), .b(n_32503), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_32584) );
ao12f80 g738973 ( .a(n_41012), .b(n_41149), .c(n_40758), .o(n_41163) );
in01f80 newInst_2669 ( .a(newNet_2668), .o(newNet_2669) );
in01f80 newInst_964 ( .a(newNet_963), .o(newNet_964) );
ao12f80 g781196 ( .a(n_45), .b(n_162), .c(n_117), .o(n_174) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_28_ ( .ck(newNet_2925), .d(FE_OCP_RBN3134_n_6567), .o(delay_add_ln22_unr5_stage3_stallmux_q_28_) );
in01f80 newInst_2873 ( .a(newNet_2740), .o(newNet_2873) );
in01f80 g739631 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .o(n_40581) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_20_ ( .ck(newNet_2285), .d(n_40498), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_) );
in01f80 FE_OCP_RBC2434_n_14072 ( .a(n_14072), .o(FE_OCP_RBN2434_n_14072) );
no02f80 g745025 ( .a(n_45185), .b(n_34397), .o(n_34830) );
in01f80 g747735 ( .a(n_33699), .o(n_33700) );
in01f80 newInst_3227 ( .a(newNet_3226), .o(newNet_3227) );
in01f80 newInst_996 ( .a(newNet_995), .o(newNet_996) );
in01f80 FE_OCP_RBC2597_n_25181 ( .a(FE_OCP_RBN2593_n_25181), .o(FE_OCP_RBN2597_n_25181) );
no02f80 g778573 ( .a(n_2441), .b(n_2082), .o(n_2465) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_0_ ( .ck(newNet_1915), .d(n_36658), .o(delay_sub_ln22_unr24_stage9_stallmux_q_0_) );
no02f80 g768081 ( .a(FE_OCP_RBN3414_n_12739), .b(n_12720), .o(n_12982) );
no02f80 g762689 ( .a(FE_OCP_RBN2142_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_12_), .o(n_18052) );
in01f80 g749014 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_), .o(n_32375) );
na02f80 g740532 ( .a(n_39668), .b(n_45530), .o(n_39674) );
ao22s80 g763162 ( .a(n_17394), .b(FE_OCP_RBN3211_n_44365), .c(n_45450), .d(delay_xor_ln22_unr12_stage5_stallmux_q_6_), .o(n_17581) );
in01f80 newInst_2795 ( .a(newNet_1881), .o(newNet_2795) );
na02f80 g746478 ( .a(n_34721), .b(n_34740), .o(n_34759) );
in01f80 newInst_403 ( .a(newNet_402), .o(newNet_403) );
na02f80 g766604 ( .a(n_13924), .b(n_13442), .o(n_13921) );
na02f80 g754848 ( .a(n_25506), .b(n_25973), .o(n_25593) );
no02f80 g738225 ( .a(n_41924), .b(n_41957), .o(n_41958) );
no02f80 g773157 ( .a(n_7612), .b(n_8135), .o(n_7646) );
oa12f80 g750969 ( .a(n_30097), .b(n_30164), .c(n_30166), .o(n_30183) );
in01f80 g776996 ( .a(n_4145), .o(n_4146) );
in01f80 newInst_1018 ( .a(newNet_1017), .o(newNet_1018) );
in01f80 newInst_585 ( .a(newNet_584), .o(newNet_585) );
in01f80 newInst_3644 ( .a(newNet_3643), .o(newNet_3644) );
no02f80 g762882 ( .a(n_17839), .b(n_17838), .o(n_17840) );
na02f80 FE_RC_3949_0 ( .a(n_32878), .b(n_33113), .o(FE_RN_1708_0) );
no02f80 g780009 ( .a(n_1269), .b(n_1026), .o(n_1282) );
na02f80 g738923 ( .a(n_41191), .b(n_40890), .o(n_41200) );
na02f80 FE_RC_2745_0 ( .a(n_12474), .b(FE_RN_1165_0), .o(n_12497) );
oa22f80 FE_RC_986_0 ( .a(n_24350), .b(n_27783), .c(n_27845), .d(n_27756), .o(n_27844) );
oa22f80 FE_RC_1274_0 ( .a(n_3029), .b(n_3807), .c(n_3615), .d(FE_OCP_RBN2607_n_3807), .o(n_3963) );
na02f80 g737698 ( .a(n_42203), .b(n_42211), .o(n_42254) );
in01f80 g761274 ( .a(n_19984), .o(n_19985) );
na02f80 g753467 ( .a(n_26878), .b(n_26917), .o(n_27019) );
ao12f80 g760559 ( .a(n_19940), .b(n_19939), .c(n_19938), .o(n_20018) );
ao12f80 g751434 ( .a(FE_OCP_RBN2192_n_28597), .b(n_28698), .c(n_27807), .o(n_28744) );
oa22f80 g762936 ( .a(n_17460), .b(n_17584), .c(n_17456), .d(n_16339), .o(n_17567) );
in01f80 g757064 ( .a(n_24110), .o(n_23830) );
no02f80 g750278 ( .a(n_29752), .b(n_28583), .o(n_29848) );
na02f80 g739235 ( .a(n_40842), .b(n_40885), .o(n_41201) );
na02f80 g749200 ( .a(n_30763), .b(n_30385), .o(n_30808) );
ao12f80 g771155 ( .a(n_9446), .b(n_9639), .c(n_9447), .o(n_9831) );
no02f80 g750482 ( .a(n_29508), .b(n_29486), .o(n_29568) );
no02f80 g767988 ( .a(n_13200), .b(n_13197), .o(n_13544) );
in01f80 newInst_1664 ( .a(newNet_1663), .o(newNet_1664) );
na02f80 g779845 ( .a(FE_OCP_RBN3247_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n_1379) );
in01f80 g750217 ( .a(n_29869), .o(n_29896) );
in01f80 g748972 ( .a(n_31153), .o(n_31154) );
ao22s80 g740818 ( .a(n_39376), .b(n_39151), .c(n_39440), .d(n_39152), .o(n_39945) );
na02f80 g777805 ( .a(n_3222), .b(n_3245), .o(n_3246) );
no02f80 g755431 ( .a(n_24657), .b(n_24310), .o(n_24728) );
ao12f80 FE_RC_1763_0 ( .a(FE_RN_503_0), .b(FE_RN_504_0), .c(n_12535), .o(n_12623) );
na02f80 g738597 ( .a(n_41608), .b(n_41324), .o(n_41661) );
in01f80 newInst_2030 ( .a(newNet_2029), .o(newNet_2030) );
in01f80 g745260 ( .a(n_34591), .o(n_34592) );
no02f80 g762037 ( .a(n_19014), .b(n_18280), .o(n_18323) );
ao12f80 g772057 ( .a(n_7568), .b(n_8621), .c(n_7581), .o(n_8747) );
oa12f80 g768443 ( .a(n_12379), .b(n_12378), .c(n_12377), .o(n_13434) );
in01f80 FE_OCP_RBC3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
na02f80 g775977 ( .a(n_5253), .b(n_47019), .o(n_5394) );
na02f80 g779083 ( .a(n_2034), .b(n_1173), .o(n_2084) );
na02f80 g776582 ( .a(n_4573), .b(n_4572), .o(n_4574) );
in01f80 newInst_3408 ( .a(newNet_204), .o(newNet_3408) );
oa12f80 g745779 ( .a(n_35374), .b(n_35373), .c(n_35372), .o(n_35845) );
in01f80 g771232 ( .a(n_9838), .o(n_9839) );
na02f80 g754236 ( .a(n_25955), .b(n_25747), .o(n_26013) );
in01f80 g779743 ( .a(n_1751), .o(n_1752) );
oa12f80 g767082 ( .a(n_13287), .b(n_13699), .c(n_13378), .o(n_13825) );
in01f80 g762049 ( .a(n_18456), .o(n_18457) );
in01f80 FE_RC_2131_0 ( .a(n_23271), .o(FE_RN_744_0) );
in01f80 g757952 ( .a(n_22313), .o(n_22349) );
oa22f80 g784344 ( .a(FE_OFN86_n_46137), .b(n_6137), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_6146), .o(n_46150) );
in01f80 g776616 ( .a(n_4313), .o(n_4314) );
na02f80 g763535 ( .a(FE_OCP_RBN1208_n_16814), .b(n_16940), .o(n_16976) );
oa22f80 g770656 ( .a(n_10068), .b(n_9987), .c(FE_OCP_RBN2824_n_10068), .d(n_10047), .o(n_10326) );
in01f80 FE_OCP_RBC2915_n_42947 ( .a(n_42947), .o(FE_OCP_RBN2915_n_42947) );
na02f80 g740255 ( .a(n_39994), .b(n_39967), .o(n_39968) );
in01f80 newInst_504 ( .a(newNet_160), .o(newNet_504) );
na02f80 g740398 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39965), .o(n_40269) );
na02f80 g775593 ( .a(n_5639), .b(n_5710), .o(n_5725) );
na02f80 g736770 ( .a(n_43521), .b(n_43307), .o(n_43560) );
in01f80 g747794 ( .a(n_33653), .o(n_33599) );
no02f80 g763904 ( .a(n_16617), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17104) );
no02f80 g739446 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n_40849) );
no02f80 g771938 ( .a(n_8895), .b(n_8833), .o(n_8926) );
in01f80 g764067 ( .a(n_17093), .o(n_17423) );
na02f80 g772695 ( .a(n_8162), .b(FE_OCP_RBN2399_FE_RN_347_0), .o(n_8219) );
oa12f80 g748641 ( .a(n_32393), .b(n_32610), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_32611) );
in01f80 g764013 ( .a(n_19418), .o(n_19645) );
na02f80 g760957 ( .a(n_19328), .b(n_18936), .o(n_19357) );
in01f80 g764704 ( .a(n_15984), .o(n_15985) );
ao22s80 g736421 ( .a(n_43729), .b(n_43550), .c(n_43728), .d(n_43549), .o(n_43771) );
no02f80 FE_RC_3146_0 ( .a(FE_RN_1396_0), .b(n_27087), .o(n_27150) );
no02f80 g756940 ( .a(n_23697), .b(n_23905), .o(n_24667) );
in01f80 fopt783161 ( .a(n_44695), .o(n_44696) );
in01f80 g763763 ( .a(n_17702), .o(n_17703) );
no02f80 g755087 ( .a(n_25688), .b(n_25195), .o(n_25800) );
in01f80 g753151 ( .a(n_27486), .o(n_27487) );
in01f80 FE_OCPC1411_n_21007 ( .a(n_21007), .o(FE_OCPN1411_n_21007) );
in01f80 g751279 ( .a(n_29993), .o(n_29756) );
na02f80 FE_RC_2196_0 ( .a(FE_OCPN1522_n_26054), .b(n_26055), .o(FE_RN_788_0) );
na02f80 g771357 ( .a(FE_OCP_RBN2521_n_8951), .b(FE_OCP_RBN3476_n_7886), .o(n_9048) );
na02f80 g758104 ( .a(n_44268), .b(FE_OCP_RBN1337_n_20941), .o(n_22261) );
na02f80 g736718 ( .a(n_43142), .b(n_43230), .o(n_43232) );
na02f80 g763154 ( .a(n_17477), .b(n_17400), .o(n_17544) );
no02f80 g738701 ( .a(FE_OCPN948_n_41382), .b(n_41494), .o(n_41879) );
in01f80 FE_OCP_RBC3498_n_8187 ( .a(n_8187), .o(FE_OCP_RBN3498_n_8187) );
oa12f80 g782643 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36950), .c(n_36992), .o(n_44037) );
no02f80 g751940 ( .a(n_28149), .b(n_28010), .o(n_28191) );
no02f80 g741946 ( .a(n_38015), .b(n_38062), .o(n_38122) );
in01f80 g766047 ( .a(n_45520), .o(n_14712) );
no02f80 g777329 ( .a(n_4675), .b(n_3501), .o(n_4901) );
in01f80 newInst_3234 ( .a(newNet_3233), .o(newNet_3234) );
ao12f80 g761351 ( .a(n_18478), .b(n_18868), .c(n_18516), .o(n_18952) );
in01f80 g740947 ( .a(n_39114), .o(n_39087) );
na02f80 g768392 ( .a(n_12528), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_), .o(n_12564) );
in01f80 newInst_2732 ( .a(newNet_358), .o(newNet_2732) );
no02f80 g768284 ( .a(n_12538), .b(n_12537), .o(n_12558) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_5_ ( .ck(newNet_2438), .d(FE_OCPUNCON1808_n_31435), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_) );
no02f80 g784601 ( .a(n_11089), .b(FE_OCP_RBN3643_n_44490), .o(n_46424) );
in01f80 g745317 ( .a(n_36167), .o(n_36168) );
ao12f80 g759821 ( .a(FE_OCP_RBN3678_n_21051), .b(n_21626), .c(n_21625), .o(n_21779) );
ao22s80 FE_RC_4109_0 ( .a(n_32099), .b(n_47205), .c(n_32100), .d(n_32279), .o(n_32394) );
no02f80 g761285 ( .a(n_18982), .b(n_18547), .o(n_19009) );
oa12f80 g737203 ( .a(n_42656), .b(n_42975), .c(n_42606), .o(n_42985) );
in01f80 FE_RC_914_0 ( .a(n_27246), .o(FE_RN_270_0) );
in01f80 g775482 ( .a(n_5841), .o(n_5795) );
no02f80 g778113 ( .a(n_2820), .b(n_2209), .o(n_2914) );
no03m80 g767725 ( .a(n_13111), .b(n_13208), .c(n_13197), .o(n_13209) );
in01f80 g769357 ( .a(n_11838), .o(n_11897) );
in01f80 g763876 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_13_), .o(n_18048) );
oa12f80 g774251 ( .a(n_6585), .b(n_6664), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n_6769) );
no02f80 g773145 ( .a(n_7743), .b(n_7794), .o(n_7922) );
na02f80 g756242 ( .a(n_24770), .b(n_24769), .o(n_24771) );
oa12f80 g751342 ( .a(n_28404), .b(n_28611), .c(n_28355), .o(n_28684) );
in01f80 g766499 ( .a(n_14144), .o(n_14145) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_3_ ( .ck(newNet_858), .d(n_40597), .o(delay_xor_ln21_unr28_stage10_stallmux_q_3_) );
in01f80 g742393 ( .a(n_37767), .o(n_37768) );
in01f80 FE_RC_2404_0 ( .a(FE_RN_947_0), .o(n_47210) );
na02f80 g765048 ( .a(n_15463), .b(n_15462), .o(n_15497) );
no02f80 g743647 ( .a(n_44831), .b(n_36071), .o(n_36467) );
no02f80 g765640 ( .a(n_14981), .b(FE_OCP_RBN2758_FE_RN_722_0), .o(n_15045) );
no02f80 g738600 ( .a(n_41422), .b(n_41421), .o(n_41423) );
no02f80 g780775 ( .a(n_540), .b(n_539), .o(n_541) );
in01f80 newInst_122 ( .a(newNet_83), .o(newNet_122) );
na02f80 g756002 ( .a(FE_OCP_RBN2525_n_24902), .b(n_24957), .o(n_25089) );
in01f80 FE_RC_3317_0 ( .a(n_17868), .o(FE_RN_1460_0) );
no02f80 FE_RC_2355_0 ( .a(n_1673), .b(FE_RN_907_0), .o(FE_RN_908_0) );
no02f80 g779540 ( .a(FE_OCP_RBN3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_2_), .o(n_1397) );
in01f80 g776315 ( .a(n_4507), .o(n_4508) );
in01f80 g759494 ( .a(n_21054), .o(n_21206) );
in01f80 newInst_753 ( .a(newNet_752), .o(newNet_753) );
no02f80 g765300 ( .a(n_15709), .b(n_15717), .o(n_16505) );
na02f80 g755031 ( .a(n_25127), .b(n_25126), .o(n_25241) );
no02f80 g737475 ( .a(n_42603), .b(n_42602), .o(n_42604) );
na02f80 g775721 ( .a(n_5159), .b(n_5204), .o(n_5212) );
na02f80 FE_RC_1649_0 ( .a(FE_OCP_RBN1379_n_20732), .b(FE_RN_460_0), .o(FE_RN_461_0) );
ao12f80 g779517 ( .a(n_1519), .b(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .o(n_1567) );
in01f80 FE_OCP_RBC2331_n_29353 ( .a(n_29353), .o(FE_OCP_RBN2331_n_29353) );
in01f80 newInst_1097 ( .a(newNet_1096), .o(newNet_1097) );
no02f80 g767063 ( .a(n_14758), .b(n_14107), .o(n_14205) );
in01f80 FE_OCP_DRV_C1556_n_19384 ( .a(FE_OCP_DRV_N1555_n_19384), .o(FE_OCP_DRV_N1556_n_19384) );
no02f80 FE_RC_1364_0 ( .a(FE_RN_407_0), .b(n_5449), .o(n_47001) );
in01f80 g755339 ( .a(n_24877), .o(n_24938) );
na02f80 g757404 ( .a(n_23400), .b(n_23382), .o(n_23383) );
in01f80 g766540 ( .a(n_13997), .o(n_13998) );
no02f80 g750840 ( .a(n_29159), .b(n_29180), .o(n_29313) );
ao22s80 FE_RC_222_0 ( .a(n_12600), .b(n_13175), .c(n_12599), .d(n_13176), .o(n_13335) );
in01f80 FE_OCPC1038_n_28318 ( .a(FE_OCPN1037_n_28318), .o(FE_OCPN1038_n_28318) );
oa12f80 g770191 ( .a(n_10818), .b(n_10817), .c(n_10816), .o(n_10868) );
no02f80 g766803 ( .a(n_13940), .b(n_13865), .o(n_14085) );
in01f80 FE_RC_4237_0 ( .a(FE_OCPN3175_n_31125), .o(FE_RN_1861_0) );
na02f80 g773966 ( .a(n_6937), .b(n_6932), .o(n_6933) );
no02f80 FE_RC_2712_0 ( .a(n_12547), .b(FE_RN_1142_0), .o(FE_RN_1143_0) );
ao12f80 g743178 ( .a(n_36907), .b(n_36908), .c(n_36906), .o(n_37744) );
in01f80 drc784099 ( .a(n_45843), .o(n_45844) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_1_ ( .ck(newNet_892), .d(n_32304), .o(delay_xor_ln21_unr21_stage8_stallmux_q_1_) );
na02f80 g745393 ( .a(n_34568), .b(n_34627), .o(n_34747) );
na02f80 g765273 ( .a(n_15116), .b(n_14758), .o(n_15118) );
in01f80 g756073 ( .a(n_24305), .o(n_24419) );
in01f80 FE_OCP_RBC3453_FE_OCPN1240_n_7721 ( .a(FE_OCPN1240_n_7721), .o(FE_OCP_RBN3453_FE_OCPN1240_n_7721) );
oa22f80 FE_RC_384_0 ( .a(n_958), .b(n_44659), .c(n_918), .d(n_44637), .o(n_1307) );
in01f80 g760422 ( .a(n_20162), .o(n_20163) );
no02f80 g753246 ( .a(n_27098), .b(n_25599), .o(n_27183) );
oa12f80 g769951 ( .a(n_10734), .b(n_10767), .c(n_10278), .o(n_10880) );
in01f80 g760036 ( .a(FE_OCP_RBN3678_n_21051), .o(n_21374) );
na02f80 g776647 ( .a(n_47009), .b(FE_OCP_RBN2465_n_4336), .o(n_4484) );
na02f80 g750688 ( .a(n_29233), .b(n_29143), .o(n_29278) );
in01f80 FE_OCP_RBC3209_n_44365 ( .a(FE_OCP_RBN3210_n_44365), .o(FE_OCP_RBN3209_n_44365) );
in01f80 FE_OCPC1524_n_45072 ( .a(FE_OCPN1523_n_45072), .o(FE_OCPN1524_n_45072) );
na02f80 g763003 ( .a(n_17579), .b(n_17618), .o(n_17671) );
oa12f80 g737861 ( .a(n_42413), .b(n_42547), .c(n_42321), .o(n_42616) );
na02f80 g746241 ( .a(n_33568), .b(n_33218), .o(n_33646) );
na02f80 g739457 ( .a(n_40663), .b(delay_add_ln22_unr27_stage10_stallmux_q_1_), .o(n_40669) );
na02f80 g763611 ( .a(n_16791), .b(FE_OCP_RBN2761_n_15200), .o(n_16879) );
na02f80 g780516 ( .a(n_1052), .b(n_761), .o(n_1054) );
oa12f80 g775303 ( .a(n_5886), .b(n_5825), .c(n_5763), .o(n_5919) );
in01f80 g774492 ( .a(n_6696), .o(n_6697) );
ao12f80 g757967 ( .a(n_23181), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_25_), .o(n_23548) );
na02f80 g736890 ( .a(n_43492), .b(n_43530), .o(n_43591) );
no02f80 g764190 ( .a(n_16444), .b(n_16434), .o(n_16496) );
no02f80 g741262 ( .a(FE_OCP_RBN2550_n_44944), .b(n_38405), .o(n_39199) );
na02f80 g766168 ( .a(n_14498), .b(FE_OCP_RBN3529_n_13765), .o(n_14576) );
na02f80 g762738 ( .a(n_17824), .b(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_17921) );
in01f80 g773992 ( .a(n_6914), .o(n_6915) );
in01f80 newInst_1682 ( .a(newNet_1681), .o(newNet_1682) );
ao12f80 g774157 ( .a(n_6753), .b(n_6668), .c(n_6676), .o(n_6754) );
in01f80 g750346 ( .a(n_29674), .o(n_29720) );
oa22f80 FE_RC_293_0 ( .a(n_20419), .b(FE_OFN751_n_45003), .c(n_45065), .d(n_20420), .o(n_20549) );
in01f80 FE_OCP_RBC3851_n_20848 ( .a(n_20848), .o(FE_OCP_RBN3851_n_20848) );
in01f80 newInst_3429 ( .a(newNet_3428), .o(newNet_3429) );
na02f80 g769081 ( .a(n_11568), .b(n_11357), .o(n_11569) );
in01f80 FE_OCP_RBC1186_n_14823 ( .a(n_14823), .o(FE_OCP_RBN1186_n_14823) );
in01f80 g778667 ( .a(n_2592), .o(n_2593) );
no02f80 g769836 ( .a(n_11128), .b(FE_OCP_RBN2769_n_9892), .o(n_11166) );
in01f80 g756739 ( .a(n_23542), .o(n_23543) );
no02f80 g759537 ( .a(n_20806), .b(n_20818), .o(n_20907) );
in01f80 g741217 ( .a(n_39269), .o(n_39270) );
ao12f80 g760385 ( .a(n_20702), .b(n_20701), .c(n_20700), .o(n_21591) );
oa12f80 g749563 ( .a(n_30487), .b(n_30486), .c(n_30485), .o(n_30573) );
no02f80 g741115 ( .a(n_38957), .b(n_38925), .o(n_38926) );
in01f80 FE_OCP_RBC1187_n_14823 ( .a(FE_OCP_RBN1186_n_14823), .o(FE_OCP_RBN1187_n_14823) );
na02f80 g763340 ( .a(n_17182), .b(n_17221), .o(n_17378) );
no02f80 g780592 ( .a(n_779), .b(n_867), .o(n_925) );
na02f80 g779331 ( .a(n_1634), .b(n_1662), .o(n_1671) );
in01f80 newInst_2331 ( .a(newNet_2330), .o(newNet_2331) );
in01f80 g772347 ( .a(n_8409), .o(n_8434) );
no02f80 g748662 ( .a(n_31166), .b(n_31162), .o(n_31308) );
no02f80 g760340 ( .a(n_20172), .b(n_20153), .o(n_20249) );
no02f80 g775292 ( .a(n_5610), .b(n_4875), .o(n_5670) );
in01f80 g775956 ( .a(n_5065), .o(n_5066) );
in01f80 g771142 ( .a(n_9578), .o(n_9674) );
in01f80 newInst_946 ( .a(newNet_945), .o(newNet_946) );
in01f80 g741301 ( .a(n_38853), .o(n_38876) );
in01f80 newInst_1175 ( .a(newNet_1174), .o(newNet_1175) );
in01f80 g772277 ( .a(n_8523), .o(n_8524) );
in01f80 g756043 ( .a(n_25081), .o(n_25052) );
in01f80 g778777 ( .a(n_2235), .o(n_2215) );
in01f80 g756032 ( .a(n_25029), .o(n_25088) );
in01f80 g768525 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_29_), .o(n_13086) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_18_ ( .ck(newNet_3631), .d(n_46974), .o(delay_add_ln22_unr11_stage5_stallmux_q_18_) );
na02f80 g784597 ( .a(n_10465), .b(FE_OCP_RBN3560_n_8809), .o(n_46420) );
no02f80 g767263 ( .a(n_13512), .b(n_13488), .o(n_13591) );
no02f80 g776333 ( .a(n_4918), .b(n_4774), .o(n_5053) );
na02f80 g739089 ( .a(n_41108), .b(n_41094), .o(n_41095) );
na02f80 g739561 ( .a(n_40633), .b(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n_40634) );
no02f80 g756457 ( .a(n_23632), .b(n_23664), .o(n_23665) );
in01f80 FE_OCP_DRV_C1571_n_29860 ( .a(n_29860), .o(FE_OCP_DRV_N1571_n_29860) );
oa12f80 g752019 ( .a(n_28100), .b(n_28099), .c(n_28098), .o(n_29155) );
ao12f80 g784800 ( .a(n_3150), .b(n_3149), .c(n_2983), .o(n_47341) );
ao22s80 FE_RC_3324_0 ( .a(n_23689), .b(n_24072), .c(n_23690), .d(n_24043), .o(n_24102) );
in01f80 FE_OCP_RBC3031_n_39942 ( .a(FE_OCP_RBN3030_n_39942), .o(FE_OCP_RBN3031_n_39942) );
in01f80 FE_RC_2363_0 ( .a(n_1748), .o(FE_RN_914_0) );
in01f80 g736959 ( .a(n_43306), .o(n_43351) );
in01f80 FE_OCP_RBC1139_n_25816 ( .a(n_25816), .o(FE_OCP_RBN1139_n_25816) );
in01f80 FE_OCP_RBC2292_n_2438 ( .a(FE_OCP_RBN2290_n_2438), .o(FE_OCP_RBN2292_n_2438) );
na02f80 g744222 ( .a(n_36183), .b(n_36138), .o(n_36289) );
in01f80 g769930 ( .a(n_11076), .o(n_11104) );
no02f80 g781136 ( .a(n_221), .b(n_264), .o(n_227) );
na02f80 g742305 ( .a(n_37837), .b(n_37836), .o(n_37842) );
na02f80 g742121 ( .a(n_38179), .b(n_38199), .o(n_38200) );
in01f80 g776815 ( .a(n_4190), .o(n_4191) );
in01f80 newInst_3358 ( .a(newNet_3357), .o(newNet_3358) );
oa12f80 g778411 ( .a(n_2429), .b(n_2428), .c(n_2427), .o(n_2664) );
no02f80 g756895 ( .a(n_23238), .b(n_23312), .o(n_23377) );
in01f80 g737083 ( .a(n_43162), .o(n_43197) );
oa22f80 g751522 ( .a(FE_OCP_RBN3407_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_29_), .c(FE_OCP_RBN2216_FE_OCPN950_n_28595), .d(n_28795), .o(n_28820) );
in01f80 g760145 ( .a(n_20570), .o(n_20571) );
no02f80 g770372 ( .a(n_10635), .b(n_10678), .o(n_10713) );
in01f80 newInst_1921 ( .a(newNet_1508), .o(newNet_1921) );
no02f80 g754019 ( .a(n_26156), .b(n_26179), .o(n_26208) );
na02f80 g756777 ( .a(n_23424), .b(delay_add_ln22_unr14_stage6_stallmux_q_12_), .o(n_23479) );
na02f80 g741636 ( .a(n_38623), .b(n_38597), .o(n_38635) );
in01f80 FE_OCP_RBC2556_n_44576 ( .a(FE_OCP_RBN3548_n_44575), .o(FE_OCP_RBN2556_n_44576) );
in01f80 FE_OCP_RBC1337_n_20941 ( .a(FE_OCP_RBN1336_n_20941), .o(FE_OCP_RBN1337_n_20941) );
in01f80 newInst_3335 ( .a(newNet_3334), .o(newNet_3335) );
in01f80 FE_RC_3385_0 ( .a(FE_RN_1468_0), .o(n_13144) );
in01f80 g771794 ( .a(n_9125), .o(n_9126) );
na02f80 g768312 ( .a(n_12530), .b(delay_add_ln22_unr8_stage4_stallmux_q_15_), .o(n_12563) );
na02f80 g745321 ( .a(n_35717), .b(n_35765), .o(n_35766) );
na02f80 g750600 ( .a(n_30394), .b(n_29936), .o(n_30441) );
na02f80 g736705 ( .a(n_43182), .b(FE_OCPN912_n_43022), .o(n_43284) );
na02f80 g758178 ( .a(n_22405), .b(n_22328), .o(n_22460) );
na02f80 FE_RC_3011_0 ( .a(FE_OCP_RBN2450_n_14114), .b(FE_OCP_RBN3622_n_15135), .o(FE_RN_1319_0) );
in01f80 g770166 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_), .o(n_11784) );
na02f80 g770724 ( .a(n_10376), .b(n_10414), .o(n_10521) );
in01f80 g774085 ( .a(n_6847), .o(n_6848) );
in01f80 newInst_1421 ( .a(newNet_1420), .o(newNet_1421) );
na02f80 g778260 ( .a(n_2615), .b(n_2587), .o(n_2588) );
oa22f80 FE_RC_26_0 ( .a(n_5095), .b(n_5561), .c(n_5096), .d(n_5562), .o(n_5693) );
no02f80 g737432 ( .a(n_42672), .b(n_42574), .o(n_42707) );
in01f80 g744967 ( .a(n_34934), .o(n_35905) );
na02f80 g778319 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_31_), .o(n_2901) );
in01f80 g778466 ( .a(n_2601), .o(n_2602) );
no02f80 g747339 ( .a(n_32600), .b(n_32438), .o(n_32551) );
no02f80 g759543 ( .a(n_20790), .b(n_44144), .o(n_20906) );
na02f80 g754920 ( .a(FE_OCP_RBN2597_n_25181), .b(n_25386), .o(n_25388) );
in01f80 newInst_292 ( .a(newNet_291), .o(newNet_292) );
ao12f80 g753588 ( .a(n_26596), .b(n_26539), .c(n_23590), .o(n_26670) );
na02f80 g741839 ( .a(n_38438), .b(n_38437), .o(n_38439) );
no02f80 g770754 ( .a(n_9819), .b(FE_OCP_RBN2478_n_8599), .o(n_9896) );
in01f80 g775023 ( .a(n_6248), .o(n_6206) );
no02f80 g748293 ( .a(n_31554), .b(n_31601), .o(n_31685) );
oa22f80 g779899 ( .a(n_44652), .b(FE_OFN794_n_45813), .c(n_44623), .d(n_1203), .o(n_1325) );
no02f80 g764403 ( .a(n_16125), .b(n_16162), .o(n_16328) );
in01f80 g753073 ( .a(n_27923), .o(n_27765) );
in01f80 newInst_1251 ( .a(newNet_1250), .o(newNet_1251) );
oa12f80 g736442 ( .a(n_43414), .b(n_43716), .c(n_43214), .o(n_43779) );
in01f80 g743630 ( .a(n_36482), .o(n_36501) );
in01f80 newInst_3592 ( .a(newNet_3591), .o(newNet_3592) );
in01f80 g752449 ( .a(n_27739), .o(n_27730) );
no02f80 g773752 ( .a(n_7279), .b(n_7260), .o(n_8174) );
in01f80 g776456 ( .a(n_4673), .o(n_4674) );
na02f80 g760123 ( .a(n_20334), .b(FE_OCP_RBN3610_FE_OCPN1797_n_20333), .o(n_20371) );
na02f80 g771456 ( .a(n_9526), .b(n_9525), .o(n_9560) );
oa12f80 g772564 ( .a(n_8360), .b(n_8359), .c(n_8358), .o(n_8426) );
in01f80 g752315 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_27_), .o(n_27860) );
na02f80 FE_RC_3161_0 ( .a(FE_OCPN1864_n_26171), .b(n_27222), .o(FE_RN_1401_0) );
oa12f80 g742868 ( .a(n_36936), .b(n_37187), .c(n_36923), .o(n_37212) );
na02f80 g781044 ( .a(sin_out_20), .b(FE_OFN3_n_43918), .o(n_307) );
na02f80 g760683 ( .a(n_19636), .b(n_19131), .o(n_19706) );
in01f80 fopt783664 ( .a(n_23044), .o(n_45312) );
in01f80 g778815 ( .a(n_3029), .o(n_3615) );
na02f80 g770411 ( .a(n_10677), .b(n_10598), .o(n_10682) );
in01f80 g767668 ( .a(n_13391), .o(n_13392) );
na02f80 g758293 ( .a(n_22288), .b(n_20649), .o(n_22409) );
no02f80 g763689 ( .a(n_16762), .b(n_16707), .o(n_16785) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_2_ ( .ck(newNet_220), .d(n_46148), .o(delay_xor_ln22_unr6_stage3_stallmux_q_2_) );
na02f80 FE_RC_902_0 ( .a(FE_RN_264_0), .b(FE_RN_265_0), .o(FE_RN_266_0) );
na02f80 g776920 ( .a(n_3979), .b(n_3849), .o(n_4010) );
in01f80 g738755 ( .a(n_41598), .o(n_41599) );
in01f80 g761204 ( .a(n_19105), .o(n_19106) );
no02f80 g753406 ( .a(n_27613), .b(n_26833), .o(n_27657) );
no02f80 g771681 ( .a(n_10073), .b(n_44516), .o(n_10124) );
na02f80 g769914 ( .a(n_10916), .b(n_44463), .o(n_10967) );
oa22f80 FE_RC_1664_0 ( .a(n_40304), .b(n_40561), .c(n_40305), .d(FE_OCP_RBN3104_n_40561), .o(n_40592) );
na02f80 g751352 ( .a(n_29036), .b(n_28647), .o(n_28774) );
na02f80 g754152 ( .a(n_25938), .b(n_23254), .o(n_25976) );
oa12f80 g770600 ( .a(n_10426), .b(n_10425), .c(n_10424), .o(n_10490) );
no02f80 g769318 ( .a(FE_OCPN858_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .o(n_11972) );
in01f80 g766210 ( .a(n_14625), .o(n_14626) );
no02f80 g778269 ( .a(n_2575), .b(n_2574), .o(n_2576) );
no02f80 g765946 ( .a(n_14721), .b(n_14581), .o(n_14753) );
in01f80 g738044 ( .a(n_42151), .o(n_42160) );
na02f80 g737669 ( .a(n_42392), .b(n_42562), .o(n_42663) );
in01f80 g738541 ( .a(n_41784), .o(n_41785) );
no02f80 g761521 ( .a(n_18801), .b(n_18760), .o(n_18899) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_14_ ( .ck(newNet_2583), .d(n_27364), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_) );
na02f80 g769988 ( .a(n_10988), .b(n_10975), .o(n_11058) );
na02f80 g759625 ( .a(n_20597), .b(n_20294), .o(n_20618) );
no02f80 g740662 ( .a(n_39481), .b(n_39207), .o(n_39498) );
ao12f80 g754830 ( .a(n_25679), .b(n_25977), .c(n_25741), .o(n_26005) );
na02f80 g766375 ( .a(n_14269), .b(n_14266), .o(n_14361) );
in01f80 newInst_628 ( .a(newNet_627), .o(newNet_628) );
in01f80 g778543 ( .a(n_2332), .o(n_2397) );
na02f80 g758945 ( .a(n_21471), .b(n_21470), .o(n_21472) );
na02f80 g742096 ( .a(FE_OCP_RBN3452_n_37945), .b(n_37574), .o(n_38163) );
na02f80 g756361 ( .a(n_24498), .b(n_23817), .o(n_24560) );
na02f80 g736835 ( .a(n_43125), .b(n_46939), .o(n_43138) );
in01f80 newInst_1706 ( .a(newNet_1705), .o(newNet_1706) );
na02f80 g778004 ( .a(n_3001), .b(n_2232), .o(n_3092) );
in01f80 FE_OCP_RBC1690_n_29491 ( .a(n_29491), .o(FE_OCP_RBN1690_n_29491) );
no02f80 g741991 ( .a(n_38088), .b(n_38087), .o(n_38108) );
oa12f80 g770255 ( .a(n_10777), .b(n_10776), .c(n_10775), .o(n_10840) );
na02f80 g771879 ( .a(n_8860), .b(n_8887), .o(n_8929) );
no02f80 g769937 ( .a(n_11058), .b(FE_OCP_RBN2748_n_9584), .o(n_11131) );
in01f80 g749627 ( .a(n_30299), .o(n_30327) );
in01f80 newInst_2953 ( .a(newNet_2952), .o(newNet_2953) );
in01f80 newInst_2922 ( .a(newNet_253), .o(newNet_2922) );
no02f80 g771535 ( .a(n_9103), .b(FE_OCP_RBN3571_n_44563), .o(n_9341) );
na02f80 g780810 ( .a(n_597), .b(beta_0), .o(n_598) );
in01f80 g775802 ( .a(n_5335), .o(n_5365) );
in01f80 g770136 ( .a(n_10762), .o(n_10763) );
oa22f80 g763870 ( .a(n_16963), .b(n_16260), .c(n_16962), .d(n_16259), .o(n_17103) );
in01f80 g777214 ( .a(n_3605), .o(n_3606) );
na02f80 g772917 ( .a(n_45875), .b(n_7318), .o(n_7868) );
in01f80 g773234 ( .a(n_7657), .o(n_7658) );
oa12f80 g736251 ( .a(n_333), .b(n_43912), .c(FE_OFN4_n_43918), .o(n_43920) );
in01f80 g771340 ( .a(n_9057), .o(n_9114) );
na02f80 g768040 ( .a(n_12914), .b(n_12964), .o(n_13162) );
in01f80 g775381 ( .a(n_46998), .o(n_5933) );
ao12f80 g777920 ( .a(n_3088), .b(n_3111), .c(n_3087), .o(n_4686) );
no02f80 g781099 ( .a(n_239), .b(n_172), .o(n_258) );
in01f80 g741284 ( .a(n_38998), .o(n_38941) );
na02f80 g778760 ( .a(n_2327), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .o(n_2413) );
in01f80 g738867 ( .a(n_41481), .o(n_41286) );
na02f80 g774309 ( .a(FE_OCP_RBN1986_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .o(n_6526) );
no02f80 g765206 ( .a(n_15257), .b(n_15340), .o(n_15413) );
ao12f80 g757370 ( .a(n_22953), .b(n_23400), .c(n_22922), .o(n_23438) );
na02f80 g755178 ( .a(n_25145), .b(n_25176), .o(n_25335) );
in01f80 g779106 ( .a(n_1974), .o(n_1975) );
na02f80 g776989 ( .a(n_4071), .b(n_4070), .o(n_4147) );
oa12f80 g772535 ( .a(n_7492), .b(n_8186), .c(n_7460), .o(n_8231) );
na02f80 FE_RC_3563_0 ( .a(n_23668), .b(n_24934), .o(FE_RN_1547_0) );
na02f80 g746953 ( .a(n_33014), .b(delay_add_ln22_unr20_stage8_stallmux_q_10_), .o(n_33079) );
oa22f80 FE_RC_3364_0 ( .a(n_36194), .b(n_36535), .c(n_36195), .d(FE_OCP_RBN3087_n_36535), .o(n_36632) );
in01f80 g769031 ( .a(n_11786), .o(n_11704) );
in01f80 newInst_1150 ( .a(newNet_1149), .o(newNet_1150) );
no02f80 g763808 ( .a(n_17100), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n_17208) );
in01f80 FE_OCP_RBC2316_n_41420 ( .a(FE_OCP_RBN2315_n_41420), .o(FE_OCP_RBN2316_n_41420) );
in01f80 g741959 ( .a(n_38166), .o(n_38140) );
in01f80 FE_OCP_RBC3592_n_8902 ( .a(n_8902), .o(FE_OCP_RBN3592_n_8902) );
in01f80 newInst_3541 ( .a(newNet_191), .o(newNet_3541) );
in01f80 g778720 ( .a(n_2390), .o(n_2391) );
in01f80 FE_OCP_RBC2652_n_14684 ( .a(n_14684), .o(FE_OCP_RBN2652_n_14684) );
oa12f80 g775060 ( .a(n_5878), .b(n_5970), .c(n_5871), .o(n_6041) );
no02f80 g754087 ( .a(n_26058), .b(n_25994), .o(n_26123) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_1_ ( .ck(newNet_2100), .d(n_4600), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_1_) );
no02f80 g745150 ( .a(n_34725), .b(n_34709), .o(n_34710) );
in01f80 newInst_2985 ( .a(newNet_2984), .o(newNet_2985) );
no02f80 g775514 ( .a(n_5849), .b(n_5891), .o(n_5892) );
oa22f80 g741092 ( .a(FE_OCP_RBN2689_n_38870), .b(n_38404), .c(FE_OCPN957_n_39096), .d(n_38434), .o(n_39274) );
na02f80 g769006 ( .a(n_11650), .b(n_11762), .o(n_11813) );
no02f80 g757603 ( .a(n_23242), .b(n_22887), .o(n_23298) );
in01f80 g754685 ( .a(n_26606), .o(n_26572) );
in01f80 FE_RC_916_0 ( .a(FE_RN_272_0), .o(n_31082) );
na02f80 g757212 ( .a(n_23535), .b(n_22979), .o(n_23566) );
oa12f80 g766147 ( .a(n_14840), .b(n_14839), .c(n_14838), .o(n_15869) );
in01f80 g751182 ( .a(n_29945), .o(n_29877) );
in01f80 newInst_3245 ( .a(newNet_3244), .o(newNet_3245) );
no02f80 FE_RC_2735_0 ( .a(n_38888), .b(n_38852), .o(FE_RN_1159_0) );
no02f80 g745695 ( .a(n_34207), .b(n_34225), .o(n_34289) );
in01f80 newInst_1978 ( .a(newNet_1977), .o(newNet_1978) );
in01f80 newInst_2619 ( .a(newNet_1545), .o(newNet_2619) );
oa12f80 g773048 ( .a(FE_OCPN940_n_7712), .b(n_7807), .c(n_7801), .o(n_7809) );
na02f80 g759760 ( .a(n_21517), .b(n_21478), .o(n_21520) );
no04s80 g762328 ( .a(n_18051), .b(n_18003), .c(n_17971), .d(n_18052), .o(n_18054) );
na02f80 g750329 ( .a(n_29684), .b(n_29671), .o(n_29704) );
no02f80 g737642 ( .a(n_42742), .b(n_42469), .o(n_42799) );
no02f80 g747740 ( .a(n_33393), .b(n_32902), .o(n_33356) );
in01f80 newInst_1904 ( .a(newNet_1903), .o(newNet_1904) );
oa12f80 g739869 ( .a(n_40048), .b(n_40199), .c(n_40254), .o(n_40347) );
in01f80 FE_OCPC3797_n_26115 ( .a(FE_OCPN3796_n_26115), .o(FE_OCPN3797_n_26115) );
na02f80 g780318 ( .a(n_950), .b(n_942), .o(n_979) );
in01f80 g775554 ( .a(n_5645), .o(n_5613) );
in01f80 FE_OCP_RBC2547_n_44944 ( .a(n_44944), .o(FE_OCP_RBN2547_n_44944) );
oa12f80 g759688 ( .a(n_21831), .b(n_21798), .c(n_21691), .o(n_21867) );
na02f80 FE_RC_3185_0 ( .a(FE_RN_1412_0), .b(FE_RN_1413_0), .o(FE_RN_1414_0) );
ao22s80 g780252 ( .a(n_974), .b(n_1203), .c(n_1046), .d(FE_OFN760_n_45813), .o(n_1088) );
na02f80 g748231 ( .a(FE_OCPN880_n_31944), .b(n_30592), .o(n_32072) );
na02f80 g748218 ( .a(n_32766), .b(n_32765), .o(n_32767) );
no02f80 g754213 ( .a(FE_OCP_RBN1202_n_25898), .b(n_23317), .o(n_25945) );
ao12f80 g749883 ( .a(n_30438), .b(n_31065), .c(n_30061), .o(n_31120) );
na02f80 FE_RC_1146_0 ( .a(FE_RN_345_0), .b(FE_RN_346_0), .o(FE_RN_347_0) );
in01f80 g742817 ( .a(n_37245), .o(n_37256) );
na02f80 g761725 ( .a(n_19339), .b(n_18663), .o(n_19369) );
no02f80 g742915 ( .a(n_36965), .b(n_36966), .o(n_37242) );
in01f80 newInst_2479 ( .a(newNet_1034), .o(newNet_2479) );
no02f80 g769069 ( .a(n_11578), .b(n_10916), .o(n_11641) );
na02f80 g737720 ( .a(FE_OCPN887_n_42367), .b(n_42158), .o(n_42746) );
in01f80 newInst_2949 ( .a(newNet_2948), .o(newNet_2949) );
no02f80 g743909 ( .a(n_35916), .b(n_35736), .o(n_35917) );
na02f80 g741330 ( .a(FE_OCP_RBN2546_n_44944), .b(n_38627), .o(n_39148) );
in01f80 g752582 ( .a(n_27634), .o(n_27645) );
in01f80 g776596 ( .a(n_4563), .o(n_4564) );
oa12f80 g765115 ( .a(n_14908), .b(n_15026), .c(n_14909), .o(n_15084) );
no02f80 FE_RC_2839_0 ( .a(FE_RN_1220_0), .b(n_19358), .o(n_19474) );
no02f80 g770385 ( .a(n_10600), .b(n_10585), .o(n_10707) );
na02f80 g736967 ( .a(n_43120), .b(n_42968), .o(n_43303) );
ao12f80 g779259 ( .a(n_1653), .b(n_1789), .c(n_1694), .o(n_1838) );
in01f80 FE_RC_2799_0 ( .a(n_8232), .o(FE_RN_1197_0) );
in01f80 FE_OCP_RBC2633_n_30170 ( .a(n_30170), .o(FE_OCP_RBN2633_n_30170) );
na02f80 g743516 ( .a(n_36549), .b(n_36750), .o(n_36550) );
na02f80 g746282 ( .a(n_33547), .b(n_33527), .o(n_33642) );
in01f80 g762188 ( .a(n_18171), .o(n_18172) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_12_ ( .ck(newNet_3258), .d(n_36388), .o(delay_add_ln22_unr23_stage9_stallmux_q_12_) );
na02f80 g742515 ( .a(n_37515), .b(n_37069), .o(n_37563) );
in01f80 newInst_1723 ( .a(newNet_1722), .o(newNet_1723) );
no02f80 g778038 ( .a(n_2861), .b(n_3020), .o(n_3021) );
oa12f80 g770638 ( .a(n_10352), .b(n_10373), .c(n_10351), .o(n_10420) );
na02f80 g781104 ( .a(n_244), .b(n_237), .o(n_238) );
oa12f80 g753651 ( .a(n_26715), .b(n_27203), .c(n_26792), .o(n_27283) );
in01f80 g777995 ( .a(n_3200), .o(n_3151) );
in01f80 g753987 ( .a(n_27033), .o(n_27034) );
in01f80 FE_RC_3188_0 ( .a(n_17780), .o(FE_RN_1416_0) );
in01f80 g779761 ( .a(n_1749), .o(n_1721) );
na02f80 g770357 ( .a(n_10687), .b(n_10686), .o(n_10688) );
na02f80 g769775 ( .a(n_11004), .b(n_44463), .o(n_11010) );
no02f80 g755396 ( .a(n_24765), .b(n_24764), .o(n_24837) );
in01f80 FE_OCP_RBC2183_FE_RN_464_0 ( .a(FE_RN_464_0), .o(FE_OCP_RBN2183_FE_RN_464_0) );
no02f80 g761930 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n_18674) );
in01f80 newInst_2259 ( .a(newNet_2258), .o(newNet_2259) );
ao12f80 g744005 ( .a(n_36881), .b(n_36882), .c(n_36880), .o(n_37022) );
in01f80 g752904 ( .a(n_28132), .o(n_28078) );
in01f80 fopt783525 ( .a(n_45137), .o(n_45136) );
no02f80 g745992 ( .a(n_33787), .b(FE_OCPN1758_n_33213), .o(n_33810) );
ao12f80 g768803 ( .a(n_12402), .b(FE_OCPN867_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .o(n_12207) );
in01f80 g778684 ( .a(n_2651), .o(n_2639) );
in01f80 g774302 ( .a(n_6770), .o(n_6771) );
in01f80 FE_RC_3489_0 ( .a(n_36999), .o(FE_RN_1504_0) );
in01f80 g759052 ( .a(n_21424), .o(n_21425) );
ao12f80 g742578 ( .a(n_37433), .b(n_37432), .c(n_37431), .o(n_37969) );
in01f80 g768032 ( .a(n_12911), .o(n_13077) );
na02f80 g745883 ( .a(n_35336), .b(n_34800), .o(n_35354) );
in01f80 g744311 ( .a(n_46246), .o(n_36851) );
in01f80 newInst_2216 ( .a(newNet_2215), .o(newNet_2216) );
no02f80 g755164 ( .a(n_25551), .b(n_24642), .o(n_25749) );
in01f80 FE_OCPC1409_n_27014 ( .a(n_27014), .o(FE_OCPN1409_n_27014) );
in01f80 newInst_2399 ( .a(newNet_2398), .o(newNet_2399) );
in01f80 newInst_1935 ( .a(newNet_1934), .o(newNet_1935) );
in01f80 g760218 ( .a(n_20309), .o(n_20268) );
in01f80 FE_OCP_RBC3251_delay_xor_ln22_unr6_stage3_stallmux_q_0_ ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(FE_OCP_RBN3251_delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
in01f80 newInst_105 ( .a(newNet_86), .o(newNet_105) );
na02f80 g738772 ( .a(n_41359), .b(n_41362), .o(n_41384) );
in01f80 g777069 ( .a(n_5333), .o(n_5334) );
no02f80 g739031 ( .a(n_41138), .b(n_41137), .o(n_41139) );
no02f80 g776057 ( .a(n_4989), .b(FE_OCP_RBN2609_n_3807), .o(n_5041) );
in01f80 g764803 ( .a(n_15708), .o(n_15762) );
na02f80 g778568 ( .a(n_2514), .b(n_2496), .o(n_2497) );
in01f80 g756811 ( .a(n_23394), .o(n_23395) );
in01f80 g758632 ( .a(n_21874), .o(n_21875) );
in01f80 g778746 ( .a(n_2212), .o(n_2213) );
in01f80 FE_RC_3922_0 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .o(FE_RN_1696_0) );
no02f80 g775817 ( .a(n_5277), .b(n_5230), .o(n_5354) );
no02f80 FE_RC_2988_0 ( .a(n_46423), .b(FE_RN_1304_0), .o(n_11221) );
ao12f80 g752053 ( .a(n_28015), .b(FE_OCPN878_n_44734), .c(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .o(n_28308) );
in01f80 g740125 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_1_), .o(n_40684) );
ao12f80 g743440 ( .a(n_37681), .b(n_37680), .c(n_46244), .o(n_37789) );
in01f80 newInst_1214 ( .a(newNet_1213), .o(newNet_1214) );
in01f80 FE_OCPC1026_n_25481 ( .a(FE_OCPN1025_n_25481), .o(FE_OCPN1026_n_25481) );
in01f80 g757609 ( .a(n_23260), .o(n_23261) );
na03f80 FE_RC_4132_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_6_), .b(n_32698), .c(n_32699), .o(n_32708) );
na02f80 g740218 ( .a(n_39996), .b(n_39938), .o(n_39997) );
na02f80 g775007 ( .a(n_6109), .b(n_5265), .o(n_6186) );
na02f80 g763602 ( .a(n_16827), .b(n_16825), .o(n_16933) );
na02f80 g746547 ( .a(n_34693), .b(n_34697), .o(n_35242) );
no02f80 g746974 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .o(n_33474) );
na02f80 g751902 ( .a(n_29285), .b(n_29242), .o(n_29581) );
in01f80 newInst_777 ( .a(newNet_272), .o(newNet_777) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_28_ ( .ck(newNet_2370), .d(FE_OCP_RBN3059_n_36515), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_28_) );
no02f80 g779774 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .o(n_1512) );
na02f80 g752203 ( .a(n_27972), .b(n_27971), .o(n_28189) );
in01f80 newInst_2280 ( .a(newNet_1642), .o(newNet_2280) );
no02f80 g775202 ( .a(n_46427), .b(n_5982), .o(n_5983) );
oa12f80 g741220 ( .a(n_39260), .b(FE_OCPN942_n_44925), .c(n_38873), .o(n_39297) );
na02f80 g773900 ( .a(n_7082), .b(n_7081), .o(n_7221) );
in01f80 g774837 ( .a(n_6389), .o(n_6390) );
no02f80 g739070 ( .a(n_41065), .b(n_40868), .o(n_41090) );
in01f80 g747127 ( .a(n_32968), .o(n_32969) );
oa12f80 g767301 ( .a(n_13653), .b(n_13652), .c(n_13651), .o(n_13714) );
in01f80 g769889 ( .a(n_11178), .o(n_11179) );
na02f80 g740683 ( .a(n_39566), .b(n_39454), .o(n_39587) );
no02f80 g747392 ( .a(n_32820), .b(n_32631), .o(n_32678) );
in01f80 g757593 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_26_), .o(n_22859) );
in01f80 g778374 ( .a(n_2770), .o(n_2771) );
no02f80 g753874 ( .a(n_26298), .b(n_26144), .o(n_26300) );
no02f80 g760576 ( .a(n_20356), .b(n_20355), .o(n_20357) );
no02f80 g740935 ( .a(n_39195), .b(n_39083), .o(n_39256) );
in01f80 newInst_27 ( .a(newNet_16), .o(newNet_27) );
ao12f80 g779392 ( .a(n_1444), .b(n_1561), .c(n_1396), .o(n_1628) );
na02f80 g784707 ( .a(n_47183), .b(n_47184), .o(n_47185) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_24_ ( .ck(newNet_2180), .d(n_1005), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_24_) );
in01f80 g745799 ( .a(n_34117), .o(n_34149) );
ao22s80 g777254 ( .a(FE_OCP_RBN3576_n_4528), .b(n_2913), .c(n_4528), .d(n_3029), .o(n_3720) );
in01f80 newInst_1784 ( .a(newNet_73), .o(newNet_1784) );
in01f80 g744570 ( .a(n_35365), .o(n_35352) );
in01f80 g737312 ( .a(n_42876), .o(n_42918) );
na02f80 g758713 ( .a(n_21665), .b(n_21684), .o(n_21689) );
na02f80 g746018 ( .a(n_33835), .b(n_33859), .o(n_33946) );
na02f80 g756492 ( .a(n_23683), .b(n_23682), .o(n_23716) );
na02f80 g752131 ( .a(n_27922), .b(n_44735), .o(n_28043) );
in01f80 newInst_2061 ( .a(newNet_2060), .o(newNet_2061) );
ao12f80 g767429 ( .a(n_13506), .b(n_13505), .c(n_13504), .o(n_13961) );
in01f80 g769984 ( .a(n_10992), .o(n_11049) );
ao12f80 g761206 ( .a(n_19988), .b(n_19904), .c(n_19845), .o(n_20041) );
ao12f80 g755307 ( .a(n_24536), .b(n_24787), .c(n_24535), .o(n_24862) );
in01f80 g776543 ( .a(n_4265), .o(n_4266) );
na02f80 g745191 ( .a(n_36283), .b(n_36221), .o(n_36284) );
na02f80 g761466 ( .a(n_19845), .b(n_19398), .o(n_19909) );
na02f80 g776700 ( .a(FE_OCP_RBN2701_n_4041), .b(n_3951), .o(n_3953) );
in01f80 FE_RC_3711_0 ( .a(n_24323), .o(FE_RN_1632_0) );
in01f80 newInst_2490 ( .a(newNet_2489), .o(newNet_2490) );
no02f80 g747544 ( .a(n_33556), .b(n_33515), .o(n_33557) );
in01f80 g780393 ( .a(n_875), .o(n_928) );
no02f80 FE_RC_2776_0 ( .a(n_38114), .b(n_38111), .o(FE_RN_1184_0) );
na02f80 g744807 ( .a(n_35098), .b(n_30587), .o(n_35141) );
no02f80 g780538 ( .a(n_692), .b(n_705), .o(n_855) );
no02f80 g736327 ( .a(n_43816), .b(n_43637), .o(n_43885) );
ao12f80 g777639 ( .a(n_3398), .b(n_3423), .c(n_3397), .o(n_3470) );
no02f80 g745590 ( .a(n_34261), .b(n_33221), .o(n_34324) );
in01f80 newInst_3496 ( .a(newNet_3495), .o(newNet_3496) );
no02f80 g756549 ( .a(n_23843), .b(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n_23993) );
ao12f80 g784694 ( .a(n_2786), .b(n_2722), .c(n_2137), .o(n_47024) );
na02f80 g778451 ( .a(n_2356), .b(n_1948), .o(n_2457) );
in01f80 newInst_887 ( .a(newNet_154), .o(newNet_887) );
na04m80 g762308 ( .a(n_17930), .b(n_18002), .c(n_17954), .d(n_17893), .o(n_18061) );
no02f80 g752796 ( .a(n_27853), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n_27854) );
oa12f80 g781134 ( .a(n_83), .b(n_214), .c(n_115), .o(n_222) );
in01f80 g780174 ( .a(n_1168), .o(n_1150) );
in01f80 g764948 ( .a(n_15547), .o(n_15548) );
no02f80 g765669 ( .a(n_15070), .b(n_15004), .o(n_15140) );
na02f80 g762791 ( .a(n_17870), .b(n_17823), .o(n_17926) );
ao12f80 g777895 ( .a(n_2902), .b(n_3149), .c(n_2956), .o(n_3236) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_4_ ( .ck(newNet_1573), .d(n_26999), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_) );
in01f80 newInst_2934 ( .a(newNet_2172), .o(newNet_2934) );
oa22f80 FE_RC_1002_0 ( .a(n_45741), .b(n_32752), .c(n_32680), .d(n_32753), .o(n_32829) );
na02f80 g739665 ( .a(n_40534), .b(n_40223), .o(n_40547) );
na02f80 g776208 ( .a(n_4338), .b(n_4264), .o(n_4558) );
in01f80 g763780 ( .a(n_46977), .o(n_16705) );
na02f80 g762201 ( .a(n_18190), .b(n_17947), .o(n_18191) );
in01f80 g749235 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n_32157) );
in01f80 FE_OCPC856_n_20367 ( .a(FE_OCPN855_n_20367), .o(FE_OCPN856_n_20367) );
no02f80 g754006 ( .a(n_26112), .b(n_25672), .o(n_26228) );
na02f80 g739430 ( .a(n_44798), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .o(n_40823) );
no02f80 g765150 ( .a(n_15343), .b(FE_OCP_DRV_N3156_n_15342), .o(n_15380) );
no02f80 g760799 ( .a(n_19473), .b(n_19440), .o(n_19605) );
no02f80 g753182 ( .a(n_25755), .b(n_27103), .o(n_27124) );
in01f80 g753223 ( .a(n_27384), .o(n_27418) );
in01f80 g761298 ( .a(n_19008), .o(n_19033) );
no02f80 g772793 ( .a(n_8137), .b(n_8159), .o(n_8273) );
na02f80 g761559 ( .a(n_18755), .b(n_18721), .o(n_18950) );
na02f80 g745750 ( .a(n_34196), .b(n_34241), .o(n_34685) );
in01f80 newInst_2269 ( .a(newNet_2268), .o(newNet_2269) );
na02f80 g751886 ( .a(n_29332), .b(n_29042), .o(n_29333) );
na02f80 g751212 ( .a(n_29771), .b(n_29760), .o(n_29761) );
oa22f80 FE_RC_4123_0 ( .a(n_33321), .b(n_33773), .c(n_33322), .d(n_33807), .o(n_33872) );
in01f80 g747947 ( .a(n_33169), .o(n_33554) );
oa22f80 g739405 ( .a(n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .c(n_44775), .d(n_40582), .o(n_40983) );
no02f80 g766361 ( .a(n_14163), .b(n_13120), .o(n_14164) );
oa12f80 g756837 ( .a(n_23333), .b(n_23334), .c(n_23332), .o(n_24682) );
in01f80 FE_OFC626_n_34445 ( .a(n_34445), .o(FE_OFN626_n_34445) );
in01f80 g778645 ( .a(n_2550), .o(n_2551) );
na02f80 FE_RC_3606_0 ( .a(FE_RN_1576_0), .b(n_20372), .o(FE_RN_677_0) );
in01f80 newInst_2323 ( .a(newNet_2322), .o(newNet_2323) );
no02f80 g766022 ( .a(n_14996), .b(n_14995), .o(n_14997) );
na02f80 g738557 ( .a(n_41503), .b(FE_OCPN948_n_41382), .o(n_41672) );
no02f80 g747694 ( .a(n_33358), .b(n_33421), .o(n_33443) );
na02f80 g775896 ( .a(n_5351), .b(n_5318), .o(n_5493) );
ms00f80 sin_out_reg_0_ ( .ck(newNet_94), .d(n_43155), .o(sin_out_0) );
in01f80 g755154 ( .a(n_25102), .o(n_25103) );
na02f80 g780504 ( .a(n_752), .b(n_814), .o(n_1195) );
no02f80 g763303 ( .a(n_16996), .b(FE_OCP_RBN2918_n_16084), .o(n_17041) );
in01f80 newInst_3097 ( .a(newNet_3096), .o(newNet_3097) );
no02f80 g747262 ( .a(n_33748), .b(n_33556), .o(n_33801) );
in01f80 FE_RC_2011_0 ( .a(n_18973), .o(FE_RN_663_0) );
na02f80 g751782 ( .a(n_28285), .b(n_28293), .o(n_28294) );
in01f80 FE_OCP_RBC1166_n_18437 ( .a(n_18437), .o(FE_OCP_RBN1166_n_18437) );
in01f80 g740117 ( .a(n_40221), .o(n_40222) );
in01f80 g761336 ( .a(n_19846), .o(n_19847) );
no04s80 FE_RC_3322_0 ( .a(n_16973), .b(n_17129), .c(n_17239), .d(FE_OCP_RBN1136_n_17040), .o(n_17342) );
in01f80 newInst_442 ( .a(newNet_441), .o(newNet_442) );
na02f80 g764151 ( .a(n_16472), .b(FE_OCP_RBN2926_n_16446), .o(n_16517) );
no02f80 g778093 ( .a(n_2924), .b(n_2533), .o(n_2960) );
ao22s80 FE_RC_956_0 ( .a(n_32057), .b(n_32324), .c(n_32058), .d(n_32343), .o(n_32427) );
na02f80 g760055 ( .a(n_20708), .b(n_20748), .o(n_20836) );
na02f80 g749542 ( .a(n_30437), .b(n_30120), .o(n_30496) );
na02f80 g736814 ( .a(n_43144), .b(n_43113), .o(n_43177) );
no02f80 g757740 ( .a(n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(n_22539) );
in01f80 FE_OCP_RBC1353_n_33584 ( .a(n_33584), .o(FE_OCP_RBN1353_n_33584) );
in01f80 FE_OCPC1788_n_36034 ( .a(FE_OCPN1787_n_36034), .o(FE_OCPN1788_n_36034) );
in01f80 FE_OCP_RBC2643_FE_RN_1198_0 ( .a(FE_RN_1198_0), .o(FE_OCP_RBN2643_FE_RN_1198_0) );
in01f80 g756572 ( .a(n_23584), .o(n_23609) );
in01f80 g748988 ( .a(n_32314), .o(n_32315) );
na02f80 FE_RC_2523_0 ( .a(n_44769), .b(FE_RN_1027_0), .o(FE_RN_1028_0) );
oa12f80 g756705 ( .a(n_23516), .b(n_23504), .c(n_23515), .o(n_23604) );
na02f80 g762623 ( .a(n_18105), .b(n_18068), .o(n_18124) );
no02f80 g754410 ( .a(n_25656), .b(n_25360), .o(n_25678) );
oa12f80 g780759 ( .a(n_566), .b(n_565), .c(n_564), .o(n_693) );
no02f80 g743470 ( .a(FE_OCP_RBN3058_n_36515), .b(n_36750), .o(n_36554) );
na02f80 g761440 ( .a(n_18761), .b(n_17661), .o(n_18875) );
na02f80 g767269 ( .a(n_13490), .b(n_13458), .o(n_13559) );
no02f80 FE_RC_377_0 ( .a(FE_RN_111_0), .b(FE_RN_112_0), .o(FE_RN_113_0) );
in01f80 g780333 ( .a(FE_OCPN1394_n_962), .o(n_1009) );
no02f80 g739996 ( .a(n_40255), .b(n_40059), .o(n_40256) );
ao12f80 g761091 ( .a(n_18396), .b(n_19088), .c(n_18394), .o(n_19184) );
no02f80 g764561 ( .a(n_15952), .b(n_15849), .o(n_16047) );
na02f80 g748044 ( .a(n_32880), .b(n_32826), .o(n_32966) );
in01f80 g743652 ( .a(n_36416), .o(n_36397) );
ao22s80 FE_RC_3867_0 ( .a(n_30259), .b(n_30623), .c(n_30260), .d(n_30605), .o(n_30731) );
no02f80 g740405 ( .a(FE_OCP_RBN3022_n_39942), .b(n_39543), .o(n_40059) );
in01f80 g758326 ( .a(n_22212), .o(n_22298) );
in01f80 g741700 ( .a(n_38579), .o(n_38580) );
no02f80 g750653 ( .a(n_29280), .b(n_28801), .o(n_29347) );
in01f80 g777590 ( .a(n_3507), .o(n_3477) );
na02f80 g776664 ( .a(n_4029), .b(n_4039), .o(n_4218) );
no02f80 g751767 ( .a(n_28301), .b(n_28300), .o(n_28302) );
na02f80 FE_RC_2332_0 ( .a(FE_RN_890_0), .b(n_6517), .o(FE_RN_891_0) );
no02f80 g748124 ( .a(n_31906), .b(n_31835), .o(n_31952) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_5_ ( .ck(newNet_214), .d(n_46153), .o(delay_xor_ln22_unr6_stage3_stallmux_q_5_) );
na02f80 g779535 ( .a(n_1527), .b(n_1780), .o(n_1528) );
na02f80 g761778 ( .a(n_18555), .b(n_18477), .o(n_18710) );
no02f80 g747868 ( .a(n_33193), .b(n_33192), .o(n_33194) );
na02f80 g770884 ( .a(n_9964), .b(n_9624), .o(n_10052) );
in01f80 newInst_3115 ( .a(newNet_1828), .o(newNet_3115) );
in01f80 g776635 ( .a(n_4352), .o(n_4353) );
ao12f80 g756528 ( .a(n_23830), .b(n_24078), .c(n_23721), .o(n_24114) );
in01f80 FE_RC_753_0 ( .a(FE_RN_236_0), .o(n_28002) );
in01f80 newInst_1574 ( .a(newNet_1347), .o(newNet_1574) );
oa12f80 g784667 ( .a(n_5928), .b(n_5902), .c(n_5761), .o(n_46997) );
na02f80 g779174 ( .a(n_1959), .b(n_1665), .o(n_1993) );
na02f80 g773733 ( .a(n_7264), .b(n_7242), .o(n_7243) );
na02f80 g762357 ( .a(FE_OCP_RBN3409_n_45120), .b(n_17860), .o(n_18578) );
oa22f80 FE_RC_1236_0 ( .a(FE_OFN84_n_46137), .b(n_6589), .c(FE_OFN806_n_46196), .d(n_6627), .o(n_46187) );
in01f80 newInst_54 ( .a(newNet_19), .o(newNet_54) );
na02f80 g778156 ( .a(n_2802), .b(n_2793), .o(n_3502) );
na02f80 g781108 ( .a(n_241), .b(n_549), .o(n_242) );
in01f80 g743973 ( .a(n_36069), .o(n_36070) );
in01f80 g736719 ( .a(n_43282), .o(n_43283) );
na02f80 g773858 ( .a(n_7073), .b(n_6869), .o(n_7118) );
oa12f80 g740970 ( .a(n_39105), .b(n_39163), .c(n_39133), .o(n_39212) );
in01f80 g742732 ( .a(n_37397), .o(n_37444) );
in01f80 newInst_3484 ( .a(newNet_2435), .o(newNet_3484) );
in01f80 newInst_1241 ( .a(newNet_366), .o(newNet_1241) );
no02f80 FE_RC_315_0 ( .a(FE_RN_95_0), .b(n_21034), .o(n_46968) );
na02f80 g765499 ( .a(n_15719), .b(n_15958), .o(n_15875) );
na02f80 g770085 ( .a(n_10761), .b(n_9114), .o(n_10825) );
in01f80 FE_RC_1051_0 ( .a(FE_RN_308_0), .o(n_15396) );
in01f80 newInst_1033 ( .a(newNet_1032), .o(newNet_1033) );
in01f80 g752837 ( .a(n_28276), .o(n_28277) );
in01f80 fopt782828 ( .a(n_44256), .o(n_44221) );
no02f80 FE_RC_4180_0 ( .a(FE_RN_1824_0), .b(FE_RN_1826_0), .o(FE_RN_1827_0) );
no02f80 g764777 ( .a(n_15649), .b(n_15696), .o(n_15738) );
ao22s80 FE_RC_210_0 ( .a(n_14198), .b(n_14246), .c(n_14153), .d(n_14248), .o(n_14450) );
no02f80 g771299 ( .a(n_9267), .b(n_9051), .o(n_9357) );
in01f80 g744113 ( .a(n_35640), .o(n_35641) );
no02f80 g770793 ( .a(n_9867), .b(n_9858), .o(n_10023) );
in01f80 FE_OCP_RBC3688_n_5130 ( .a(n_5130), .o(FE_OCP_RBN3688_n_5130) );
in01f80 g740729 ( .a(n_39446), .o(n_39447) );
in01f80 g757970 ( .a(n_22086), .o(n_22110) );
oa12f80 g744502 ( .a(n_35403), .b(n_35402), .c(n_35414), .o(n_35426) );
na02f80 g750394 ( .a(n_29624), .b(n_29615), .o(n_29646) );
na02f80 g757261 ( .a(n_23137), .b(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(n_23133) );
no02f80 g763514 ( .a(FE_OCP_RBN3079_n_16977), .b(FE_OCPN869_n_16086), .o(n_17117) );
no02f80 g745381 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35845), .o(n_35882) );
no02f80 g745099 ( .a(n_35613), .b(n_34706), .o(n_34895) );
in01f80 g744641 ( .a(n_35343), .o(n_35344) );
no02f80 g776704 ( .a(n_4076), .b(n_3912), .o(n_4077) );
in01f80 FE_OCP_RBC3000_n_42959 ( .a(n_42959), .o(FE_OCP_RBN3000_n_42959) );
na02f80 g754161 ( .a(n_25975), .b(n_25506), .o(n_26022) );
in01f80 g740535 ( .a(n_39683), .o(n_39684) );
no02f80 g756321 ( .a(n_24587), .b(n_23936), .o(n_24585) );
no02f80 g771991 ( .a(n_44570), .b(n_10137), .o(n_8916) );
in01f80 newInst_2013 ( .a(newNet_2012), .o(newNet_2013) );
no02f80 g778616 ( .a(n_2350), .b(n_2330), .o(n_2959) );
oa22f80 g743078 ( .a(n_36014), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .d(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_37313) );
no02f80 g757988 ( .a(n_22098), .b(n_22134), .o(n_22135) );
ao12f80 g741074 ( .a(n_38887), .b(FE_OCPN957_n_39096), .c(n_38862), .o(n_39301) );
no02f80 g779604 ( .a(n_1367), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1405) );
in01f80 g736747 ( .a(n_43465), .o(n_43466) );
in01f80 newInst_3523 ( .a(newNet_3522), .o(newNet_3523) );
na02f80 g767779 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_26_), .o(n_13000) );
in01f80 FE_OCPC1033_n_28420 ( .a(n_28420), .o(FE_OCPN1033_n_28420) );
in01f80 FE_RC_1738_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(FE_RN_485_0) );
oa12f80 g746560 ( .a(n_33052), .b(n_33254), .c(n_33012), .o(n_33306) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_22_ ( .ck(newNet_2847), .d(n_11856), .o(delay_add_ln22_unr8_stage4_stallmux_q_22_) );
no02f80 g743492 ( .a(n_36609), .b(n_36580), .o(n_36667) );
oa12f80 g784679 ( .a(n_4095), .b(n_4026), .c(n_4000), .o(n_47009) );
in01f80 newInst_2869 ( .a(newNet_2868), .o(newNet_2869) );
in01f80 newInst_1201 ( .a(newNet_1200), .o(newNet_1201) );
na02f80 g769849 ( .a(n_11176), .b(n_11211), .o(n_11261) );
in01f80 newInst_2365 ( .a(newNet_2364), .o(newNet_2365) );
na02f80 g750551 ( .a(n_29419), .b(n_29260), .o(n_29476) );
no02f80 g740425 ( .a(FE_OCP_RBN3026_n_39942), .b(FE_OCP_RBN2896_n_39575), .o(n_40247) );
na02f80 FE_RC_2666_0 ( .a(n_4133), .b(n_3954), .o(FE_RN_1114_0) );
no02f80 g753478 ( .a(n_26784), .b(n_26749), .o(n_26827) );
no02f80 g751164 ( .a(n_29944), .b(n_29709), .o(n_30089) );
in01f80 fopt782981 ( .a(n_12065), .o(n_44451) );
in01f80 newInst_1309 ( .a(newNet_1308), .o(newNet_1309) );
na02f80 g754026 ( .a(n_26978), .b(n_26863), .o(n_26979) );
ao12f80 g750164 ( .a(n_29794), .b(n_29793), .c(n_29792), .o(n_31303) );
no02f80 g745704 ( .a(n_34199), .b(n_34247), .o(n_34273) );
in01f80 g777446 ( .a(FE_OCP_RBN2583_n_3734), .o(n_3912) );
na02f80 g770230 ( .a(n_10709), .b(FE_OCPN955_n_44460), .o(n_10710) );
oa22f80 g778936 ( .a(n_2214), .b(n_1984), .c(n_2257), .d(n_1983), .o(n_2297) );
na02f80 g767956 ( .a(n_12811), .b(n_12832), .o(n_12857) );
no04s80 FE_RC_3704_0 ( .a(n_32602), .b(n_32600), .c(n_32547), .d(n_32625), .o(n_32626) );
in01f80 g764733 ( .a(n_15895), .o(n_15896) );
no02f80 g746302 ( .a(n_33635), .b(n_33233), .o(n_33674) );
na02f80 g741900 ( .a(n_38338), .b(n_38017), .o(n_38205) );
no02f80 g776630 ( .a(n_4235), .b(n_4209), .o(n_4302) );
in01f80 newInst_1698 ( .a(newNet_1697), .o(newNet_1698) );
no02f80 g778605 ( .a(n_2654), .b(n_2661), .o(n_3280) );
oa12f80 g738230 ( .a(n_41663), .b(n_41940), .c(n_41558), .o(n_41966) );
oa12f80 g777822 ( .a(n_3243), .b(n_3239), .c(n_3241), .o(n_3299) );
no02f80 g765228 ( .a(n_15569), .b(n_15483), .o(n_15637) );
ao12f80 g759239 ( .a(n_20531), .b(n_20926), .c(n_20535), .o(n_20945) );
in01f80 g740012 ( .a(n_39849), .o(n_39874) );
in01f80 g768714 ( .a(n_12068), .o(n_12064) );
in01f80 newInst_1504 ( .a(newNet_1113), .o(newNet_1504) );
in01f80 g777280 ( .a(n_4731), .o(n_4732) );
in01f80 g753138 ( .a(n_27492), .o(n_27493) );
in01f80 g775340 ( .a(n_5966), .o(n_5967) );
oa12f80 g746512 ( .a(n_34421), .b(n_34420), .c(n_34419), .o(n_34814) );
in01f80 g747402 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n_32623) );
na02f80 g765298 ( .a(n_15874), .b(n_15870), .o(n_15923) );
no02f80 g777333 ( .a(n_3637), .b(n_3472), .o(n_3748) );
na02f80 g769678 ( .a(n_11256), .b(n_44511), .o(n_11299) );
na02f80 g760189 ( .a(n_20304), .b(n_20288), .o(n_20400) );
no02f80 g773481 ( .a(n_7526), .b(n_7256), .o(n_7544) );
no02f80 g752760 ( .a(n_27437), .b(n_27121), .o(n_27439) );
no02f80 g767815 ( .a(n_13241), .b(n_13271), .o(n_13790) );
oa12f80 g760722 ( .a(n_20202), .b(n_20201), .c(n_20200), .o(n_21835) );
in01f80 FE_OCP_RBC2123_n_45224 ( .a(FE_OCP_RBN2122_n_45224), .o(FE_OCP_RBN2123_n_45224) );
in01f80 g776571 ( .a(n_4321), .o(n_4322) );
oa12f80 g762176 ( .a(n_18169), .b(n_18194), .c(n_18168), .o(n_19807) );
no02f80 g743588 ( .a(n_36532), .b(n_36531), .o(n_36533) );
na02f80 g773525 ( .a(n_7440), .b(delay_add_ln22_unr5_stage3_stallmux_q_22_), .o(n_8406) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_4_ ( .ck(newNet_1472), .d(n_31690), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_) );
no02f80 g759068 ( .a(n_21494), .b(FE_OCP_DRV_N1600_n_21493), .o(n_21529) );
na02f80 g743893 ( .a(n_35868), .b(n_35830), .o(n_35987) );
na02f80 g764367 ( .a(n_16225), .b(n_46421), .o(n_16369) );
in01f80 g757296 ( .a(n_23173), .o(n_23132) );
na02f80 g780487 ( .a(n_675), .b(n_674), .o(n_676) );
na02f80 g768058 ( .a(FE_OCPN860_n_12880), .b(n_12738), .o(n_12963) );
no02f80 g763503 ( .a(n_16814), .b(FE_OCPN3180_FE_OCP_RBN2744_n_15319), .o(n_16837) );
oa22f80 FE_RC_1188_0 ( .a(n_18457), .b(n_19041), .c(n_18456), .d(n_19059), .o(n_19219) );
no03m80 FE_RC_2455_0 ( .a(n_13350), .b(n_13378), .c(n_13379), .o(FE_RN_983_0) );
in01f80 newInst_2645 ( .a(newNet_2644), .o(newNet_2645) );
no02f80 g777810 ( .a(n_3250), .b(n_2759), .o(n_3383) );
na02f80 g775042 ( .a(n_6009), .b(n_5726), .o(n_6048) );
oa12f80 g739872 ( .a(n_40039), .b(n_40298), .c(n_39973), .o(n_40381) );
no02f80 g771650 ( .a(n_8938), .b(n_8912), .o(n_9086) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_29_ ( .ck(newNet_2831), .d(n_12212), .o(delay_add_ln22_unr8_stage4_stallmux_q_29_) );
na02f80 g741722 ( .a(n_38458), .b(n_38350), .o(n_38504) );
no02f80 g759056 ( .a(n_21490), .b(FE_OCP_RBN2951_n_21489), .o(n_21630) );
in01f80 g749056 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .o(n_32271) );
in01f80 newInst_424 ( .a(newNet_61), .o(newNet_424) );
no02f80 g760228 ( .a(n_20244), .b(n_20243), .o(n_20303) );
no02f80 g753095 ( .a(n_27145), .b(n_27118), .o(n_27187) );
na02f80 g767045 ( .a(FE_OCP_RBN3529_n_13765), .b(n_13934), .o(n_14035) );
oa12f80 g736344 ( .a(n_43326), .b(n_43789), .c(n_43361), .o(n_43829) );
in01f80 FE_OCP_RBC3546_n_44575 ( .a(n_44575), .o(FE_OCP_RBN3546_n_44575) );
no02f80 FE_RC_3109_0 ( .a(n_26846), .b(n_26970), .o(FE_RN_1376_0) );
na02f80 g752484 ( .a(n_27685), .b(n_27709), .o(n_27771) );
in01f80 newInst_3036 ( .a(newNet_851), .o(newNet_3036) );
na02f80 g758126 ( .a(n_44267), .b(n_21265), .o(n_22258) );
in01f80 g766908 ( .a(n_13907), .o(n_13908) );
in01f80 g758975 ( .a(n_22030), .o(n_22119) );
in01f80 g745370 ( .a(n_35890), .o(n_35848) );
in01f80 g753605 ( .a(n_27367), .o(n_27368) );
in01f80 g779452 ( .a(n_2001), .o(n_2002) );
in01f80 g775366 ( .a(n_5805), .o(n_5806) );
no02f80 g748109 ( .a(n_32838), .b(n_32837), .o(n_32839) );
na02f80 g776050 ( .a(n_47005), .b(FE_OCP_RBN2534_n_47018), .o(n_5108) );
no02f80 g777793 ( .a(n_3375), .b(n_3308), .o(n_3413) );
in01f80 newInst_1967 ( .a(newNet_624), .o(newNet_1967) );
na02f80 g750660 ( .a(n_29278), .b(FE_OFN788_n_25834), .o(n_29380) );
in01f80 FE_RC_2087_0 ( .a(FE_RN_716_0), .o(n_14511) );
na02f80 FE_RC_4251_0 ( .a(n_26872), .b(FE_RN_1870_0), .o(n_26963) );
in01f80 newInst_1645 ( .a(newNet_1644), .o(newNet_1645) );
na02f80 g752813 ( .a(n_27788), .b(n_27882), .o(n_27907) );
in01f80 FE_OCP_RBC3651_n_39249 ( .a(n_39249), .o(FE_OCP_RBN3651_n_39249) );
no02f80 g777885 ( .a(n_3275), .b(n_3274), .o(n_3309) );
na02f80 g742658 ( .a(n_37401), .b(n_37418), .o(n_37505) );
in01f80 fopt782902 ( .a(n_44347), .o(n_44346) );
in01f80 g780931 ( .a(n_489), .o(n_475) );
in01f80 newInst_3123 ( .a(newNet_3122), .o(newNet_3123) );
in01f80 newInst_135 ( .a(newNet_134), .o(newNet_135) );
no02f80 g778323 ( .a(n_2869), .b(delay_add_ln22_unr2_stage2_stallmux_q_28_), .o(n_3857) );
na02f80 g775348 ( .a(n_5786), .b(n_5767), .o(n_5830) );
no02f80 g751845 ( .a(n_29172), .b(n_28919), .o(n_29148) );
na02f80 g777314 ( .a(FE_OCP_RBN2692_FE_OCPN843_n_3912), .b(n_4142), .o(n_4215) );
ao12f80 g752730 ( .a(n_27906), .b(n_27956), .c(n_27928), .o(n_28052) );
in01f80 newInst_2930 ( .a(newNet_2929), .o(newNet_2930) );
in01f80 g780866 ( .a(n_363), .o(n_364) );
oa12f80 g777924 ( .a(n_2655), .b(n_3111), .c(n_3108), .o(n_3112) );
na02f80 g759334 ( .a(n_21070), .b(n_20519), .o(n_21177) );
no02f80 g784786 ( .a(FE_OCP_RBN3085_n_31819), .b(n_30733), .o(n_47272) );
na02f80 g772515 ( .a(n_8433), .b(n_8009), .o(n_8469) );
oa12f80 g758665 ( .a(n_21622), .b(n_22395), .c(n_21561), .o(n_22485) );
na02f80 g742713 ( .a(n_37444), .b(n_44038), .o(n_37454) );
no02f80 g767055 ( .a(FE_OCP_RBN3529_n_13765), .b(n_13961), .o(n_13972) );
in01f80 g741554 ( .a(n_38667), .o(n_38678) );
no02f80 g761483 ( .a(n_19649), .b(n_19758), .o(n_19792) );
na02f80 g744231 ( .a(n_46203), .b(n_46214), .o(n_36841) );
in01f80 g741918 ( .a(n_38146), .o(n_38147) );
na02f80 g775501 ( .a(n_5486), .b(n_5442), .o(n_5496) );
in01f80 g737398 ( .a(n_42790), .o(n_42808) );
in01f80 g743709 ( .a(n_36325), .o(n_36326) );
no02f80 FE_RC_2360_0 ( .a(n_18769), .b(n_18724), .o(FE_RN_912_0) );
in01f80 g743263 ( .a(n_36831), .o(n_36842) );
in01f80 newInst_768 ( .a(newNet_487), .o(newNet_768) );
no02f80 g775193 ( .a(n_46996), .b(n_6030), .o(n_6069) );
in01f80 g752914 ( .a(n_28128), .o(n_28174) );
in01f80 g748571 ( .a(n_32676), .o(n_32677) );
na02f80 g736934 ( .a(n_43038), .b(n_43106), .o(n_43149) );
ao12f80 g750629 ( .a(n_29374), .b(n_29373), .c(n_29372), .o(n_29441) );
oa12f80 g736474 ( .a(n_43375), .b(n_43664), .c(n_43272), .o(n_43726) );
ao12f80 g738906 ( .a(n_41278), .b(n_41277), .c(n_41276), .o(n_41316) );
no02f80 g772857 ( .a(n_8067), .b(n_8066), .o(n_8068) );
oa12f80 g765365 ( .a(n_15867), .b(n_16245), .c(n_15823), .o(n_16253) );
in01f80 g775252 ( .a(n_5938), .o(n_5939) );
oa22f80 g763313 ( .a(n_16916), .b(FE_OFN767_n_15670), .c(n_16872), .d(n_16339), .o(n_17004) );
in01f80 g769626 ( .a(n_11409), .o(n_11490) );
na02f80 g755189 ( .a(n_24993), .b(n_25019), .o(n_25098) );
ao12f80 g778076 ( .a(n_2561), .b(n_2924), .c(n_2501), .o(n_2991) );
na02f80 g749620 ( .a(n_31644), .b(n_31643), .o(n_31645) );
oa12f80 g782636 ( .a(FE_OCP_RBN3444_n_37945), .b(n_37985), .c(n_37638), .o(n_44029) );
in01f80 g740584 ( .a(n_39629), .o(n_39630) );
in01f80 newInst_2360 ( .a(newNet_1028), .o(newNet_2360) );
na02f80 g746949 ( .a(n_32857), .b(n_32381), .o(n_32941) );
na02f80 g765329 ( .a(n_13785), .b(n_15048), .o(n_15081) );
oa22f80 g739826 ( .a(n_40263), .b(n_40019), .c(n_40264), .d(n_40018), .o(n_40385) );
in01f80 g780679 ( .a(n_666), .o(n_679) );
na02f80 g756709 ( .a(n_23482), .b(n_23112), .o(n_23483) );
no02f80 g754799 ( .a(n_26034), .b(n_25408), .o(n_26163) );
oa12f80 g746729 ( .a(n_32821), .b(n_32980), .c(n_32788), .o(n_33039) );
na02f80 g774373 ( .a(n_6783), .b(n_6782), .o(n_7473) );
no02f80 g760201 ( .a(FE_OCPN1261_n_20242), .b(n_19641), .o(n_20366) );
in01f80 g756782 ( .a(n_23397), .o(n_23429) );
na02f80 g779305 ( .a(n_1636), .b(n_47027), .o(n_1736) );
no02f80 g752966 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .o(n_28198) );
in01f80 newInst_3013 ( .a(newNet_3012), .o(newNet_3013) );
in01f80 FE_OCP_RBC2256_n_37844 ( .a(FE_OCP_RBN2255_n_37844), .o(FE_OCP_RBN2256_n_37844) );
oa12f80 g751779 ( .a(n_28910), .b(n_28911), .c(n_28909), .o(n_29799) );
in01f80 newInst_2132 ( .a(newNet_2131), .o(newNet_2132) );
oa12f80 g738612 ( .a(n_41528), .b(n_41713), .c(n_41286), .o(n_42162) );
ao12f80 g774233 ( .a(n_6758), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln22_unr6_stage3_stallmux_q_9_), .o(n_6882) );
no02f80 g778598 ( .a(n_2652), .b(n_3108), .o(n_3087) );
no02f80 g774328 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .o(n_6633) );
no02f80 g758859 ( .a(n_21764), .b(n_21763), .o(n_21783) );
no02f80 g747448 ( .a(n_32593), .b(n_32568), .o(n_32630) );
no02f80 g778392 ( .a(FE_OCP_RBN2266_n_2430), .b(n_2461), .o(n_2462) );
no02f80 g765144 ( .a(n_16100), .b(FE_OFN764_n_15670), .o(n_16101) );
na02f80 g761877 ( .a(n_18512), .b(n_18511), .o(n_18546) );
in01f80 g744891 ( .a(n_35134), .o(n_35095) );
in01f80 g780706 ( .a(n_635), .o(n_636) );
in01f80 fopt784719 ( .a(n_11035), .o(n_47200) );
in01f80 FE_OCP_RBC3633_n_20568 ( .a(FE_OCP_RBN3632_n_20568), .o(FE_OCP_RBN3633_n_20568) );
na02f80 g767931 ( .a(n_12816), .b(n_11524), .o(n_12955) );
in01f80 g776399 ( .a(n_4466), .o(n_4467) );
na02f80 g770874 ( .a(n_9851), .b(n_44818), .o(n_9866) );
ao12f80 g756315 ( .a(n_24515), .b(n_24514), .c(n_24513), .o(n_24605) );
in01f80 g779523 ( .a(n_2359), .o(n_2360) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_12_ ( .ck(newNet_521), .d(n_22973), .o(delay_xor_ln22_unr15_stage6_stallmux_q_12_) );
in01f80 g744711 ( .a(n_36571), .o(n_36572) );
ao12f80 g780687 ( .a(n_651), .b(n_650), .c(n_649), .o(n_859) );
in01f80 g749138 ( .a(n_30877), .o(n_30878) );
in01f80 g744916 ( .a(n_34982), .o(n_35980) );
oa12f80 g754583 ( .a(n_26641), .b(n_26896), .c(n_26605), .o(n_26926) );
na02f80 g777661 ( .a(n_3458), .b(n_3457), .o(n_3459) );
in01f80 g750769 ( .a(n_29217), .o(n_29231) );
in01f80 g780615 ( .a(n_913), .o(n_914) );
in01f80 g750993 ( .a(n_28963), .o(n_28964) );
no03m80 FE_RC_786_0 ( .a(n_33567), .b(n_33642), .c(n_47249), .o(n_33647) );
in01f80 g776879 ( .a(n_4099), .o(n_4100) );
in01f80 g753599 ( .a(n_26748), .o(n_26749) );
na02f80 g760648 ( .a(n_19663), .b(n_18119), .o(n_19708) );
oa22f80 g757230 ( .a(n_23042), .b(n_23204), .c(n_23191), .d(n_23205), .o(n_24425) );
no02f80 g751953 ( .a(n_28836), .b(n_28923), .o(n_29223) );
no02f80 g777771 ( .a(n_3299), .b(n_47020), .o(n_3325) );
in01f80 g738642 ( .a(FE_OCP_RBN2313_n_41420), .o(n_41540) );
no02f80 g778163 ( .a(n_2715), .b(n_2714), .o(n_2716) );
in01f80 FE_RC_2934_0 ( .a(FE_OCP_RBN1164_n_13726), .o(FE_RN_1279_0) );
in01f80 g740641 ( .a(n_39577), .o(n_39576) );
in01f80 g765878 ( .a(n_14903), .o(n_14919) );
no02f80 g749755 ( .a(n_29905), .b(n_29904), .o(n_29906) );
na02f80 g753392 ( .a(n_46422), .b(n_26961), .o(n_27012) );
in01f80 FE_RC_312_0 ( .a(n_20963), .o(FE_RN_93_0) );
in01f80 FE_OCP_RBC2966_n_26231 ( .a(FE_OCP_RBN2963_n_26231), .o(FE_OCP_RBN2966_n_26231) );
in01f80 FE_OCP_RBC2172_n_32892 ( .a(FE_OCP_RBN2170_n_32892), .o(FE_OCP_RBN2172_n_32892) );
in01f80 newInst_1318 ( .a(newNet_1317), .o(newNet_1318) );
oa12f80 g758625 ( .a(n_21646), .b(n_21964), .c(n_21647), .o(n_21987) );
no02f80 g764706 ( .a(n_15801), .b(n_15799), .o(n_15942) );
no02f80 g766728 ( .a(n_14139), .b(n_13903), .o(n_14220) );
in01f80 g752648 ( .a(n_27555), .o(n_27556) );
na02f80 g777133 ( .a(n_3654), .b(n_3679), .o(n_3790) );
in01f80 g780261 ( .a(n_1018), .o(n_975) );
no02f80 g737348 ( .a(n_42833), .b(n_42399), .o(n_42842) );
in01f80 g757635 ( .a(n_22897), .o(n_22856) );
in01f80 g751065 ( .a(n_28869), .o(n_28870) );
na02f80 g781071 ( .a(cos_out_13), .b(FE_OFN2_n_43918), .o(n_346) );
na02f80 g769760 ( .a(n_11123), .b(n_11122), .o(n_11124) );
oa12f80 g765746 ( .a(n_14718), .b(n_14862), .c(n_14717), .o(n_14942) );
na02f80 g742222 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38290), .o(n_38323) );
ao12f80 g748777 ( .a(n_32461), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n_33121) );
in01f80 g756028 ( .a(n_25033), .o(n_24999) );
na02f80 g781304 ( .a(n_46055), .b(beta_7), .o(n_118) );
in01f80 g766768 ( .a(n_13694), .o(n_13663) );
in01f80 g753906 ( .a(n_26421), .o(n_26422) );
in01f80 FE_RC_84_0 ( .a(n_17339), .o(FE_RN_25_0) );
na02f80 g757386 ( .a(n_22942), .b(n_22941), .o(n_23019) );
in01f80 g744365 ( .a(n_46219), .o(n_36816) );
na02f80 g767845 ( .a(n_12853), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_21_), .o(n_12986) );
in01f80 g771398 ( .a(n_9721), .o(n_9722) );
in01f80 g763269 ( .a(n_17283), .o(n_17274) );
in01f80 g778826 ( .a(n_3029), .o(n_3297) );
na02f80 g755404 ( .a(n_24762), .b(n_24761), .o(n_24763) );
no02f80 g780819 ( .a(n_364), .b(n_371), .o(n_380) );
in01f80 FE_RC_4019_0 ( .a(FE_RN_1746_0), .o(n_20689) );
na02f80 FE_RC_2483_0 ( .a(n_9728), .b(n_9693), .o(FE_RN_1002_0) );
ao12f80 g756408 ( .a(n_23720), .b(n_23742), .c(n_23719), .o(n_23792) );
na02f80 g755558 ( .a(n_24571), .b(n_24532), .o(n_24648) );
in01f80 newInst_500 ( .a(newNet_255), .o(newNet_500) );
na02f80 g771529 ( .a(n_9470), .b(n_9327), .o(n_9521) );
in01f80 newInst_2190 ( .a(newNet_1667), .o(newNet_2190) );
in01f80 g768266 ( .a(n_12602), .o(n_12603) );
ao12f80 g755780 ( .a(n_25257), .b(n_25256), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25371) );
no02f80 g763853 ( .a(n_16638), .b(FE_OCP_RBN2694_n_15083), .o(n_16715) );
in01f80 g766743 ( .a(n_13944), .o(n_13909) );
no02f80 g761153 ( .a(n_20037), .b(n_20036), .o(n_20038) );
in01f80 g778570 ( .a(n_2503), .o(n_2504) );
oa12f80 g751015 ( .a(n_29907), .b(n_29886), .c(n_29818), .o(n_29887) );
no02f80 g776325 ( .a(n_4766), .b(n_4728), .o(n_5156) );
in01f80 g774757 ( .a(n_6398), .o(n_6399) );
na02f80 g770153 ( .a(n_10711), .b(n_10253), .o(n_10760) );
na02f80 g737433 ( .a(n_42705), .b(n_42451), .o(n_42706) );
in01f80 g765521 ( .a(n_15924), .o(n_15866) );
na02f80 g778974 ( .a(n_2101), .b(n_1741), .o(n_2144) );
na02f80 g757190 ( .a(n_23197), .b(n_23196), .o(n_23234) );
no03m80 g763758 ( .a(n_17354), .b(n_17426), .c(n_17425), .o(n_17499) );
in01f80 newInst_1334 ( .a(newNet_1333), .o(newNet_1334) );
in01f80 g749601 ( .a(n_30572), .o(n_30592) );
na02f80 g781240 ( .a(n_106), .b(n_128), .o(n_138) );
in01f80 FE_OCP_RBC2377_n_29480 ( .a(FE_OCP_RBN2376_n_29480), .o(FE_OCP_RBN2377_n_29480) );
na02f80 g745801 ( .a(n_44100), .b(n_34118), .o(n_34130) );
in01f80 g778521 ( .a(n_2614), .o(n_2694) );
no02f80 g745295 ( .a(n_35934), .b(n_35888), .o(n_35964) );
no02f80 g761968 ( .a(n_18705), .b(n_18589), .o(n_18706) );
in01f80 FE_OCP_RBC1685_n_18986 ( .a(n_18986), .o(FE_OCP_RBN1685_n_18986) );
na02f80 g745818 ( .a(n_44104), .b(n_33605), .o(n_34203) );
na02f80 g769246 ( .a(FE_OCP_RBN3094_n_11475), .b(n_10480), .o(n_11624) );
in01f80 g755660 ( .a(n_24612), .o(n_24632) );
oa22f80 g762174 ( .a(n_18138), .b(n_18108), .c(n_18095), .d(n_18107), .o(n_19801) );
na02f80 g763104 ( .a(n_17409), .b(FE_OCP_RBN3211_n_44365), .o(n_17458) );
in01f80 g746809 ( .a(n_33321), .o(n_33322) );
no02f80 g742131 ( .a(n_38310), .b(n_38249), .o(n_38353) );
no02f80 g741598 ( .a(n_38601), .b(n_38778), .o(n_38617) );
ao12f80 g751299 ( .a(n_29655), .b(n_29654), .c(n_29653), .o(n_29942) );
in01f80 g759413 ( .a(n_20825), .o(n_20826) );
no02f80 g743377 ( .a(n_36584), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36635) );
na02f80 g738395 ( .a(n_41679), .b(n_41694), .o(n_41705) );
na02f80 g755747 ( .a(n_25112), .b(n_25058), .o(n_25111) );
in01f80 g778655 ( .a(n_2437), .o(n_3245) );
na02f80 g775159 ( .a(n_5953), .b(n_5914), .o(n_6047) );
in01f80 FE_OCPC1385_n_470 ( .a(n_470), .o(FE_OCPN1385_n_470) );
na02f80 g778398 ( .a(n_2457), .b(n_2463), .o(n_2464) );
no02f80 g754934 ( .a(FE_OCP_RBN2594_n_25181), .b(FE_OCPN3164_n_24117), .o(n_25239) );
na02f80 g743025 ( .a(n_37104), .b(n_37102), .o(n_37105) );
na02f80 g756937 ( .a(n_23672), .b(n_23810), .o(n_23724) );
na02f80 FE_RC_1793_0 ( .a(FE_RN_528_0), .b(n_34440), .o(n_34493) );
in01f80 newInst_514 ( .a(newNet_513), .o(newNet_514) );
in01f80 newInst_189 ( .a(newNet_188), .o(newNet_189) );
no02f80 g761454 ( .a(n_19609), .b(n_18778), .o(n_19714) );
na02f80 g744226 ( .a(n_36088), .b(n_36058), .o(n_36234) );
in01f80 FE_OCP_RBC2187_n_37686 ( .a(FE_OCP_RBN2186_n_37686), .o(FE_OCP_RBN2187_n_37686) );
in01f80 newInst_633 ( .a(newNet_632), .o(newNet_633) );
in01f80 newInst_499 ( .a(newNet_171), .o(newNet_499) );
no02f80 g750298 ( .a(n_30786), .b(n_30785), .o(n_30787) );
no02f80 g751885 ( .a(n_29308), .b(n_29071), .o(n_29072) );
no02f80 g738951 ( .a(n_41166), .b(n_41165), .o(n_41167) );
no03m80 FE_RC_3767_0 ( .a(n_10276), .b(n_10507), .c(n_10486), .o(n_10599) );
no02f80 FE_RC_2593_0 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_3_), .b(n_6804), .o(FE_RN_1073_0) );
no02f80 g775980 ( .a(n_5123), .b(n_4723), .o(n_5161) );
in01f80 FE_RC_1694_0 ( .a(n_25645), .o(FE_RN_468_0) );
oa22f80 g772041 ( .a(n_8900), .b(n_8166), .c(n_8852), .d(n_8167), .o(n_10122) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_24_ ( .ck(newNet_712), .d(n_46188), .o(delay_xor_ln21_unr6_stage3_stallmux_q_24_) );
na02f80 g741511 ( .a(n_38728), .b(n_38733), .o(n_38765) );
na02f80 g736583 ( .a(n_43335), .b(n_43385), .o(n_43450) );
no02f80 g765247 ( .a(n_15297), .b(n_15142), .o(n_15455) );
in01f80 FE_OCP_RBC2152_n_22822 ( .a(n_22822), .o(FE_OCP_RBN2152_n_22822) );
in01f80 g743002 ( .a(n_37357), .o(n_37160) );
in01f80 g739792 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_13_), .o(n_40493) );
na02f80 g765013 ( .a(n_15641), .b(n_15606), .o(n_15607) );
in01f80 FE_OCP_RBC1718_n_20090 ( .a(n_20090), .o(FE_OCP_RBN1718_n_20090) );
no02f80 g748076 ( .a(n_32841), .b(n_32840), .o(n_32842) );
in01f80 fopt783288 ( .a(n_44867), .o(n_44866) );
na02f80 g743194 ( .a(n_36918), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .o(n_36943) );
in01f80 newInst_826 ( .a(newNet_194), .o(newNet_826) );
ao12f80 g758965 ( .a(n_21356), .b(n_21540), .c(FE_OCP_RBN3683_FE_RN_770_0), .o(n_21609) );
in01f80 g774118 ( .a(n_7177), .o(n_7178) );
in01f80 g754626 ( .a(n_27366), .o(n_27536) );
in01f80 g742925 ( .a(n_37207), .o(n_37208) );
in01f80 FE_RC_3974_0 ( .a(n_29561), .o(FE_RN_1721_0) );
no02f80 g740767 ( .a(n_39294), .b(n_39216), .o(n_39450) );
in01f80 newInst_3263 ( .a(newNet_3262), .o(newNet_3263) );
ms00f80 cos_out_reg_23_ ( .ck(newNet_3716), .d(n_43869), .o(cos_out_23) );
ao22s80 FE_RC_3766_0 ( .a(n_14403), .b(n_14474), .c(n_14404), .d(n_14448), .o(n_14641) );
in01f80 FE_OCP_RBC2523_n_8951 ( .a(FE_OCP_RBN2522_n_8951), .o(FE_OCP_RBN2523_n_8951) );
na02f80 g741310 ( .a(FE_OCP_RBN2549_n_44944), .b(n_38873), .o(n_39260) );
in01f80 g766836 ( .a(n_13645), .o(n_13711) );
in01f80 FE_OCP_RBC2220_n_12888 ( .a(n_12888), .o(FE_OCP_RBN2220_n_12888) );
in01f80 g744677 ( .a(n_35288), .o(n_35289) );
oa12f80 g774125 ( .a(n_6675), .b(n_6674), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n_7364) );
no02f80 g749291 ( .a(n_30670), .b(n_30294), .o(n_30765) );
na02f80 g753077 ( .a(n_27126), .b(n_27157), .o(n_27190) );
no02f80 g746921 ( .a(FE_OCP_RBN3384_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_24_), .o(n_33231) );
in01f80 g738686 ( .a(n_41877), .o(n_41878) );
na02f80 g771204 ( .a(n_9424), .b(FE_OCP_RBN2643_FE_RN_1198_0), .o(n_9543) );
oa22f80 g742159 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37398), .c(n_44887), .d(n_37910), .o(n_38334) );
no02f80 g742241 ( .a(FE_OCP_RBN2240_n_44881), .b(n_37697), .o(n_38157) );
na02f80 g769106 ( .a(n_11673), .b(n_11649), .o(n_11806) );
oa12f80 g755382 ( .a(n_24763), .b(n_24762), .c(n_24761), .o(n_26468) );
in01f80 g765037 ( .a(n_15464), .o(n_15465) );
no02f80 g745584 ( .a(n_34297), .b(n_33426), .o(n_34316) );
na02f80 g772050 ( .a(n_8893), .b(n_8855), .o(n_8998) );
na02f80 g768498 ( .a(n_12338), .b(FE_OCPN1002_n_45660), .o(n_12384) );
no02f80 g767608 ( .a(n_13047), .b(n_13138), .o(n_13190) );
in01f80 g760748 ( .a(n_19635), .o(n_19636) );
in01f80 g778715 ( .a(n_2491), .o(n_2654) );
no02f80 g753278 ( .a(n_27167), .b(FE_OCP_RBN2909_n_26173), .o(n_27294) );
in01f80 g741649 ( .a(n_38587), .o(n_38598) );
in01f80 newInst_3538 ( .a(newNet_1248), .o(newNet_3538) );
na02f80 FE_RC_2291_0 ( .a(FE_RN_860_0), .b(n_45524), .o(FE_RN_861_0) );
no02f80 g753941 ( .a(FE_OCP_RBN2893_n_26152), .b(n_23466), .o(n_26223) );
ao12f80 g748360 ( .a(n_32749), .b(n_32748), .c(n_32747), .o(n_33415) );
in01f80 FE_OCP_RBC3844_FE_RN_1242_0 ( .a(FE_RN_1242_0), .o(FE_OCP_RBN3844_FE_RN_1242_0) );
in01f80 g743314 ( .a(n_36778), .o(n_36779) );
no02f80 g776412 ( .a(n_4381), .b(n_4328), .o(n_4472) );
na03f80 FE_RC_2549_0 ( .a(n_37368), .b(n_37142), .c(n_37369), .o(n_37401) );
in01f80 g751975 ( .a(n_28863), .o(n_28907) );
no02f80 g781342 ( .a(n_47), .b(n_46055), .o(n_86) );
in01f80 FE_OCPC3182_FE_OCP_RBN2831_n_10198 ( .a(FE_OCPN3181_FE_OCP_RBN2831_n_10198), .o(FE_OCPN3182_FE_OCP_RBN2831_n_10198) );
no02f80 g759528 ( .a(n_20768), .b(FE_OCP_RBN2664_n_20333), .o(n_20819) );
na02f80 g736894 ( .a(n_43486), .b(n_43184), .o(n_43587) );
in01f80 newInst_2080 ( .a(newNet_2079), .o(newNet_2080) );
ao12f80 g772351 ( .a(n_7466), .b(n_8407), .c(n_7501), .o(n_8504) );
no02f80 g741148 ( .a(n_39120), .b(FE_OCP_RBN2604_n_39126), .o(n_39186) );
no02f80 g738565 ( .a(n_41607), .b(n_41724), .o(n_41762) );
in01f80 newInst_1548 ( .a(newNet_1264), .o(newNet_1548) );
na02f80 g778389 ( .a(n_2511), .b(n_1835), .o(n_2626) );
ao12f80 g741462 ( .a(n_38768), .b(n_38767), .c(n_38766), .o(n_38794) );
in01f80 g773459 ( .a(n_7545), .o(n_7546) );
in01f80 g738198 ( .a(n_41991), .o(n_42423) );
no02f80 g745531 ( .a(n_34816), .b(n_34846), .o(n_34896) );
in01f80 newInst_918 ( .a(newNet_433), .o(newNet_918) );
no02f80 FE_RC_2689_0 ( .a(n_9012), .b(n_9190), .o(FE_RN_1126_0) );
in01f80 g775370 ( .a(FE_OCP_RBN2979_n_5656), .o(n_5703) );
no02f80 g774746 ( .a(n_6319), .b(n_6328), .o(n_6329) );
oa22f80 g774397 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_), .c(FE_OCPN895_n_6521), .d(n_6761), .o(n_6956) );
in01f80 FE_RC_625_0 ( .a(n_32553), .o(FE_RN_192_0) );
oa12f80 g740906 ( .a(n_39287), .b(n_39286), .c(n_39285), .o(n_39371) );
no02f80 g779407 ( .a(n_1537), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_), .o(n_1538) );
in01f80 g737945 ( .a(n_42341), .o(n_42342) );
in01f80 FE_OCP_RBC1216_n_20595 ( .a(n_20595), .o(FE_OCP_RBN1216_n_20595) );
na02f80 g777104 ( .a(n_3752), .b(n_3700), .o(n_3943) );
ao12f80 g779310 ( .a(n_1692), .b(n_1691), .c(n_1690), .o(n_2405) );
na02f80 g775774 ( .a(n_5332), .b(n_5145), .o(n_5410) );
in01f80 g769698 ( .a(n_11294), .o(n_11310) );
na02f80 g759919 ( .a(n_21051), .b(n_20156), .o(n_21253) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_28_ ( .ck(newNet_3027), .d(n_1066), .o(delay_add_ln22_unr2_stage2_stallmux_q_28_) );
no02f80 g768659 ( .a(n_12249), .b(n_12260), .o(n_12250) );
na02f80 g738417 ( .a(n_41632), .b(n_41631), .o(n_41633) );
na02f80 g759961 ( .a(n_20709), .b(n_20456), .o(n_20787) );
in01f80 g754956 ( .a(n_25904), .o(n_25977) );
in01f80 g770827 ( .a(n_10032), .o(n_10033) );
na02f80 FE_RC_3097_0 ( .a(FE_RN_1368_0), .b(FE_OCP_RBN3712_n_31466), .o(n_31548) );
in01f80 newInst_3342 ( .a(newNet_3341), .o(newNet_3342) );
oa12f80 g772456 ( .a(n_8302), .b(n_44351), .c(n_8303), .o(n_8381) );
in01f80 g776936 ( .a(n_4065), .o(n_4066) );
ao12f80 g764634 ( .a(n_15787), .b(n_16450), .c(n_15783), .o(n_16509) );
in01f80 g739182 ( .a(n_40894), .o(n_41206) );
ao22s80 g768378 ( .a(n_12481), .b(n_12315), .c(n_12450), .d(n_12314), .o(n_13510) );
na02f80 g750122 ( .a(FE_OCP_RBN3567_n_29857), .b(FE_OCP_RBN2236_n_29055), .o(n_30049) );
in01f80 newInst_2460 ( .a(newNet_2459), .o(newNet_2460) );
in01f80 newInst_660 ( .a(newNet_88), .o(newNet_660) );
ao12f80 g769018 ( .a(n_11420), .b(n_11434), .c(n_11454), .o(n_11535) );
na02f80 g764255 ( .a(n_16458), .b(n_16429), .o(n_16489) );
in01f80 FE_RC_1934_0 ( .a(n_18848), .o(FE_RN_615_0) );
na02f80 g763185 ( .a(n_17438), .b(n_17437), .o(n_17439) );
oa22f80 FE_RC_3250_0 ( .a(n_10615), .b(n_10661), .c(n_10616), .d(n_10660), .o(n_10784) );
in01f80 g779458 ( .a(n_1491), .o(n_1492) );
in01f80 g762695 ( .a(n_17947), .o(n_17948) );
no02f80 g741140 ( .a(n_39041), .b(n_39040), .o(n_39042) );
no02f80 g770837 ( .a(n_47260), .b(n_9930), .o(n_9947) );
in01f80 g758525 ( .a(n_21968), .o(n_21990) );
in01f80 FE_OCP_RBC2462_n_3076 ( .a(n_3076), .o(FE_OCP_RBN2462_n_3076) );
in01f80 FE_OCP_RBC2208_n_12907 ( .a(FE_OCP_RBN2207_n_12907), .o(FE_OCP_RBN2208_n_12907) );
na02f80 g771275 ( .a(n_9531), .b(n_9406), .o(n_9532) );
in01f80 FE_RC_3632_0 ( .a(FE_RN_1592_0), .o(n_24404) );
na02f80 g779320 ( .a(n_1639), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_), .o(n_1729) );
no02f80 g772730 ( .a(n_8259), .b(n_8258), .o(n_8300) );
ao22s80 FE_RC_568_0 ( .a(n_30640), .b(n_30866), .c(n_30621), .d(n_30865), .o(n_31046) );
in01f80 newInst_3564 ( .a(newNet_3563), .o(newNet_3564) );
in01f80 g757040 ( .a(n_23909), .o(n_23831) );
in01f80 FE_RC_3057_0 ( .a(n_26797), .o(FE_RN_1340_0) );
na02f80 g776999 ( .a(n_4128), .b(n_4059), .o(n_4198) );
no02f80 g772442 ( .a(n_8443), .b(n_8254), .o(n_8496) );
in01f80 newInst_581 ( .a(newNet_580), .o(newNet_581) );
in01f80 g771772 ( .a(n_9229), .o(n_9230) );
oa22f80 g769309 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .c(n_10812), .d(FE_OCPN1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_12442) );
oa12f80 g736639 ( .a(n_321), .b(n_43151), .c(FE_OFN5_n_43918), .o(n_43288) );
na02f80 g758232 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .o(n_22808) );
in01f80 g737516 ( .a(n_43121), .o(n_43494) );
no02f80 g764682 ( .a(n_15797), .b(n_14452), .o(n_16080) );
no02f80 g780691 ( .a(n_653), .b(n_652), .o(n_654) );
na02f80 g784605 ( .a(n_12686), .b(n_12406), .o(n_46933) );
in01f80 g758228 ( .a(n_22699), .o(n_22653) );
in01f80 drc784079 ( .a(n_45821), .o(n_45824) );
na02f80 g744995 ( .a(n_34797), .b(n_34338), .o(n_34880) );
in01f80 fopt783556 ( .a(n_45153), .o(n_45155) );
in01f80 newInst_1132 ( .a(newNet_756), .o(newNet_1132) );
in01f80 g774445 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_26_), .o(n_6631) );
na02f80 g738421 ( .a(n_41583), .b(n_41629), .o(n_41630) );
ao12f80 g766519 ( .a(n_46984), .b(n_14115), .c(n_12868), .o(n_14116) );
ao12f80 g756520 ( .a(n_23851), .b(n_23783), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n_23964) );
na02f80 g764782 ( .a(n_15595), .b(n_14419), .o(n_15628) );
no02f80 g755332 ( .a(n_24920), .b(n_24919), .o(n_24882) );
na02f80 g744756 ( .a(n_35200), .b(n_35141), .o(n_35221) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_21_ ( .ck(newNet_3316), .d(n_32255), .o(delay_add_ln22_unr20_stage8_stallmux_q_21_) );
na02f80 g749197 ( .a(n_30818), .b(FE_OCPN1410_n_27014), .o(n_30936) );
na02f80 g771947 ( .a(FE_OFN754_n_44461), .b(n_9544), .o(n_9693) );
in01f80 g780406 ( .a(n_851), .o(n_807) );
no02f80 g756641 ( .a(n_23518), .b(n_23556), .o(n_23797) );
in01f80 newInst_2246 ( .a(newNet_545), .o(newNet_2246) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_6_ ( .ck(newNet_548), .d(n_17224), .o(delay_xor_ln22_unr12_stage5_stallmux_q_6_) );
no02f80 g738531 ( .a(FE_OCP_RBN2312_n_41420), .b(n_41542), .o(n_41640) );
no02f80 g779035 ( .a(n_2063), .b(n_2062), .o(n_2064) );
in01f80 FE_OCPC1014_n_32820 ( .a(n_32820), .o(FE_OCPN1014_n_32820) );
na02f80 g736688 ( .a(n_43401), .b(n_43350), .o(n_43437) );
ao12f80 g773953 ( .a(n_7254), .b(n_7217), .c(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .o(n_7441) );
in01f80 newInst_3029 ( .a(newNet_3028), .o(newNet_3029) );
na02f80 g743041 ( .a(n_37106), .b(n_37148), .o(n_37496) );
in01f80 fopt782740 ( .a(n_17688), .o(n_44150) );
no02f80 g738031 ( .a(n_42148), .b(n_42158), .o(n_42159) );
oa22f80 FE_RC_1490_0 ( .a(n_24350), .b(n_27771), .c(n_27845), .d(n_27744), .o(n_27819) );
oa22f80 FE_RC_1488_0 ( .a(n_24059), .b(n_27728), .c(n_27796), .d(n_27706), .o(n_27750) );
in01f80 g773571 ( .a(n_8444), .o(n_7458) );
in01f80 g766503 ( .a(n_14028), .o(n_14029) );
in01f80 fopt783271 ( .a(n_33873), .o(n_44842) );
in01f80 g741251 ( .a(n_39026), .o(n_39027) );
na02f80 g751603 ( .a(FE_OCP_RBN3404_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n_28773) );
na02f80 g773895 ( .a(n_6941), .b(n_6748), .o(n_6997) );
ao12f80 g743753 ( .a(n_35754), .b(n_36109), .c(n_35873), .o(n_36275) );
no02f80 g776649 ( .a(n_4229), .b(n_4228), .o(n_4557) );
no02f80 g763123 ( .a(n_17251), .b(n_17225), .o(n_17515) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_26_ ( .ck(newNet_3216), .d(n_36581), .o(delay_add_ln22_unr23_stage9_stallmux_q_26_) );
in01f80 g761009 ( .a(n_19323), .o(n_19324) );
no02f80 g740757 ( .a(n_39384), .b(n_39078), .o(n_39411) );
no02f80 g761831 ( .a(n_18481), .b(n_18479), .o(n_18482) );
in01f80 g748609 ( .a(n_31336), .o(n_31383) );
no02f80 g776006 ( .a(n_4749), .b(n_4769), .o(n_4936) );
in01f80 g769133 ( .a(n_11739), .o(n_11740) );
ao12f80 g773054 ( .a(n_7629), .b(n_7636), .c(n_7628), .o(n_8021) );
na02f80 g761743 ( .a(n_18709), .b(n_18684), .o(n_18855) );
no02f80 FE_RC_3229_0 ( .a(FE_RN_1430_0), .b(FE_OCP_RBN3578_n_8774), .o(FE_RN_1432_0) );
ms00f80 sin_out_reg_27_ ( .ck(newNet_39), .d(n_43917), .o(sin_out_27) );
na02f80 g758319 ( .a(n_22249), .b(FE_OCP_RBN3219_n_21358), .o(n_22293) );
no02f80 g770947 ( .a(n_9748), .b(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .o(n_9909) );
in01f80 FE_RC_2738_0 ( .a(FE_RN_1161_0), .o(n_9570) );
no02f80 FE_RC_2105_0 ( .a(n_20372), .b(FE_OCP_RBN1695_n_19206), .o(FE_RN_727_0) );
oa12f80 g758910 ( .a(n_21569), .b(n_21642), .c(n_21487), .o(n_21705) );
in01f80 newInst_751 ( .a(newNet_750), .o(newNet_751) );
na02f80 g779737 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .o(n_1613) );
in01f80 g762122 ( .a(n_18205), .o(n_18206) );
na02f80 g781063 ( .a(sin_out_29), .b(FE_OFN4_n_43918), .o(n_333) );
no02f80 g748313 ( .a(n_31555), .b(n_31599), .o(n_31607) );
in01f80 g777959 ( .a(n_3114), .o(n_3083) );
in01f80 newInst_1110 ( .a(newNet_1109), .o(newNet_1110) );
na02f80 g780524 ( .a(n_842), .b(n_776), .o(n_825) );
in01f80 g742537 ( .a(n_37597), .o(n_37760) );
na02f80 g767769 ( .a(n_13317), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_), .o(n_13421) );
in01f80 g768489 ( .a(n_12423), .o(n_12457) );
ao12f80 g752295 ( .a(n_27999), .b(FE_OCP_RBN2126_n_44734), .c(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .o(n_28028) );
in01f80 g737896 ( .a(n_42247), .o(n_42248) );
na02f80 g739718 ( .a(n_40539), .b(n_40437), .o(n_40561) );
no02f80 g758887 ( .a(n_21661), .b(n_21577), .o(n_21578) );
in01f80 g743700 ( .a(n_36408), .o(n_36409) );
no02f80 g742424 ( .a(n_37720), .b(n_37670), .o(n_37721) );
ao22s80 FE_RC_3835_0 ( .a(n_35946), .b(n_36431), .c(n_35945), .d(n_36445), .o(n_36489) );
in01f80 newInst_2912 ( .a(newNet_2911), .o(newNet_2912) );
oa12f80 g748495 ( .a(n_31494), .b(n_31589), .c(FE_OCP_RBN2972_n_31239), .o(n_31718) );
ao12f80 g749749 ( .a(n_31092), .b(n_31091), .c(n_31090), .o(n_31481) );
na02f80 g743622 ( .a(n_36381), .b(n_35899), .o(n_36400) );
na02f80 FE_RC_2597_0 ( .a(n_2878), .b(n_2877), .o(FE_RN_1076_0) );
ao12f80 g746989 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_13_), .c(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n_33380) );
na02f80 g753402 ( .a(n_27010), .b(n_27009), .o(n_27057) );
oa12f80 g736428 ( .a(n_336), .b(n_43760), .c(n_43918), .o(n_43817) );
in01f80 FE_RC_4168_0 ( .a(n_18519), .o(FE_RN_1817_0) );
in01f80 g742972 ( .a(n_36974), .o(n_37071) );
in01f80 g749004 ( .a(n_31099), .o(n_31100) );
in01f80 newInst_831 ( .a(newNet_479), .o(newNet_831) );
in01f80 g743823 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n_35989) );
oa12f80 g772942 ( .a(n_7963), .b(n_8000), .c(n_8058), .o(n_8088) );
no02f80 g780876 ( .a(n_377), .b(n_393), .o(n_416) );
na02f80 FE_RC_2758_0 ( .a(FE_RN_1173_0), .b(n_18602), .o(n_18650) );
in01f80 g3 ( .a(n_44030), .o(n_44031) );
in01f80 newInst_90 ( .a(newNet_89), .o(newNet_90) );
in01f80 g761629 ( .a(n_18918), .o(n_18973) );
no02f80 g779626 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_22_), .o(n_1998) );
in01f80 FE_OCP_RBC3556_n_44575 ( .a(FE_OCP_RBN3553_n_44575), .o(FE_OCP_RBN3556_n_44575) );
no02f80 g754557 ( .a(n_26550), .b(n_26549), .o(n_26574) );
in01f80 FE_RC_2194_0 ( .a(n_31463), .o(FE_RN_787_0) );
in01f80 g762884 ( .a(n_17794), .o(n_17795) );
na02f80 g741182 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39324), .o(n_39425) );
na02f80 g776432 ( .a(n_4525), .b(n_4255), .o(n_4593) );
in01f80 FE_RC_3459_0 ( .a(FE_RN_1487_0), .o(FE_RN_1486_0) );
in01f80 g770568 ( .a(n_10314), .o(n_10315) );
in01f80 g741565 ( .a(n_38673), .o(n_38674) );
oa12f80 g758631 ( .a(n_21680), .b(n_21811), .c(n_21741), .o(n_21900) );
no02f80 g772913 ( .a(n_7901), .b(n_7926), .o(n_8051) );
oa22f80 FE_RC_3446_0 ( .a(n_23880), .b(n_24489), .c(n_23879), .d(n_24490), .o(n_24612) );
na02f80 g772230 ( .a(n_8611), .b(n_7610), .o(n_8668) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_9_ ( .ck(newNet_388), .d(n_32569), .o(delay_xor_ln22_unr21_stage8_stallmux_q_9_) );
ao22s80 g780854 ( .a(n_521), .b(n_241), .c(n_420), .d(n_235), .o(n_604) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_4_ ( .ck(newNet_1931), .d(n_36829), .o(delay_sub_ln21_unr24_stage9_stallmux_q_4_) );
no02f80 g777825 ( .a(n_3244), .b(n_3269), .o(n_3328) );
na02f80 g781038 ( .a(sin_out_14), .b(FE_OFN3_n_43918), .o(n_312) );
na04m80 g773943 ( .a(n_6831), .b(n_6801), .c(n_6802), .d(n_6645), .o(n_6883) );
oa12f80 g754875 ( .a(n_25885), .b(n_25884), .c(n_25883), .o(n_26604) );
na02f80 g777269 ( .a(n_3545), .b(n_3029), .o(n_3679) );
no02f80 g736955 ( .a(FE_OCPN912_n_43022), .b(n_46938), .o(n_43362) );
in01f80 newInst_1104 ( .a(newNet_293), .o(newNet_1104) );
in01f80 g765180 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_2_), .o(n_17229) );
oa12f80 g774946 ( .a(n_6007), .b(n_6118), .c(n_5982), .o(n_6181) );
in01f80 g776002 ( .a(n_5196), .o(n_5273) );
oa22f80 g759817 ( .a(n_21714), .b(n_21597), .c(n_21691), .d(n_21562), .o(n_21855) );
in01f80 newInst_2091 ( .a(newNet_2090), .o(newNet_2091) );
in01f80 FE_OCP_RBC1091_n_45224 ( .a(FE_OCP_RBN3269_n_45224), .o(FE_OCP_RBN1091_n_45224) );
in01f80 newInst_251 ( .a(newNet_250), .o(newNet_251) );
in01f80 newInst_194 ( .a(newNet_193), .o(newNet_194) );
na02f80 g753590 ( .a(n_26755), .b(n_26754), .o(n_26776) );
na02f80 g774312 ( .a(n_6518), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6607) );
no02f80 g738168 ( .a(n_42033), .b(n_42032), .o(n_42034) );
in01f80 newInst_1762 ( .a(newNet_907), .o(newNet_1762) );
in01f80 g762978 ( .a(n_17592), .o(n_17593) );
ao22s80 FE_RC_3757_0 ( .a(n_6616), .b(n_6635), .c(FE_OCP_RBN2110_n_6616), .d(n_6636), .o(n_6798) );
in01f80 FE_OCP_RBC3033_n_43000 ( .a(n_43000), .o(FE_OCP_RBN3033_n_43000) );
in01f80 FE_OCPC946_n_1780 ( .a(FE_OCPN945_n_1780), .o(FE_OCPN946_n_1780) );
in01f80 FE_OCP_RBC1991_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_ ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(FE_OCP_RBN1991_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
na02f80 g781322 ( .a(n_46055), .b(beta_15), .o(n_42) );
no02f80 g768120 ( .a(n_12589), .b(n_12400), .o(n_12616) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_22_ ( .ck(newNet_3139), .d(n_40512), .o(delay_add_ln22_unr27_stage10_stallmux_q_22_) );
no02f80 FE_RC_3058_0 ( .a(FE_RN_1339_0), .b(FE_RN_1340_0), .o(FE_RN_1341_0) );
no02f80 g777372 ( .a(n_5494), .b(n_4797), .o(n_4863) );
in01f80 g771241 ( .a(n_9502), .o(n_9565) );
na02f80 g780883 ( .a(n_457), .b(n_493), .o(n_497) );
in01f80 newInst_2654 ( .a(newNet_2653), .o(newNet_2654) );
in01f80 g771667 ( .a(n_9264), .o(n_9265) );
na02f80 g757653 ( .a(n_22632), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n_22633) );
in01f80 fopt782751 ( .a(n_38788), .o(n_44166) );
oa22f80 FE_RC_1422_0 ( .a(n_30584), .b(n_30747), .c(n_30651), .d(n_27014), .o(n_30769) );
na02f80 g777844 ( .a(n_3204), .b(n_2385), .o(n_3206) );
in01f80 newInst_1925 ( .a(newNet_1450), .o(newNet_1925) );
no02f80 g781117 ( .a(n_229), .b(n_228), .o(n_230) );
na02f80 g775096 ( .a(n_6036), .b(n_5889), .o(n_6121) );
no02f80 FE_RC_3596_0 ( .a(n_13310), .b(FE_RN_1569_0), .o(FE_RN_1570_0) );
na02f80 FE_RC_3073_0 ( .a(FE_RN_1351_0), .b(FE_RN_1349_0), .o(FE_RN_1352_0) );
in01f80 g761175 ( .a(n_19641), .o(n_20369) );
in01f80 FE_RC_2938_0 ( .a(n_29442), .o(FE_RN_1282_0) );
no02f80 g762095 ( .a(n_18266), .b(delay_add_ln22_unr11_stage5_stallmux_q_19_), .o(n_18278) );
in01f80 newInst_1139 ( .a(newNet_1138), .o(newNet_1139) );
in01f80 g779444 ( .a(n_1474), .o(n_1475) );
no02f80 g777183 ( .a(n_5147), .b(n_5090), .o(n_5174) );
na02f80 g772023 ( .a(FE_OCP_RBN2518_n_8762), .b(n_8561), .o(n_8798) );
oa12f80 g738279 ( .a(n_41866), .b(n_41865), .c(n_41864), .o(n_42562) );
oa12f80 g762910 ( .a(n_17988), .b(n_17987), .c(n_17986), .o(n_18064) );
oa12f80 g760049 ( .a(n_20254), .b(n_21050), .c(n_20218), .o(n_21138) );
in01f80 g747994 ( .a(n_32109), .o(n_32110) );
in01f80 FE_RC_3514_0 ( .a(FE_RN_1518_0), .o(FE_OCPN988_n_28353) );
in01f80 FE_OCP_RBC1697_n_19206 ( .a(FE_OCP_RBN1696_n_19206), .o(FE_OCP_RBN1697_n_19206) );
no02f80 g750853 ( .a(n_29137), .b(FE_OCP_RBN1152_n_29053), .o(n_29180) );
na02f80 FE_RC_2052_0 ( .a(FE_RN_688_0), .b(FE_RN_692_0), .o(FE_RN_693_0) );
na02f80 g741988 ( .a(n_37914), .b(n_37981), .o(n_37982) );
in01f80 g755248 ( .a(n_24989), .o(n_25016) );
no02f80 g743113 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .o(n_37108) );
in01f80 newInst_3134 ( .a(newNet_3133), .o(newNet_3134) );
na02f80 g755735 ( .a(n_25112), .b(n_25089), .o(n_25113) );
na02f80 g753989 ( .a(n_26976), .b(n_26552), .o(n_27003) );
oa12f80 g751859 ( .a(n_28222), .b(n_28221), .c(n_28220), .o(n_28223) );
in01f80 g774932 ( .a(n_6259), .o(n_6260) );
in01f80 g752260 ( .a(n_27939), .o(n_27940) );
na02f80 g738914 ( .a(n_41195), .b(n_41014), .o(n_41261) );
in01f80 newInst_2536 ( .a(newNet_2535), .o(newNet_2536) );
oa22f80 g762065 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_31_), .c(FE_OCP_RBN2205_n_18242), .d(n_17852), .o(n_18669) );
ao22s80 FE_RC_1199_0 ( .a(n_15369), .b(n_15906), .c(n_15370), .d(n_15820), .o(n_16084) );
in01f80 g756612 ( .a(n_23708), .o(n_23765) );
no02f80 g741018 ( .a(n_38931), .b(n_38870), .o(n_39015) );
in01f80 g741782 ( .a(n_38474), .o(n_38453) );
in01f80 newInst_3162 ( .a(newNet_3161), .o(newNet_3162) );
in01f80 g770397 ( .a(n_10405), .o(n_10445) );
oa12f80 g746641 ( .a(n_32988), .b(n_33204), .c(n_32954), .o(n_33254) );
in01f80 newInst_3660 ( .a(newNet_3659), .o(newNet_3660) );
no02f80 g781296 ( .a(beta_31), .b(beta_13), .o(n_82) );
in01f80 FE_OCPC1401_n_9642 ( .a(n_9642), .o(FE_OCPN1401_n_9642) );
oa22f80 g746867 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .c(FE_OCP_RBN2171_n_32892), .d(n_32362), .o(n_33470) );
in01f80 g777583 ( .a(n_3638), .o(n_3698) );
na02f80 g746830 ( .a(n_33079), .b(n_33078), .o(n_33100) );
na02f80 g779163 ( .a(n_1911), .b(n_1758), .o(n_1948) );
in01f80 g775322 ( .a(n_5971), .o(n_5935) );
in01f80 g772470 ( .a(n_10214), .o(n_8514) );
ao12f80 g761755 ( .a(n_19233), .b(n_19232), .c(n_19231), .o(n_19793) );
in01f80 g772937 ( .a(n_7931), .o(n_7932) );
in01f80 g754270 ( .a(n_25940), .o(n_25974) );
no02f80 g742071 ( .a(FE_OCP_RBN3446_n_37945), .b(n_37575), .o(n_38106) );
ao22s80 g769573 ( .a(n_11383), .b(n_11360), .c(n_11400), .d(n_11359), .o(n_11495) );
oa22f80 g779859 ( .a(n_44652), .b(n_1163), .c(n_44623), .d(n_1151), .o(n_1315) );
oa22f80 FE_RC_1210_0 ( .a(n_13321), .b(n_13838), .c(n_13320), .d(n_13812), .o(n_13960) );
in01f80 g745313 ( .a(n_35992), .o(n_35993) );
in01f80 newInst_3241 ( .a(newNet_3240), .o(newNet_3241) );
no02f80 g769567 ( .a(n_11327), .b(n_11279), .o(n_11336) );
in01f80 newInst_3718 ( .a(newNet_3717), .o(newNet_3718) );
in01f80 FE_OCPC850_n_2306 ( .a(FE_OCPN849_n_2306), .o(FE_OCPN850_n_2306) );
no02f80 FE_RC_2347_0 ( .a(FE_RN_900_0), .b(n_33004), .o(n_33048) );
in01f80 g736779 ( .a(n_43396), .o(n_43397) );
in01f80 FE_OCPC3784_FE_OCP_RBN2831_n_10198 ( .a(FE_OCP_RBN2831_n_10198), .o(FE_OCPN3784_FE_OCP_RBN2831_n_10198) );
na02f80 g773495 ( .a(n_7445), .b(delay_add_ln22_unr5_stage3_stallmux_q_23_), .o(n_7465) );
na02f80 g748768 ( .a(n_31352), .b(n_31298), .o(n_31375) );
no02f80 g772004 ( .a(n_44568), .b(FE_OCP_RBN3559_n_8809), .o(n_8925) );
na02f80 g746595 ( .a(n_34612), .b(n_34613), .o(n_34699) );
oa22f80 g748858 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .c(n_32034), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32806) );
no02f80 g743060 ( .a(n_37144), .b(n_37029), .o(n_37173) );
in01f80 newInst_2557 ( .a(newNet_2556), .o(newNet_2557) );
ao22s80 g743858 ( .a(n_46250), .b(n_36851), .c(n_36980), .d(n_46246), .o(n_37224) );
na02f80 g750465 ( .a(n_30552), .b(n_30520), .o(n_30521) );
oa12f80 g751204 ( .a(n_29944), .b(n_29999), .c(n_29509), .o(n_29990) );
in01f80 g771384 ( .a(n_9446), .o(n_9464) );
in01f80 FE_OCP_RBC3449_n_37945 ( .a(FE_OCP_RBN3445_n_37945), .o(FE_OCP_RBN3449_n_37945) );
in01f80 newInst_2020 ( .a(newNet_1024), .o(newNet_2020) );
na02f80 g767435 ( .a(n_13338), .b(n_13400), .o(n_13339) );
in01f80 g762045 ( .a(n_18539), .o(n_18540) );
in01f80 g772807 ( .a(n_8159), .o(n_8170) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_2_ ( .ck(newNet_1081), .d(n_9518), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_) );
in01f80 g753366 ( .a(n_27287), .o(n_27377) );
na02f80 g767789 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n_12930) );
in01f80 g754493 ( .a(n_26772), .o(n_26773) );
oa22f80 g740331 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39969), .c(FE_OCP_RBN3021_n_39942), .d(n_39519), .o(n_40394) );
no02f80 g736394 ( .a(n_43747), .b(n_43434), .o(n_43775) );
in01f80 g776535 ( .a(n_4485), .o(n_4486) );
na02f80 g754870 ( .a(n_25301), .b(n_25357), .o(n_25426) );
in01f80 FE_RC_3300_0 ( .a(FE_RN_1452_0), .o(FE_RN_1451_0) );
in01f80 FE_OCPC867_n_45697 ( .a(FE_OCPN866_n_45697), .o(FE_OCPN867_n_45697) );
oa12f80 g757783 ( .a(n_23087), .b(n_23010), .c(n_22697), .o(n_23155) );
na02f80 g776354 ( .a(n_4634), .b(n_4186), .o(n_4703) );
no02f80 g772744 ( .a(n_8127), .b(n_46991), .o(n_8165) );
in01f80 g766646 ( .a(n_13947), .o(n_13981) );
in01f80 g741176 ( .a(n_39242), .o(n_39243) );
in01f80 FE_OCP_RBC3057_n_36506 ( .a(n_36506), .o(FE_OCP_RBN3057_n_36506) );
oa12f80 g754736 ( .a(n_25287), .b(n_26161), .c(n_25312), .o(n_26238) );
na02f80 g756542 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23883) );
in01f80 g750877 ( .a(n_29062), .o(n_29292) );
oa12f80 g742580 ( .a(n_37430), .b(n_37429), .c(n_37428), .o(n_37493) );
no02f80 g740407 ( .a(FE_OCP_RBN3022_n_39942), .b(n_39605), .o(n_40303) );
in01f80 g759268 ( .a(n_20979), .o(n_20978) );
in01f80 FE_RC_1111_0 ( .a(FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_RN_334_0) );
oa12f80 g771410 ( .a(n_9607), .b(n_9606), .c(n_9605), .o(n_9782) );
na02f80 g758291 ( .a(FE_OCPN992_n_22249), .b(n_20688), .o(n_22372) );
in01f80 g761883 ( .a(n_18433), .o(n_18468) );
oa12f80 g773843 ( .a(n_7112), .b(n_7111), .c(n_7110), .o(n_7163) );
no02f80 g771840 ( .a(n_9771), .b(n_9734), .o(n_10686) );
in01f80 newInst_1458 ( .a(newNet_1457), .o(newNet_1458) );
no02f80 g753087 ( .a(FE_OCPN3186_FE_OCP_RBN1140_n_25816), .b(n_27124), .o(n_27156) );
in01f80 newInst_3003 ( .a(newNet_2718), .o(newNet_3003) );
in01f80 g769884 ( .a(n_11177), .o(n_11151) );
oa12f80 g760522 ( .a(n_19897), .b(n_19896), .c(n_19895), .o(n_21728) );
no02f80 g759610 ( .a(n_20646), .b(n_20289), .o(n_20728) );
in01f80 g750269 ( .a(n_30840), .o(n_30923) );
in01f80 FE_OCPC3789_n_15708 ( .a(FE_OCPN3788_n_15708), .o(FE_OCPN3789_n_15708) );
in01f80 g754374 ( .a(n_25889), .o(n_25907) );
ao12f80 g752705 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .b(n_27997), .c(n_27988), .o(n_27998) );
oa22f80 FE_RC_1196_0 ( .a(FE_OCP_RBN2395_n_8288), .b(n_8602), .c(FE_OCP_RBN2394_n_8288), .d(n_8601), .o(n_8753) );
in01f80 newInst_3277 ( .a(newNet_3276), .o(newNet_3277) );
na02f80 g751633 ( .a(n_28422), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .o(n_28465) );
in01f80 newInst_1887 ( .a(newNet_1886), .o(newNet_1887) );
ao12f80 g742684 ( .a(n_37107), .b(n_37407), .c(n_37148), .o(n_37501) );
na02f80 g767074 ( .a(n_13598), .b(n_12586), .o(n_13669) );
ao22s80 FE_RC_292_0 ( .a(n_45024), .b(n_21216), .c(n_45023), .d(n_21203), .o(n_21390) );
in01f80 FE_RC_3660_0 ( .a(FE_RN_1605_0), .o(FE_RN_1607_0) );
ao12f80 g757102 ( .a(n_23114), .b(n_44068), .c(delay_xor_ln22_unr15_stage6_stallmux_q_15_), .o(n_23142) );
na02f80 g774843 ( .a(n_6343), .b(n_6302), .o(n_6435) );
in01f80 g747437 ( .a(n_33533), .o(n_33574) );
in01f80 newInst_2583 ( .a(newNet_2582), .o(newNet_2583) );
in01f80 g773806 ( .a(n_7201), .o(n_7202) );
in01f80 FE_OFC832_n_18287 ( .a(n_18287), .o(FE_OFN832_n_18287) );
no02f80 g746345 ( .a(n_33561), .b(n_33560), .o(n_33562) );
oa12f80 g775317 ( .a(n_5530), .b(n_5554), .c(n_5365), .o(n_5674) );
na02f80 g772624 ( .a(n_8244), .b(n_8250), .o(n_8332) );
in01f80 g739733 ( .a(n_40501), .o(n_40502) );
in01f80 newInst_1836 ( .a(newNet_1835), .o(newNet_1836) );
oa12f80 g765111 ( .a(FE_OFN764_n_15670), .b(n_16100), .c(n_16099), .o(n_16133) );
in01f80 g740931 ( .a(n_39113), .o(n_39146) );
no02f80 g774510 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n_6815) );
in01f80 FE_RC_650_0 ( .a(n_6932), .o(FE_RN_207_0) );
oa12f80 g741826 ( .a(n_38414), .b(n_38413), .c(n_38412), .o(n_38884) );
no02f80 g743016 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_27_), .o(n_36998) );
no02f80 g774018 ( .a(n_6946), .b(n_6945), .o(n_6947) );
na02f80 g783823 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_2_), .b(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n_45507) );
in01f80 newInst_868 ( .a(newNet_867), .o(newNet_868) );
no02f80 g760417 ( .a(n_20076), .b(n_20265), .o(n_20126) );
no02f80 g760318 ( .a(n_20238), .b(n_20225), .o(n_20325) );
no02f80 g756395 ( .a(n_24014), .b(n_24011), .o(n_24013) );
na02f80 g748816 ( .a(n_32485), .b(n_32415), .o(n_32530) );
no02f80 g774496 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .o(n_6877) );
ao12f80 g764474 ( .a(n_16180), .b(n_16179), .c(n_16107), .o(n_16316) );
oa12f80 g761944 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n_18431) );
in01f80 g773218 ( .a(n_7960), .o(n_7961) );
na02f80 g762238 ( .a(n_18186), .b(n_18213), .o(n_18238) );
in01f80 g752755 ( .a(n_27104), .o(n_27128) );
na02f80 g754038 ( .a(n_26204), .b(n_26149), .o(n_26245) );
in01f80 g746890 ( .a(n_33107), .o(n_33058) );
in01f80 g743137 ( .a(n_36983), .o(n_36984) );
in01f80 g767315 ( .a(n_13430), .o(n_13431) );
na02f80 g750731 ( .a(n_29327), .b(n_25738), .o(n_29270) );
na02f80 g749942 ( .a(n_30051), .b(FE_OCP_RBN2236_n_29055), .o(n_30078) );
in01f80 FE_OCP_RBC3415_n_12739 ( .a(n_12739), .o(FE_OCP_RBN3415_n_12739) );
oa12f80 g775566 ( .a(n_5216), .b(n_5551), .c(n_5153), .o(n_5624) );
in01f80 g770195 ( .a(n_10799), .o(n_10885) );
no02f80 FE_RC_2504_0 ( .a(FE_RN_1016_0), .b(n_8215), .o(n_8283) );
na02f80 g780462 ( .a(FE_OFN759_n_45813), .b(FE_OFN50_n_1045), .o(n_815) );
oa12f80 g756885 ( .a(n_23743), .b(n_23955), .c(n_23954), .o(n_23988) );
no02f80 g750330 ( .a(n_29681), .b(FE_OCP_RBN2445_n_29684), .o(n_29717) );
oa12f80 g769831 ( .a(n_10953), .b(n_10971), .c(n_10941), .o(n_11113) );
no02f80 g771827 ( .a(n_9770), .b(n_9828), .o(n_9829) );
in01f80 newInst_3071 ( .a(newNet_3070), .o(newNet_3071) );
na02f80 g748810 ( .a(n_32450), .b(n_32412), .o(n_33042) );
na02f80 g776232 ( .a(n_4626), .b(n_4625), .o(n_4657) );
no02f80 FE_RC_1641_0 ( .a(FE_RN_458_0), .b(n_23068), .o(n_23189) );
oa22f80 g784567 ( .a(FE_OFN801_n_46285), .b(n_11369), .c(FE_OCP_RBN3044_n_46337), .d(n_11338), .o(n_46388) );
na02f80 g773984 ( .a(n_6900), .b(n_6899), .o(n_6901) );
in01f80 g757663 ( .a(n_23242), .o(n_23243) );
in01f80 newInst_2681 ( .a(newNet_412), .o(newNet_2681) );
no02f80 g772847 ( .a(n_7822), .b(n_7379), .o(n_7903) );
no02f80 g780901 ( .a(n_357), .b(n_501), .o(n_358) );
no02f80 g760894 ( .a(n_19283), .b(n_19335), .o(n_19434) );
na02f80 g773182 ( .a(FE_OCP_RBN2229_n_7598), .b(n_7925), .o(n_7701) );
in01f80 g741046 ( .a(n_39077), .o(n_39078) );
ao12f80 g779492 ( .a(n_1861), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_17_), .o(n_1876) );
no02f80 g752729 ( .a(n_27549), .b(n_27548), .o(n_27550) );
in01f80 g744761 ( .a(n_36498), .o(n_36499) );
no02f80 g754229 ( .a(n_25931), .b(n_23254), .o(n_26128) );
in01f80 g748353 ( .a(n_31912), .o(n_31913) );
oa12f80 g775677 ( .a(n_4739), .b(n_5432), .c(n_4598), .o(n_5552) );
na02f80 g769975 ( .a(n_11008), .b(n_10801), .o(n_11032) );
no02f80 g765245 ( .a(n_15491), .b(n_15519), .o(n_15635) );
no02f80 g768537 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_16_), .o(n_12370) );
oa22f80 g771315 ( .a(n_9137), .b(n_9178), .c(n_9177), .d(n_9138), .o(n_9411) );
na02f80 g753329 ( .a(n_27057), .b(n_27025), .o(n_27071) );
in01f80 newInst_805 ( .a(newNet_804), .o(newNet_805) );
no02f80 g758987 ( .a(n_21202), .b(n_21239), .o(n_21289) );
in01f80 newInst_2717 ( .a(newNet_2716), .o(newNet_2717) );
in01f80 g777567 ( .a(n_3938), .o(n_4046) );
ao12f80 g775789 ( .a(n_4975), .b(n_4916), .c(n_5026), .o(n_5084) );
in01f80 FE_OCP_RBC2513_n_8533 ( .a(n_8533), .o(FE_OCP_RBN2513_n_8533) );
no02f80 g762246 ( .a(n_18453), .b(n_18585), .o(n_18586) );
in01f80 newInst_114 ( .a(newNet_113), .o(newNet_114) );
oa12f80 g750031 ( .a(n_30953), .b(n_30952), .c(n_30951), .o(n_31038) );
no02f80 g769360 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_), .o(n_11896) );
no02f80 g768922 ( .a(FE_OCP_RBN2123_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_10_), .o(n_11888) );
no02f80 g766056 ( .a(n_14645), .b(n_14376), .o(n_14647) );
in01f80 g762312 ( .a(n_18078), .o(n_18079) );
in01f80 g759247 ( .a(n_21218), .o(n_21264) );
na02f80 g758316 ( .a(FE_OCP_RBN1846_n_22068), .b(FE_OCP_RBN1378_n_20889), .o(n_22149) );
ao12f80 g763953 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_8_), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n_17426) );
in01f80 newInst_3107 ( .a(newNet_3106), .o(newNet_3107) );
in01f80 g767247 ( .a(n_13623), .o(n_13624) );
no02f80 g752944 ( .a(n_27722), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .o(n_27763) );
in01f80 g774728 ( .a(n_6371), .o(n_6380) );
no02f80 g745364 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35720), .o(n_35937) );
na02f80 g749038 ( .a(n_31123), .b(n_31122), .o(n_31124) );
in01f80 newInst_1949 ( .a(newNet_1948), .o(newNet_1949) );
in01f80 FE_OCP_RBC2446_n_29684 ( .a(n_29684), .o(FE_OCP_RBN2446_n_29684) );
no02f80 g757300 ( .a(n_44066), .b(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .o(n_23308) );
na02f80 g779230 ( .a(n_1812), .b(n_1555), .o(n_1862) );
no02f80 g764417 ( .a(n_16095), .b(n_14420), .o(n_16236) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_4_ ( .ck(newNet_2443), .d(n_31397), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_) );
in01f80 FE_OCPC1766_n_33447 ( .a(FE_OCPN1765_n_33447), .o(FE_OCPN1766_n_33447) );
no02f80 g769057 ( .a(n_11594), .b(n_45224), .o(n_11691) );
in01f80 FE_OCP_RBC1170_n_13756 ( .a(FE_OCP_RBN3478_n_13756), .o(FE_OCP_RBN1170_n_13756) );
in01f80 g751546 ( .a(n_28474), .o(n_28451) );
no02f80 g774001 ( .a(n_6752), .b(n_6609), .o(n_6841) );
in01f80 g753546 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n_27453) );
na02f80 g765797 ( .a(n_14926), .b(n_14929), .o(n_14976) );
in01f80 FE_OCP_RBC2234_n_33648 ( .a(n_33648), .o(FE_OCP_RBN2234_n_33648) );
in01f80 newInst_2427 ( .a(newNet_2426), .o(newNet_2427) );
in01f80 g777235 ( .a(n_3686), .o(n_3687) );
no02f80 g756717 ( .a(n_23502), .b(delay_add_ln22_unr14_stage6_stallmux_q_14_), .o(n_23556) );
in01f80 FE_OCP_RBC3471_n_7886 ( .a(FE_OCP_RBN3469_n_7886), .o(FE_OCP_RBN3471_n_7886) );
na02f80 g748295 ( .a(n_31683), .b(n_31657), .o(n_31684) );
no02f80 g776797 ( .a(n_4281), .b(n_4280), .o(n_4446) );
na02f80 g749192 ( .a(n_30711), .b(FE_OCPN1410_n_27014), .o(n_30749) );
na02f80 g750951 ( .a(n_30039), .b(n_29821), .o(n_30105) );
in01f80 FE_OCP_RBC3727_FE_RN_1787_0 ( .a(FE_RN_1787_0), .o(FE_OCP_RBN3727_FE_RN_1787_0) );
na02f80 g738081 ( .a(n_42096), .b(n_42095), .o(n_42097) );
na02f80 g746487 ( .a(n_34529), .b(n_34499), .o(n_34553) );
no02f80 g774032 ( .a(n_6776), .b(n_6594), .o(n_6840) );
na02f80 g756841 ( .a(n_23362), .b(n_23350), .o(n_23424) );
in01f80 newInst_477 ( .a(newNet_476), .o(newNet_477) );
no02f80 g748889 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_), .o(n_32413) );
na02f80 g764373 ( .a(n_16219), .b(n_16368), .o(n_16390) );
in01f80 g755715 ( .a(n_24465), .o(n_24466) );
oa12f80 g771180 ( .a(n_9560), .b(n_9794), .c(n_9656), .o(n_9822) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_8_ ( .ck(newNet_2042), .d(n_5408), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_) );
no02f80 g747420 ( .a(n_32388), .b(n_44962), .o(n_32435) );
no02f80 g748333 ( .a(FE_OCP_RBN3083_n_31819), .b(n_30594), .o(n_31860) );
in01f80 newInst_3270 ( .a(newNet_3269), .o(newNet_3270) );
no02f80 g772657 ( .a(n_8163), .b(n_7743), .o(n_8184) );
oa22f80 g770345 ( .a(n_10712), .b(FE_OCP_RBN3607_n_8981), .c(n_10630), .d(FE_OFN349_n_8981), .o(n_10746) );
na02f80 g751593 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_24_), .o(n_28647) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_23_ ( .ck(newNet_2381), .d(n_36449), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_) );
in01f80 g738075 ( .a(n_42128), .o(n_42129) );
no02f80 FE_RC_1192_0 ( .a(n_13599), .b(FE_RN_362_0), .o(n_13724) );
in01f80 g777778 ( .a(n_3396), .o(n_3440) );
no02f80 g773682 ( .a(n_7933), .b(n_7795), .o(n_7388) );
in01f80 newInst_3693 ( .a(newNet_3692), .o(newNet_3693) );
no02f80 g761062 ( .a(n_19210), .b(n_18820), .o(n_19274) );
no02f80 g740396 ( .a(FE_OCP_RBN3021_n_39942), .b(n_39910), .o(n_40206) );
na02f80 FE_RC_3730_0 ( .a(FE_RN_1640_0), .b(FE_RN_1641_0), .o(FE_RN_1642_0) );
in01f80 newInst_556 ( .a(newNet_555), .o(newNet_556) );
in01f80 g752537 ( .a(n_27648), .o(n_27649) );
in01f80 g743029 ( .a(n_37155), .o(n_37156) );
na02f80 g772523 ( .a(n_8454), .b(n_8453), .o(n_8535) );
in01f80 FE_OCP_RBC3392_n_37557 ( .a(n_37557), .o(FE_OCP_RBN3392_n_37557) );
oa12f80 g759448 ( .a(n_21886), .b(n_21885), .c(n_21884), .o(n_21931) );
na02f80 g772358 ( .a(n_8603), .b(n_8515), .o(n_8604) );
in01f80 g745945 ( .a(n_33985), .o(n_33986) );
in01f80 newInst_2578 ( .a(newNet_2577), .o(newNet_2578) );
na02f80 g764308 ( .a(n_16328), .b(n_14805), .o(n_16374) );
no02f80 g774364 ( .a(n_6741), .b(n_6625), .o(n_7242) );
no02f80 g774290 ( .a(n_6816), .b(n_6815), .o(n_6817) );
ao22s80 FE_RC_1329_0 ( .a(n_34335), .b(n_34829), .c(n_34334), .d(n_34793), .o(n_34934) );
in01f80 g746714 ( .a(n_33204), .o(n_33162) );
na02f80 g749707 ( .a(n_30056), .b(n_30023), .o(n_30024) );
na02f80 g743962 ( .a(n_35699), .b(n_35749), .o(n_35750) );
ao12f80 g776141 ( .a(n_4799), .b(n_4951), .c(n_4673), .o(n_4990) );
in01f80 newInst_2317 ( .a(newNet_2316), .o(newNet_2317) );
in01f80 newInst_992 ( .a(newNet_991), .o(newNet_992) );
ao22s80 g779878 ( .a(n_1282), .b(n_902), .c(n_44650), .d(n_934), .o(n_1356) );
oa12f80 g773222 ( .a(n_7233), .b(n_7542), .c(n_7204), .o(n_7636) );
in01f80 g768237 ( .a(n_12753), .o(n_12709) );
in01f80 g737756 ( .a(n_42679), .o(n_42680) );
na02f80 g754929 ( .a(n_25481), .b(n_24774), .o(n_25694) );
no02f80 g763022 ( .a(n_17484), .b(n_17023), .o(n_17559) );
in01f80 g778278 ( .a(n_2669), .o(n_2670) );
na02f80 g738016 ( .a(n_42150), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42165) );
in01f80 newInst_202 ( .a(newNet_201), .o(newNet_202) );
no02f80 g748006 ( .a(n_33004), .b(n_32506), .o(n_33029) );
na02f80 g749520 ( .a(n_31815), .b(n_31287), .o(n_31857) );
no03m80 g747088 ( .a(n_33997), .b(n_34020), .c(n_33671), .o(n_34104) );
na02f80 g762100 ( .a(n_18177), .b(n_18176), .o(n_18178) );
in01f80 newInst_30 ( .a(newNet_29), .o(newNet_30) );
in01f80 g779045 ( .a(n_2346), .o(n_2870) );
no02f80 g756868 ( .a(n_23905), .b(n_23907), .o(n_24006) );
na02f80 g763939 ( .a(n_16624), .b(n_16599), .o(n_16642) );
in01f80 newInst_1040 ( .a(newNet_1039), .o(newNet_1040) );
in01f80 g750141 ( .a(n_29862), .o(n_29863) );
na02f80 g745577 ( .a(n_34291), .b(n_34293), .o(n_34320) );
na02f80 g759754 ( .a(n_21516), .b(n_21404), .o(n_21480) );
na02f80 g759552 ( .a(n_20767), .b(n_20464), .o(n_20817) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_24_ ( .ck(newNet_3041), .d(n_1190), .o(delay_add_ln22_unr2_stage2_stallmux_q_24_) );
in01f80 newInst_3528 ( .a(newNet_1543), .o(newNet_3528) );
oa12f80 g754751 ( .a(n_26135), .b(n_26161), .c(n_26134), .o(n_26734) );
in01f80 fopt783333 ( .a(n_44920), .o(n_44877) );
in01f80 fopt782723 ( .a(n_44102), .o(n_44104) );
in01f80 FE_OCP_RBC2947_n_10722 ( .a(n_10722), .o(FE_OCP_RBN2947_n_10722) );
na02f80 g736668 ( .a(n_43473), .b(n_43006), .o(n_43474) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_9_ ( .ck(newNet_2333), .d(n_35922), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_) );
no02f80 g779209 ( .a(n_1837), .b(delay_add_ln22_unr2_stage2_stallmux_q_9_), .o(n_1856) );
na02f80 FE_RC_4164_0 ( .a(n_12574), .b(n_13059), .o(FE_RN_1814_0) );
no02f80 g771957 ( .a(FE_OCP_RBN3571_n_44563), .b(n_9223), .o(n_9308) );
na02f80 g740414 ( .a(FE_OCP_RBN3022_n_39942), .b(n_40028), .o(n_40100) );
in01f80 g736594 ( .a(n_43446), .o(n_43447) );
no02f80 g772010 ( .a(FE_OCPN903_n_44581), .b(n_9321), .o(n_9385) );
in01f80 drc784145 ( .a(n_45891), .o(n_45894) );
in01f80 g742851 ( .a(n_37251), .o(n_37286) );
no02f80 g741725 ( .a(n_46417), .b(n_38213), .o(n_38535) );
na02f80 g765334 ( .a(FE_OCP_RBN2708_n_15135), .b(FE_OCP_RBN2455_n_14157), .o(n_15452) );
na02f80 g768502 ( .a(n_12342), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_9_), .o(n_12385) );
in01f80 newInst_1893 ( .a(newNet_1892), .o(newNet_1893) );
in01f80 newInst_1489 ( .a(newNet_1488), .o(newNet_1489) );
oa22f80 g762676 ( .a(n_18183), .b(n_17703), .c(n_18184), .d(n_17702), .o(n_18251) );
na02f80 g752920 ( .a(n_27722), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_), .o(n_27812) );
in01f80 g768399 ( .a(n_12500), .o(n_12501) );
no02f80 g756821 ( .a(n_24076), .b(n_24059), .o(n_24355) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_12_ ( .ck(newNet_2122), .d(n_5841), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_12_) );
in01f80 FE_OCP_RBC2650_n_9042 ( .a(n_9042), .o(FE_OCP_RBN2650_n_9042) );
na02f80 g747871 ( .a(n_33128), .b(n_33127), .o(n_33129) );
in01f80 newInst_273 ( .a(newNet_78), .o(newNet_273) );
na02f80 g774476 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(n_6564) );
in01f80 g776061 ( .a(n_4683), .o(n_4684) );
na02f80 g743677 ( .a(n_36328), .b(n_35683), .o(n_36394) );
no02f80 FE_RC_2073_0 ( .a(n_30577), .b(n_30173), .o(FE_RN_707_0) );
no02f80 g763823 ( .a(n_17362), .b(n_17422), .o(n_17958) );
in01f80 g772258 ( .a(n_8831), .o(n_8832) );
ao12f80 g765372 ( .a(n_16135), .b(n_15874), .c(n_15564), .o(n_16352) );
in01f80 g742496 ( .a(n_37609), .o(n_37582) );
no02f80 g740653 ( .a(n_39584), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39603) );
na02f80 g768130 ( .a(n_12662), .b(n_12085), .o(n_12703) );
in01f80 newInst_3587 ( .a(newNet_3586), .o(newNet_3587) );
na02f80 g764832 ( .a(n_15792), .b(FE_OFN823_n_15791), .o(n_15934) );
in01f80 g768115 ( .a(n_12633), .o(n_12634) );
na02f80 g762252 ( .a(n_18579), .b(n_18622), .o(n_18661) );
na02f80 g769786 ( .a(n_11139), .b(n_11063), .o(n_11174) );
in01f80 g771162 ( .a(n_9621), .o(n_9715) );
in01f80 FE_OCPC843_n_3912 ( .a(n_3912), .o(FE_OCPN843_n_3912) );
in01f80 newInst_741 ( .a(newNet_402), .o(newNet_741) );
no02f80 g753120 ( .a(n_27213), .b(n_27172), .o(n_27264) );
in01f80 newInst_1848 ( .a(newNet_1281), .o(newNet_1848) );
na02f80 g768282 ( .a(n_12641), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .o(n_12697) );
na02f80 g754850 ( .a(n_25486), .b(n_25424), .o(n_25509) );
no02f80 g761042 ( .a(n_19211), .b(FE_OFN779_n_17093), .o(n_19565) );
no02f80 g776683 ( .a(n_3787), .b(n_3838), .o(n_5603) );
no02f80 g737489 ( .a(n_42636), .b(n_42644), .o(n_42665) );
in01f80 newInst_703 ( .a(newNet_702), .o(newNet_703) );
in01f80 g753407 ( .a(n_27611), .o(n_27612) );
in01f80 g741768 ( .a(n_38553), .o(n_38514) );
oa22f80 g751935 ( .a(n_28919), .b(n_28134), .c(n_28897), .d(n_28993), .o(n_29245) );
in01f80 g756932 ( .a(n_23906), .o(n_23907) );
na02f80 g752510 ( .a(n_27659), .b(n_27465), .o(n_27685) );
in01f80 g749553 ( .a(n_30428), .o(n_30427) );
in01f80 newInst_1789 ( .a(newNet_1788), .o(newNet_1789) );
na02f80 g759101 ( .a(n_21092), .b(n_21016), .o(n_21132) );
no02f80 g773662 ( .a(n_7323), .b(n_7322), .o(n_7324) );
in01f80 newInst_144 ( .a(newNet_143), .o(newNet_144) );
na02f80 g760067 ( .a(n_20606), .b(n_20573), .o(n_20670) );
na02f80 FE_RC_3586_0 ( .a(FE_RN_1563_0), .b(n_44174), .o(n_35615) );
in01f80 newInst_3156 ( .a(newNet_2799), .o(newNet_3156) );
no02f80 g767996 ( .a(n_12630), .b(n_12653), .o(n_13889) );
in01f80 FE_OCPC3758_n_2346 ( .a(n_2346), .o(FE_OCPN3758_n_2346) );
in01f80 g759580 ( .a(n_20821), .o(n_20850) );
ao12f80 g755275 ( .a(n_25521), .b(n_25638), .c(n_25548), .o(n_25607) );
oa12f80 g748732 ( .a(n_31035), .b(n_31086), .c(n_31138), .o(n_31141) );
na02f80 g778525 ( .a(n_2369), .b(n_2351), .o(n_2352) );
in01f80 g777720 ( .a(n_3313), .o(n_3331) );
in01f80 FE_RC_2987_0 ( .a(n_11144), .o(FE_RN_1304_0) );
oa22f80 g752593 ( .a(n_27591), .b(n_27270), .c(n_27590), .d(n_27271), .o(n_27665) );
in01f80 fopt783450 ( .a(n_45012), .o(n_45010) );
in01f80 g737675 ( .a(n_42754), .o(n_42755) );
ao12f80 g765865 ( .a(n_15246), .b(n_15245), .c(n_15244), .o(n_15711) );
in01f80 g752170 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .o(n_27922) );
in01f80 FE_OCP_RBC2873_n_10477 ( .a(n_10477), .o(FE_OCP_RBN2873_n_10477) );
in01f80 newInst_987 ( .a(newNet_19), .o(newNet_987) );
no02f80 g749761 ( .a(n_31224), .b(n_31223), .o(n_31225) );
na02f80 FE_RC_4146_0 ( .a(FE_RN_1801_0), .b(n_44721), .o(FE_RN_1802_0) );
in01f80 FE_RC_1340_0 ( .a(n_4416), .o(FE_RN_399_0) );
in01f80 FE_OCP_RBC3418_n_12739 ( .a(FE_OCP_RBN3416_n_12739), .o(FE_OCP_RBN3418_n_12739) );
in01f80 FE_RC_3094_0 ( .a(FE_RN_1367_0), .o(n_26190) );
in01f80 newInst_2372 ( .a(newNet_2371), .o(newNet_2372) );
in01f80 newInst_200 ( .a(newNet_199), .o(newNet_200) );
in01f80 g773666 ( .a(n_7300), .o(n_7301) );
na02f80 g780212 ( .a(n_1042), .b(n_1111), .o(n_1128) );
in01f80 g762966 ( .a(n_17765), .o(n_17744) );
no02f80 g772785 ( .a(FE_OCP_RBN2383_n_8342), .b(FE_OCPN940_n_7712), .o(n_8176) );
in01f80 newInst_2411 ( .a(newNet_2410), .o(newNet_2411) );
oa12f80 g764555 ( .a(n_16510), .b(n_16509), .c(n_16508), .o(n_16549) );
in01f80 g778307 ( .a(n_2849), .o(n_2894) );
no02f80 g757266 ( .a(n_23495), .b(n_22926), .o(n_23527) );
oa12f80 g769994 ( .a(n_10811), .b(n_10874), .c(n_10748), .o(n_10948) );
in01f80 g768431 ( .a(n_12413), .o(n_12449) );
in01f80 FE_RC_2387_0 ( .a(n_42443), .o(FE_RN_934_0) );
na03f80 FE_RC_1290_0 ( .a(n_3184), .b(n_3216), .c(n_3187), .o(n_3272) );
no02f80 g780804 ( .a(n_468), .b(n_467), .o(n_469) );
in01f80 g765974 ( .a(n_14789), .o(n_14811) );
in01f80 newInst_492 ( .a(newNet_491), .o(newNet_492) );
na02f80 FE_RC_2208_0 ( .a(FE_RN_794_0), .b(n_27554), .o(n_27568) );
na02f80 g740225 ( .a(n_40056), .b(FE_OCP_RBN3027_n_39942), .o(n_40134) );
no02f80 g763896 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_16_), .o(n_17464) );
no02f80 g749444 ( .a(FE_OCP_RBN2755_n_30558), .b(n_30577), .o(n_30579) );
no02f80 g771923 ( .a(n_8876), .b(n_8916), .o(n_8995) );
no02f80 g759789 ( .a(n_21694), .b(FE_OCP_RBN3678_n_21051), .o(n_21778) );
no02f80 g736339 ( .a(n_43833), .b(n_43646), .o(n_43846) );
no02f80 g769327 ( .a(FE_OCPN858_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .o(n_11974) );
na02f80 g762449 ( .a(n_18351), .b(n_18350), .o(n_18352) );
in01f80 g774351 ( .a(n_6651), .o(n_6539) );
in01f80 g757823 ( .a(n_22511), .o(n_22531) );
in01f80 g743188 ( .a(n_36878), .o(n_36879) );
no02f80 g762655 ( .a(n_18256), .b(n_18255), .o(n_18257) );
na02f80 g752168 ( .a(n_28008), .b(n_27975), .o(n_28086) );
na02f80 g776801 ( .a(n_4263), .b(n_4155), .o(n_4236) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_13_ ( .ck(newNet_749), .d(n_46166), .o(delay_xor_ln21_unr6_stage3_stallmux_q_13_) );
na02f80 g777695 ( .a(n_3407), .b(n_2759), .o(n_3408) );
na02f80 g742439 ( .a(n_37658), .b(n_36948), .o(n_37738) );
oa22f80 g748193 ( .a(n_31497), .b(n_31471), .c(n_31498), .d(n_31472), .o(n_31561) );
in01f80 g780742 ( .a(n_596), .o(n_601) );
na02f80 g748648 ( .a(n_32610), .b(n_32589), .o(n_32590) );
in01f80 g769348 ( .a(n_11711), .o(n_11797) );
oa12f80 g756954 ( .a(n_23620), .b(n_23619), .c(n_23618), .o(n_23701) );
na02f80 g768106 ( .a(FE_OCP_RBN2219_n_12698), .b(n_12734), .o(n_12736) );
no02f80 g756870 ( .a(n_23990), .b(n_23951), .o(n_24706) );
na02f80 g762640 ( .a(n_17932), .b(n_17931), .o(n_17999) );
oa12f80 g770660 ( .a(n_10289), .b(n_10353), .c(n_10288), .o(n_10392) );
in01f80 newInst_590 ( .a(newNet_589), .o(newNet_590) );
in01f80 g748199 ( .a(n_32180), .o(n_32181) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_11_ ( .ck(newNet_758), .d(n_46159), .o(delay_xor_ln21_unr6_stage3_stallmux_q_11_) );
na02f80 g770700 ( .a(n_9941), .b(FE_OCP_RBN2474_n_8664), .o(n_10022) );
na02f80 g760547 ( .a(n_19894), .b(n_19893), .o(n_20106) );
no02f80 g758327 ( .a(n_22187), .b(FE_OCP_RBN1378_n_20889), .o(n_22212) );
in01f80 newInst_396 ( .a(newNet_395), .o(newNet_396) );
in01f80 newInst_1742 ( .a(newNet_1741), .o(newNet_1742) );
in01f80 g750606 ( .a(n_29422), .o(n_29475) );
na02f80 g777729 ( .a(n_3338), .b(n_2759), .o(n_3339) );
no02f80 g779546 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_26_), .o(n_2108) );
in01f80 newInst_2786 ( .a(newNet_2785), .o(newNet_2786) );
in01f80 FE_OCP_RBC1839_n_19528 ( .a(n_19528), .o(FE_OCP_RBN1839_n_19528) );
na02f80 g765652 ( .a(n_14988), .b(FE_OCP_RBN2503_n_13896), .o(n_14989) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_7_ ( .ck(newNet_1924), .d(n_36895), .o(delay_sub_ln21_unr24_stage9_stallmux_q_7_) );
na02f80 g754417 ( .a(n_25704), .b(n_25412), .o(n_25705) );
no02f80 g743620 ( .a(n_36483), .b(n_36010), .o(n_36485) );
no02f80 g760961 ( .a(FE_OCP_RBN1345_n_19270), .b(n_19218), .o(n_19331) );
oa22f80 g752663 ( .a(n_27314), .b(n_27225), .c(n_27313), .d(n_27224), .o(n_27443) );
no02f80 g755325 ( .a(n_24883), .b(n_24897), .o(n_24884) );
na02f80 g770677 ( .a(n_10072), .b(n_44464), .o(n_10104) );
na02f80 g738710 ( .a(n_41716), .b(n_41482), .o(n_41875) );
in01f80 g741159 ( .a(n_38966), .o(n_38924) );
no02f80 g767530 ( .a(n_13382), .b(n_12995), .o(n_13393) );
in01f80 newInst_541 ( .a(newNet_540), .o(newNet_541) );
in01f80 g778208 ( .a(n_2747), .o(n_2801) );
no02f80 g773761 ( .a(n_7241), .b(n_7046), .o(n_7279) );
no02f80 g771845 ( .a(n_44516), .b(n_10079), .o(n_10123) );
no02f80 g746393 ( .a(n_33410), .b(FE_OCP_RBN2178_n_33022), .o(n_33489) );
na03f80 g742649 ( .a(n_37215), .b(n_37376), .c(n_36974), .o(n_37459) );
na02f80 g773635 ( .a(n_7389), .b(n_7386), .o(n_7387) );
ao22s80 FE_RC_232_0 ( .a(FE_OCP_RBN2249_n_13017), .b(n_14069), .c(n_14070), .d(FE_OCP_RBN2250_n_13017), .o(n_14249) );
no02f80 g764884 ( .a(n_15790), .b(n_15724), .o(n_15886) );
no02f80 g764864 ( .a(n_15623), .b(n_15622), .o(n_15649) );
in01f80 g746114 ( .a(n_35765), .o(n_35217) );
na02f80 g759747 ( .a(n_20502), .b(n_45010), .o(n_20587) );
ao22s80 FE_RC_226_0 ( .a(FE_OCP_RBN3399_n_12751), .b(n_12578), .c(n_12751), .d(n_12577), .o(n_12902) );
oa12f80 g736374 ( .a(n_312), .b(n_43785), .c(FE_OFN3_n_43918), .o(n_43824) );
in01f80 g742981 ( .a(n_37079), .o(n_36971) );
in01f80 newInst_2335 ( .a(newNet_908), .o(newNet_2335) );
in01f80 g774766 ( .a(n_6471), .o(n_6472) );
na02f80 g743521 ( .a(FE_OCP_RBN1326_n_36489), .b(n_36750), .o(n_36519) );
oa12f80 g762902 ( .a(n_17993), .b(n_17994), .c(n_17992), .o(n_18420) );
oa22f80 g740781 ( .a(n_39430), .b(n_39185), .c(n_39493), .d(n_39186), .o(n_39531) );
no02f80 g768346 ( .a(n_12584), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .o(n_12947) );
in01f80 g774730 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_21_), .o(n_7401) );
na02f80 g753141 ( .a(n_27303), .b(n_27339), .o(n_27459) );
na02f80 g748930 ( .a(n_31154), .b(n_31070), .o(n_31199) );
in01f80 newInst_2990 ( .a(newNet_2989), .o(newNet_2990) );
oa12f80 g776674 ( .a(n_3651), .b(n_3822), .c(n_3749), .o(n_3992) );
oa22f80 g737957 ( .a(n_42169), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .c(n_42170), .d(n_42196), .o(n_42187) );
ao12f80 g741086 ( .a(n_39034), .b(n_39033), .c(n_39032), .o(n_39800) );
no02f80 g776902 ( .a(n_3681), .b(n_2946), .o(n_3723) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_23_ ( .ck(newNet_2469), .d(n_32471), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_) );
na02f80 g764270 ( .a(n_16389), .b(n_16424), .o(n_16511) );
in01f80 FE_OCPC1749_n_27223 ( .a(n_27223), .o(FE_OCPN1749_n_27223) );
in01f80 g752715 ( .a(n_27241), .o(n_27242) );
no02f80 g743309 ( .a(n_36674), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36710) );
no02f80 g748407 ( .a(n_31730), .b(n_30729), .o(n_31731) );
no02f80 g763526 ( .a(FE_OCP_RBN3082_n_16977), .b(n_16117), .o(n_16978) );
no02f80 FE_RC_1792_0 ( .a(n_34162), .b(n_34522), .o(FE_RN_528_0) );
oa22f80 FE_RC_1717_0 ( .a(n_17336), .b(n_17440), .c(n_17753), .d(n_17334), .o(n_17476) );
na02f80 g745517 ( .a(n_34381), .b(n_34380), .o(n_34382) );
in01f80 FE_RC_410_0 ( .a(n_13257), .o(FE_RN_120_0) );
na02f80 g777699 ( .a(n_3403), .b(n_3006), .o(n_3458) );
na02f80 g768261 ( .a(n_12673), .b(n_12672), .o(n_12733) );
na02f80 g749966 ( .a(n_29984), .b(n_29890), .o(n_30012) );
no02f80 g748754 ( .a(n_31058), .b(n_30965), .o(n_31087) );
in01f80 newInst_2892 ( .a(newNet_1633), .o(newNet_2892) );
in01f80 g738803 ( .a(n_41478), .o(n_41525) );
no02f80 g760308 ( .a(n_20214), .b(n_20125), .o(n_20227) );
na02f80 g772501 ( .a(n_8344), .b(n_8403), .o(n_8404) );
in01f80 g766736 ( .a(n_13806), .o(n_13807) );
oa12f80 g772766 ( .a(n_8142), .b(n_8141), .c(n_8140), .o(n_9790) );
na02f80 g763294 ( .a(n_17329), .b(n_17328), .o(n_17330) );
na02f80 g760090 ( .a(n_20340), .b(FE_OCP_RBN1694_n_19052), .o(n_20341) );
ao12f80 g758157 ( .a(n_22690), .b(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_9_), .o(n_22726) );
in01f80 FE_OCP_RBC2516_n_8657 ( .a(n_8657), .o(FE_OCP_RBN2516_n_8657) );
no02f80 g780020 ( .a(n_1258), .b(n_1020), .o(n_1266) );
no03m80 g756176 ( .a(n_24132), .b(n_24792), .c(n_24151), .o(n_24904) );
in01f80 g758332 ( .a(n_22291), .o(n_22417) );
in01f80 FE_OCP_RBC2133_n_45508 ( .a(n_45508), .o(FE_OCP_RBN2133_n_45508) );
na02f80 g775077 ( .a(n_6052), .b(n_5174), .o(n_6111) );
in01f80 g759222 ( .a(n_21012), .o(n_21013) );
na02f80 FE_RC_3636_0 ( .a(FE_RN_1594_0), .b(n_30324), .o(FE_RN_1595_0) );
na02f80 g762749 ( .a(n_17913), .b(n_17966), .o(n_18041) );
in01f80 FE_OCP_RBC3687_n_5105 ( .a(n_5105), .o(FE_OCP_RBN3687_n_5105) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_18_ ( .ck(newNet_647), .d(n_46353), .o(delay_xor_ln21_unr9_stage4_stallmux_q_18_) );
in01f80 g776472 ( .a(n_4398), .o(n_4399) );
no02f80 g766030 ( .a(n_14716), .b(n_13563), .o(n_14717) );
no02f80 g744151 ( .a(n_36095), .b(n_36000), .o(n_36139) );
in01f80 g778031 ( .a(n_3102), .o(n_3103) );
no02f80 g749346 ( .a(n_30674), .b(n_30701), .o(n_30824) );
in01f80 g749331 ( .a(n_30747), .o(n_30651) );
na02f80 g759999 ( .a(n_20752), .b(n_20664), .o(n_20753) );
oa22f80 FE_RC_3794_0 ( .a(n_38722), .b(n_38751), .c(n_38720), .d(n_38750), .o(n_38800) );
no02f80 g749687 ( .a(n_31192), .b(n_31294), .o(n_31258) );
no02f80 FE_RC_2888_0 ( .a(FE_RN_1249_0), .b(n_14535), .o(FE_RN_1250_0) );
no02f80 g763431 ( .a(n_17454), .b(n_17022), .o(n_17268) );
in01f80 g758507 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_11_), .o(n_23376) );
in01f80 g764125 ( .a(n_46979), .o(n_16634) );
in01f80 newInst_1008 ( .a(newNet_1007), .o(newNet_1008) );
in01f80 FE_OCP_RBC2367_n_24408 ( .a(n_24408), .o(FE_OCP_RBN2367_n_24408) );
oa12f80 g747233 ( .a(n_32694), .b(n_32693), .c(n_32692), .o(n_33917) );
ao12f80 g764924 ( .a(n_15644), .b(n_15676), .c(n_15531), .o(n_15680) );
in01f80 g738236 ( .a(n_41955), .o(n_42276) );
oa12f80 g755908 ( .a(n_25307), .b(n_25160), .c(n_25251), .o(n_25710) );
in01f80 FE_OCP_RBC3356_delay_xor_ln22_unr28_stage10_stallmux_q_0_ ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(FE_OCP_RBN3356_delay_xor_ln22_unr28_stage10_stallmux_q_0_) );
no02f80 g776513 ( .a(n_4385), .b(n_4308), .o(n_4386) );
in01f80 g738672 ( .a(n_41688), .o(n_41657) );
in01f80 FE_OCP_RBC2171_n_32892 ( .a(FE_OCP_RBN2170_n_32892), .o(FE_OCP_RBN2171_n_32892) );
in01f80 newInst_1163 ( .a(newNet_24), .o(newNet_1163) );
no02f80 g757926 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n_23055) );
in01f80 newInst_2298 ( .a(newNet_2297), .o(newNet_2298) );
oa22f80 g745079 ( .a(n_36180), .b(n_35767), .c(n_36179), .d(n_35768), .o(n_36286) );
na02f80 g747626 ( .a(n_33464), .b(n_33419), .o(n_33997) );
na02f80 FE_RC_521_0 ( .a(FE_RN_162_0), .b(FE_RN_163_0), .o(FE_RN_164_0) );
in01f80 g754391 ( .a(n_25843), .o(n_25869) );
in01f80 FE_RC_2959_0 ( .a(n_39822), .o(FE_RN_1292_0) );
no02f80 g778062 ( .a(n_2994), .b(FE_OCP_RBN3486_n_2438), .o(n_2995) );
oa22f80 g784349 ( .a(FE_OCP_RBN3078_FE_OFN807_n_46195), .b(n_6267), .c(FE_OFN774_n_46137), .d(n_6245), .o(n_46155) );
in01f80 g738328 ( .a(n_42209), .o(n_42267) );
no02f80 g757086 ( .a(n_23235), .b(n_23234), .o(n_23236) );
oa22f80 g749822 ( .a(n_31311), .b(n_31256), .c(n_31530), .d(n_31211), .o(n_31564) );
in01f80 newInst_1011 ( .a(newNet_248), .o(newNet_1011) );
in01f80 g739351 ( .a(n_40674), .o(n_40689) );
oa12f80 g741745 ( .a(n_38492), .b(n_38491), .c(n_38490), .o(n_38564) );
in01f80 g777579 ( .a(n_3700), .o(n_3788) );
oa22f80 g747775 ( .a(n_33372), .b(n_33316), .c(n_33571), .d(n_33310), .o(n_33912) );
in01f80 g766464 ( .a(n_14225), .o(n_14265) );
no02f80 g737420 ( .a(n_42736), .b(n_42361), .o(n_42737) );
ao22s80 FE_RC_823_0 ( .a(FE_OCP_RBN2339_n_29385), .b(n_28803), .c(n_28802), .d(n_29385), .o(n_29480) );
in01f80 FE_OCPC1483_n_18953 ( .a(n_18953), .o(FE_OCPN1483_n_18953) );
in01f80 g748139 ( .a(n_31948), .o(n_31949) );
no02f80 g748914 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_), .o(n_32408) );
na02f80 g771005 ( .a(n_9960), .b(n_10034), .o(n_10139) );
in01f80 g739063 ( .a(n_41119), .o(n_41085) );
in01f80 g767697 ( .a(n_13156), .o(n_13157) );
no02f80 g760549 ( .a(n_19916), .b(n_18288), .o(n_20077) );
in01f80 g749220 ( .a(n_30849), .o(n_30871) );
na02f80 g756861 ( .a(n_23334), .b(n_23249), .o(n_23348) );
no02f80 g784768 ( .a(n_44102), .b(FE_OCP_RBN2269_n_33803), .o(n_47254) );
oa12f80 g744660 ( .a(n_35889), .b(n_36555), .c(n_35934), .o(n_36599) );
ao12f80 g762464 ( .a(n_17710), .b(n_45524), .c(n_17611), .o(n_18386) );
in01f80 FE_RC_4157_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(FE_RN_1809_0) );
no02f80 g778504 ( .a(n_2336), .b(n_2373), .o(n_2520) );
in01f80 g765500 ( .a(n_15928), .o(n_15822) );
in01f80 g766443 ( .a(n_14191), .o(n_14152) );
in01f80 g744790 ( .a(n_35146), .o(n_35147) );
in01f80 g774201 ( .a(n_7161), .o(n_7162) );
in01f80 FE_RC_1544_0 ( .a(n_28226), .o(FE_RN_435_0) );
in01f80 newInst_1083 ( .a(newNet_1082), .o(newNet_1083) );
na02f80 g775619 ( .a(n_5458), .b(n_4606), .o(n_5472) );
oa22f80 FE_RC_1267_0 ( .a(n_38234), .b(n_38546), .c(n_38233), .d(n_38547), .o(n_38592) );
in01f80 g773701 ( .a(n_7309), .o(n_7310) );
in01f80 newInst_782 ( .a(newNet_93), .o(newNet_782) );
in01f80 g753474 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_5_), .o(n_28220) );
in01f80 fopt783930 ( .a(n_27639), .o(n_45638) );
na02f80 g746694 ( .a(n_33290), .b(n_33217), .o(n_33340) );
in01f80 g741003 ( .a(n_39163), .o(n_39158) );
in01f80 newInst_311 ( .a(newNet_310), .o(newNet_311) );
no02f80 g773611 ( .a(n_7377), .b(n_6863), .o(n_7413) );
no02f80 g744980 ( .a(n_34994), .b(n_34625), .o(n_34992) );
no02f80 g747303 ( .a(n_32706), .b(n_32527), .o(n_32597) );
no02f80 g769746 ( .a(n_11124), .b(n_11125), .o(n_11209) );
in01f80 g744321 ( .a(n_35545), .o(n_35546) );
no02f80 g768786 ( .a(n_12097), .b(n_12069), .o(n_12177) );
in01f80 g763867 ( .a(n_16757), .o(n_16725) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_14_ ( .ck(newNet_512), .d(n_22949), .o(delay_xor_ln22_unr15_stage6_stallmux_q_14_) );
no02f80 FE_RC_4028_0 ( .a(FE_RN_1749_0), .b(n_15900), .o(FE_RN_1750_0) );
no02f80 g776250 ( .a(n_4847), .b(n_4368), .o(n_4913) );
in01f80 newInst_172 ( .a(newNet_171), .o(newNet_172) );
oa12f80 g784646 ( .a(n_16703), .b(n_16640), .c(n_16656), .o(n_46976) );
na02f80 g765402 ( .a(n_15177), .b(n_15170), .o(n_15296) );
in01f80 newInst_2768 ( .a(newNet_2767), .o(newNet_2768) );
in01f80 g778554 ( .a(n_2392), .o(n_2361) );
na02f80 g753773 ( .a(FE_OCP_RBN2968_n_26398), .b(FE_OCP_RBN2939_n_26276), .o(n_26471) );
no02f80 g778703 ( .a(n_2235), .b(n_2234), .o(n_2258) );
na02f80 g763166 ( .a(n_17402), .b(n_17285), .o(n_17483) );
in01f80 g782659 ( .a(n_44053), .o(n_44054) );
in01f80 g755302 ( .a(n_24898), .o(n_24899) );
na02f80 g750132 ( .a(n_29840), .b(n_28776), .o(n_29984) );
na02f80 g748979 ( .a(n_31073), .b(FE_OCPN1452_n_27518), .o(n_31105) );
oa12f80 g766687 ( .a(n_14562), .b(n_14529), .c(n_14527), .o(n_14619) );
in01f80 g761686 ( .a(n_18650), .o(n_18759) );
in01f80 FE_OCP_RBC2866_n_39640 ( .a(n_39640), .o(FE_OCP_RBN2866_n_39640) );
no02f80 g755182 ( .a(n_25115), .b(n_23893), .o(n_25175) );
no02f80 g760622 ( .a(n_19776), .b(n_19837), .o(n_19896) );
no02f80 g758949 ( .a(n_21640), .b(FE_OCP_DRV_N1602_n_21639), .o(n_21676) );
no02f80 g776163 ( .a(n_4933), .b(n_4348), .o(n_5012) );
in01f80 g742197 ( .a(n_38227), .o(n_38228) );
na02f80 g738690 ( .a(n_41716), .b(n_41494), .o(n_41826) );
in01f80 g761667 ( .a(n_18754), .o(n_18755) );
no02f80 g758747 ( .a(n_21621), .b(n_21508), .o(n_21665) );
ao22s80 g771917 ( .a(n_44575), .b(n_8514), .c(n_44566), .d(n_10214), .o(n_9035) );
no02f80 g753191 ( .a(n_27103), .b(n_25909), .o(n_27121) );
in01f80 g771742 ( .a(n_8850), .o(n_8851) );
no02f80 g760816 ( .a(n_19474), .b(n_19202), .o(n_19475) );
no02f80 FE_RC_1415_0 ( .a(FE_RN_413_0), .b(n_15728), .o(n_46981) );
na02f80 g777065 ( .a(n_3833), .b(n_3604), .o(n_4034) );
in01f80 newInst_726 ( .a(newNet_725), .o(newNet_726) );
oa12f80 g765954 ( .a(n_14573), .b(n_14673), .c(n_14572), .o(n_14771) );
na02f80 g751795 ( .a(n_28286), .b(n_28285), .o(n_28425) );
in01f80 FE_OCPC964_n_27287 ( .a(FE_OCPN963_n_27287), .o(FE_OCPN964_n_27287) );
in01f80 g768884 ( .a(n_11929), .o(n_11876) );
na02f80 g768684 ( .a(n_12098), .b(n_10371), .o(n_12253) );
no02f80 g752185 ( .a(n_27944), .b(n_44735), .o(n_28064) );
na02f80 g752137 ( .a(n_28116), .b(n_28115), .o(n_28181) );
in01f80 g779356 ( .a(n_1638), .o(n_1639) );
na02f80 g772586 ( .a(n_8332), .b(n_8355), .o(n_8439) );
in01f80 g767090 ( .a(n_13532), .o(n_13533) );
oa22f80 FE_RC_3248_0 ( .a(n_20671), .b(n_21088), .c(n_20670), .d(FE_OCP_RBN1218_n_21088), .o(n_21238) );
in01f80 FE_RC_1334_0 ( .a(n_4647), .o(FE_RN_396_0) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_28_ ( .ck(newNet_2634), .d(FE_OCP_RBN3118_n_22755), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_) );
no02f80 g772872 ( .a(n_7958), .b(n_7942), .o(n_8100) );
in01f80 g759700 ( .a(n_21865), .o(n_21866) );
na02f80 g760586 ( .a(n_19812), .b(n_19785), .o(n_19842) );
no02f80 g756017 ( .a(n_25026), .b(n_24768), .o(n_25220) );
in01f80 newInst_1972 ( .a(newNet_1971), .o(newNet_1972) );
no02f80 g771533 ( .a(n_9335), .b(n_9390), .o(n_9483) );
no02f80 g776820 ( .a(n_3732), .b(n_3722), .o(n_4041) );
in01f80 newInst_2078 ( .a(newNet_933), .o(newNet_2078) );
in01f80 g756597 ( .a(n_23740), .o(n_23676) );
na02f80 g746546 ( .a(n_34886), .b(n_34938), .o(n_34962) );
no02f80 g779577 ( .a(n_1783), .b(n_1739), .o(n_2120) );
no02f80 g751797 ( .a(n_28232), .b(n_28234), .o(n_28233) );
no02f80 g737512 ( .a(n_42455), .b(n_42213), .o(n_42498) );
na02f80 g744593 ( .a(n_35276), .b(n_35297), .o(n_35368) );
na02f80 g745159 ( .a(n_35554), .b(n_34628), .o(n_34918) );
in01f80 g778653 ( .a(n_2450), .o(n_2451) );
na02f80 g754030 ( .a(n_26974), .b(n_26865), .o(n_26975) );
no02f80 g776076 ( .a(n_4927), .b(n_4371), .o(n_4945) );
no02f80 g740499 ( .a(n_39702), .b(n_39685), .o(n_39703) );
no02f80 FE_RC_2844_0 ( .a(n_47200), .b(n_11166), .o(FE_RN_1224_0) );
in01f80 FE_OCP_RBC2540_n_8781 ( .a(n_8781), .o(FE_OCP_RBN2540_n_8781) );
oa22f80 g742702 ( .a(n_37348), .b(n_37064), .c(n_37349), .d(n_37063), .o(n_37882) );
in01f80 g773887 ( .a(n_7769), .o(n_7105) );
in01f80 g776347 ( .a(n_4592), .o(n_4541) );
in01f80 g775891 ( .a(n_4916), .o(n_4968) );
na02f80 g763579 ( .a(n_16988), .b(n_16900), .o(n_17129) );
no02f80 g744839 ( .a(n_34960), .b(n_30545), .o(n_35012) );
na02f80 g738412 ( .a(n_41638), .b(n_41637), .o(n_41639) );
no02f80 g768830 ( .a(n_12005), .b(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n_11966) );
ao22s80 g736542 ( .a(n_43651), .b(n_43622), .c(n_43659), .d(n_43621), .o(n_43708) );
na02f80 g777052 ( .a(n_3582), .b(n_2848), .o(n_3632) );
oa12f80 g748611 ( .a(n_31302), .b(n_31301), .c(n_31308), .o(n_31363) );
no02f80 g761088 ( .a(n_20038), .b(n_19787), .o(n_20068) );
in01f80 FE_OCP_RBC3733_n_31819 ( .a(FE_OCP_RBN3086_n_31819), .o(FE_OCP_RBN3733_n_31819) );
no02f80 g741694 ( .a(n_38564), .b(n_38562), .o(n_38565) );
in01f80 newInst_872 ( .a(newNet_871), .o(newNet_872) );
na02f80 g757500 ( .a(n_22865), .b(FE_OCP_RBN3822_n_44061), .o(n_22866) );
ao12f80 g750957 ( .a(n_28526), .b(n_28871), .c(n_28530), .o(n_28968) );
na02f80 g769093 ( .a(n_11518), .b(n_11598), .o(n_11638) );
in01f80 FE_RC_1566_0 ( .a(n_28332), .o(FE_RN_444_0) );
na02f80 FE_RC_2221_0 ( .a(FE_RN_803_0), .b(n_33274), .o(FE_RN_804_0) );
na02f80 g770508 ( .a(n_10481), .b(n_10471), .o(n_10472) );
no02f80 g759177 ( .a(n_21266), .b(n_21214), .o(n_21348) );
no02f80 FE_RC_4051_0 ( .a(n_35746), .b(FE_RN_1761_0), .o(n_36208) );
na02f80 g766119 ( .a(n_14895), .b(n_14296), .o(n_14993) );
na02f80 g768004 ( .a(n_12809), .b(n_12732), .o(n_12819) );
na02f80 FE_RC_3044_0 ( .a(n_35360), .b(n_35377), .o(FE_RN_1333_0) );
in01f80 newInst_2306 ( .a(newNet_2305), .o(newNet_2306) );
na02f80 g753416 ( .a(n_27007), .b(FE_OCP_RBN2938_n_26456), .o(n_27039) );
na02f80 g764625 ( .a(n_16447), .b(n_16024), .o(n_16504) );
in01f80 newInst_2996 ( .a(newNet_465), .o(newNet_2996) );
in01f80 newInst_2165 ( .a(newNet_1826), .o(newNet_2165) );
ao22s80 g779115 ( .a(n_2003), .b(n_1824), .c(n_2025), .d(n_1825), .o(n_2066) );
oa22f80 g767730 ( .a(n_12799), .b(n_11943), .c(n_12798), .d(n_12747), .o(n_14676) );
in01f80 newInst_3432 ( .a(newNet_3241), .o(newNet_3432) );
in01f80 g774962 ( .a(n_6218), .o(n_6219) );
oa12f80 g760560 ( .a(n_19882), .b(n_19854), .c(n_19833), .o(n_20007) );
in01f80 g762804 ( .a(n_17782), .o(n_17756) );
na02f80 g746906 ( .a(n_33015), .b(n_31855), .o(n_33077) );
na02f80 g776917 ( .a(n_3773), .b(n_3884), .o(n_3850) );
na02f80 g756053 ( .a(n_25160), .b(n_25138), .o(n_25306) );
in01f80 g766812 ( .a(n_15482), .o(n_15513) );
no02f80 FE_RC_2881_0 ( .a(FE_OCP_RBN3651_n_39249), .b(n_39479), .o(FE_RN_1246_0) );
no02f80 g776628 ( .a(n_4221), .b(n_4240), .o(n_4315) );
na02f80 g768793 ( .a(n_11956), .b(n_11955), .o(n_11962) );
in01f80 newInst_293 ( .a(newNet_292), .o(newNet_293) );
na02f80 g746132 ( .a(n_33732), .b(n_33777), .o(n_33831) );
in01f80 g771164 ( .a(FE_OCP_RBN2748_n_9584), .o(n_9620) );
no02f80 g761347 ( .a(n_18954), .b(n_18953), .o(n_19035) );
na02f80 g764109 ( .a(n_16556), .b(n_16557), .o(n_16605) );
in01f80 FE_RC_2235_0 ( .a(n_23058), .o(FE_RN_815_0) );
na03f80 g779183 ( .a(n_1601), .b(n_1869), .c(n_1580), .o(n_1928) );
ao12f80 g768624 ( .a(n_12250), .b(n_12249), .c(n_12260), .o(n_12321) );
na02f80 g762731 ( .a(n_17721), .b(n_17778), .o(n_17804) );
in01f80 FE_RC_3183_0 ( .a(n_6716), .o(FE_RN_1412_0) );
in01f80 g778532 ( .a(n_2729), .o(n_2730) );
oa12f80 g747653 ( .a(n_33299), .b(n_33298), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_33337) );
in01f80 newInst_3366 ( .a(newNet_3365), .o(newNet_3366) );
in01f80 FE_OCPC1258_n_25353 ( .a(n_25353), .o(FE_OCPN1258_n_25353) );
in01f80 g779241 ( .a(n_1835), .o(n_1836) );
oa22f80 FE_RC_586_0 ( .a(n_32975), .b(n_33428), .c(n_32974), .d(n_33427), .o(n_33503) );
in01f80 FE_OCP_RBC1335_n_20941 ( .a(n_20941), .o(FE_OCP_RBN1335_n_20941) );
oa22f80 FE_RC_1427_0 ( .a(n_22801), .b(n_22701), .c(n_22580), .d(n_22622), .o(n_22742) );
in01f80 g765988 ( .a(n_14721), .o(n_14746) );
in01f80 g755365 ( .a(n_24787), .o(n_24836) );
ao12f80 g778636 ( .a(n_2660), .b(n_3029), .c(n_2611), .o(n_3453) );
no02f80 g775080 ( .a(n_5948), .b(n_5986), .o(n_6037) );
ao12f80 g752155 ( .a(n_28039), .b(FE_OCP_RBN2126_n_44734), .c(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .o(n_28062) );
no02f80 g748831 ( .a(n_31036), .b(n_31086), .o(n_31139) );
no02f80 g774091 ( .a(n_6798), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_), .o(n_6885) );
in01f80 FE_RC_1078_0 ( .a(FE_RN_320_0), .o(n_12579) );
na02f80 g742083 ( .a(FE_OCP_RBN3442_n_37945), .b(n_37392), .o(n_38237) );
no02f80 g781129 ( .a(n_222), .b(n_217), .o(n_218) );
in01f80 g763126 ( .a(n_17862), .o(n_17903) );
in01f80 g776626 ( .a(n_4166), .o(n_4167) );
no02f80 g750079 ( .a(n_29869), .b(n_29417), .o(n_30294) );
oa12f80 g772984 ( .a(n_7797), .b(n_7796), .c(n_7795), .o(n_7934) );
in01f80 g763914 ( .a(n_17159), .o(n_17099) );
in01f80 g739118 ( .a(n_41048), .o(n_41029) );
na02f80 g766887 ( .a(n_14303), .b(n_14215), .o(n_14339) );
na02f80 g776343 ( .a(n_4672), .b(n_4750), .o(n_4880) );
oa12f80 g760561 ( .a(n_20330), .b(n_20329), .c(n_20328), .o(n_21294) );
na02f80 g761139 ( .a(n_19150), .b(n_18742), .o(n_19210) );
na02f80 g761660 ( .a(n_18717), .b(n_18277), .o(n_18796) );
in01f80 newInst_540 ( .a(newNet_503), .o(newNet_540) );
no02f80 g741964 ( .a(n_38042), .b(n_38229), .o(n_38260) );
in01f80 g759866 ( .a(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24624) );
na02f80 g738295 ( .a(n_41888), .b(n_41887), .o(n_41889) );
no02f80 g746941 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_11_), .o(n_33225) );
na02f80 g754506 ( .a(n_26452), .b(n_26415), .o(n_26453) );
oa12f80 g742167 ( .a(n_38306), .b(FE_OCP_RBN2241_n_44881), .c(n_37620), .o(n_38490) );
na02f80 g744028 ( .a(n_44256), .b(n_34263), .o(n_35707) );
na02f80 g784402 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .o(n_46214) );
in01f80 FE_RC_1049_0 ( .a(n_14619), .o(FE_RN_306_0) );
no02f80 g759685 ( .a(n_21722), .b(n_21672), .o(n_21723) );
na02f80 g767865 ( .a(n_12728), .b(delay_add_ln22_unr8_stage4_stallmux_q_21_), .o(n_12836) );
ao22s80 FE_RC_3232_0 ( .a(n_19889), .b(n_19998), .c(n_19863), .d(n_19997), .o(n_20070) );
na02f80 FE_RC_2282_0 ( .a(FE_RN_852_0), .b(n_28539), .o(FE_RN_853_0) );
na02f80 FE_RC_849_0 ( .a(n_29479), .b(n_29480), .o(FE_RN_253_0) );
ao12f80 g762809 ( .a(n_17388), .b(n_17694), .c(n_17035), .o(n_17695) );
na02f80 g769077 ( .a(n_45301), .b(n_11451), .o(n_11519) );
no02f80 g780571 ( .a(n_713), .b(n_757), .o(n_818) );
in01f80 FE_OFC775_n_46137 ( .a(FE_OFN773_n_46137), .o(FE_OFN775_n_46137) );
ao12f80 g749094 ( .a(n_30741), .b(n_30773), .c(FE_OCPN1786_n_30134), .o(n_30885) );
na02f80 g769568 ( .a(n_11424), .b(n_11395), .o(n_11429) );
in01f80 newInst_1211 ( .a(newNet_1210), .o(newNet_1211) );
no02f80 g750816 ( .a(n_29062), .b(n_25738), .o(n_29096) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_21_ ( .ck(newNet_2557), .d(n_27655), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_) );
no02f80 g764818 ( .a(n_15627), .b(n_15622), .o(n_15701) );
no02f80 g739427 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .o(n_40724) );
ao12f80 g745987 ( .a(n_34032), .b(n_33978), .c(n_33940), .o(n_34048) );
oa12f80 g766811 ( .a(n_13704), .b(n_13743), .c(n_13800), .o(n_13803) );
in01f80 g751240 ( .a(n_29944), .o(n_30097) );
oa22f80 FE_RC_1183_0 ( .a(FE_OFN803_n_46285), .b(n_12211), .c(FE_OFN771_n_46337), .d(n_12151), .o(n_46342) );
in01f80 g755175 ( .a(n_25069), .o(n_25070) );
na02f80 g743831 ( .a(n_37190), .b(n_37021), .o(n_37191) );
na02f80 g761288 ( .a(n_19034), .b(n_18550), .o(n_19080) );
in01f80 newInst_1048 ( .a(newNet_899), .o(newNet_1048) );
na02f80 g761328 ( .a(n_19849), .b(n_19763), .o(n_20355) );
in01f80 newInst_3242 ( .a(newNet_3241), .o(newNet_3242) );
no02f80 g738953 ( .a(n_41226), .b(n_41225), .o(n_41227) );
in01f80 g761212 ( .a(n_19135), .o(n_19136) );
in01f80 newInst_693 ( .a(newNet_692), .o(newNet_693) );
na02f80 g749030 ( .a(n_31022), .b(n_30992), .o(n_31077) );
in01f80 FE_OCP_RBC1677_n_44847 ( .a(n_44847), .o(FE_OCP_RBN1677_n_44847) );
in01f80 FE_OCP_RBC2176_n_1864 ( .a(n_1864), .o(FE_OCP_RBN2176_n_1864) );
ao22s80 FE_RC_1339_0 ( .a(FE_OCPN960_n_3951), .b(FE_OCP_RBN2818_n_4458), .c(FE_OCP_RBN2691_FE_OCPN843_n_3912), .d(n_4458), .o(n_4654) );
in01f80 newInst_173 ( .a(newNet_25), .o(newNet_173) );
in01f80 FE_OCP_RBC2811_n_15433 ( .a(FE_OCP_RBN2810_n_15433), .o(FE_OCP_RBN2811_n_15433) );
in01f80 g765610 ( .a(n_15021), .o(n_15156) );
oa22f80 FE_RC_3970_0 ( .a(n_13497), .b(n_13555), .c(n_13554), .d(n_13562), .o(n_13647) );
ao12f80 g779484 ( .a(n_1695), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .o(n_1923) );
in01f80 FE_OCP_RBC3284_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3284_n_44365) );
oa22f80 g752851 ( .a(n_27164), .b(n_27923), .c(n_27948), .d(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(n_28434) );
in01f80 g769941 ( .a(n_11156), .o(n_11157) );
in01f80 g773777 ( .a(n_7270), .o(n_7280) );
in01f80 g771471 ( .a(n_9603), .o(n_9604) );
in01f80 FE_OCP_RBC1989_delay_xor_ln23_unr6_stage3_stallmux_q ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .o(FE_OCP_RBN1989_delay_xor_ln23_unr6_stage3_stallmux_q) );
ao22s80 g736600 ( .a(n_43238), .b(n_43596), .c(n_43239), .d(n_43595), .o(n_43655) );
in01f80 g752502 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_20_), .o(n_27669) );
na02f80 g753883 ( .a(n_27031), .b(n_26886), .o(n_27053) );
no02f80 g760567 ( .a(n_19841), .b(n_19736), .o(n_19924) );
na02f80 g745634 ( .a(n_35479), .b(n_35478), .o(n_35480) );
na02f80 g740372 ( .a(n_39793), .b(n_39112), .o(n_39807) );
no02f80 g768790 ( .a(n_12021), .b(delay_add_ln22_unr8_stage4_stallmux_q_3_), .o(n_12041) );
no02f80 g778536 ( .a(n_2937), .b(n_2842), .o(n_3448) );
na02f80 g776218 ( .a(n_4535), .b(n_4666), .o(n_4620) );
in01f80 FE_RC_2116_0 ( .a(n_24341), .o(FE_RN_734_0) );
na02f80 g737196 ( .a(FE_OCP_RBN3001_n_42959), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_42988) );
oa12f80 g766912 ( .a(n_12683), .b(n_13459), .c(n_12658), .o(n_13560) );
in01f80 g772870 ( .a(n_8024), .o(n_8025) );
oa12f80 g738125 ( .a(n_42024), .b(n_42031), .c(n_42023), .o(n_42052) );
no03m80 g752158 ( .a(n_28215), .b(n_28634), .c(n_28326), .o(n_28688) );
in01f80 g744147 ( .a(n_36004), .o(n_36005) );
no02f80 g750679 ( .a(n_29390), .b(n_29412), .o(n_30703) );
no02f80 g770368 ( .a(n_10536), .b(n_10547), .o(n_10615) );
in01f80 FE_OCP_RBC2653_n_14684 ( .a(n_14684), .o(FE_OCP_RBN2653_n_14684) );
no02f80 FE_RC_314_0 ( .a(FE_RN_93_0), .b(FE_RN_94_0), .o(FE_RN_95_0) );
na02f80 g744012 ( .a(n_36298), .b(n_36267), .o(n_36361) );
in01f80 newInst_1969 ( .a(newNet_276), .o(newNet_1969) );
no02f80 g750593 ( .a(n_29329), .b(n_28848), .o(n_29405) );
in01f80 g776258 ( .a(n_4782), .o(n_4783) );
in01f80 g778011 ( .a(n_3030), .o(n_3069) );
in01f80 FE_RC_2773_0 ( .a(FE_RN_1182_0), .o(n_9077) );
in01f80 g756010 ( .a(n_25140), .o(n_25141) );
na02f80 g776591 ( .a(n_4518), .b(n_4553), .o(n_4519) );
in01f80 g752230 ( .a(n_27941), .o(n_27942) );
na02f80 g739314 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_26_), .o(n_40887) );
ao12f80 g777011 ( .a(n_2728), .b(n_3635), .c(n_2790), .o(n_3636) );
in01f80 g746596 ( .a(n_34740), .o(n_34692) );
in01f80 g744374 ( .a(n_46214), .o(n_36811) );
in01f80 g758960 ( .a(n_21360), .o(n_22331) );
in01f80 newInst_1006 ( .a(newNet_1005), .o(newNet_1006) );
no02f80 g738694 ( .a(n_41716), .b(n_41438), .o(n_41807) );
in01f80 g742918 ( .a(n_37118), .o(n_37119) );
no02f80 g758925 ( .a(n_21605), .b(n_21495), .o(n_21646) );
no02f80 FE_RC_2264_0 ( .a(FE_RN_836_0), .b(FE_RN_839_0), .o(FE_RN_840_0) );
no02f80 g769036 ( .a(FE_OCP_RBN3267_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_4_), .o(n_11918) );
in01f80 g770881 ( .a(n_10053), .o(n_10054) );
na02f80 g760733 ( .a(n_19605), .b(n_18099), .o(n_19704) );
in01f80 FE_OCP_RBC3590_n_47014 ( .a(FE_OCP_RBN3589_n_47014), .o(FE_OCP_RBN3590_n_47014) );
oa12f80 g739126 ( .a(n_40933), .b(n_40964), .c(n_40902), .o(n_40999) );
na02f80 FE_RC_71_0 ( .a(FE_RN_20_0), .b(n_18433), .o(n_18645) );
oa12f80 g737551 ( .a(n_42373), .b(n_42398), .c(n_42387), .o(n_42472) );
oa22f80 FE_RC_605_0 ( .a(n_34304), .b(n_34729), .c(n_34305), .d(n_34715), .o(n_34836) );
ao12f80 g746523 ( .a(n_34473), .b(n_34644), .c(n_34643), .o(n_34668) );
in01f80 g773245 ( .a(n_7605), .o(n_7606) );
in01f80 g751297 ( .a(n_30083), .o(n_29691) );
in01f80 newInst_3589 ( .a(newNet_3588), .o(newNet_3589) );
in01f80 g773401 ( .a(n_7621), .o(n_7622) );
in01f80 g775104 ( .a(n_6067), .o(n_6068) );
in01f80 g774846 ( .a(n_6238), .o(n_6239) );
no02f80 g774964 ( .a(n_6165), .b(FE_OCP_RBN2931_n_5307), .o(n_6198) );
in01f80 newInst_168 ( .a(newNet_167), .o(newNet_168) );
na02f80 g740496 ( .a(n_39736), .b(n_39749), .o(n_39793) );
in01f80 g752592 ( .a(n_27665), .o(n_27644) );
na02f80 g781230 ( .a(n_103), .b(beta_31), .o(n_85) );
in01f80 g752118 ( .a(n_28939), .o(n_28689) );
in01f80 g761469 ( .a(n_20196), .o(n_20197) );
no02f80 g774820 ( .a(n_6240), .b(n_6191), .o(n_6241) );
ao12f80 g752215 ( .a(n_28238), .b(n_28538), .c(n_28154), .o(n_28620) );
na02f80 g746960 ( .a(FE_OCP_RBN2169_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n_33210) );
no02f80 g776319 ( .a(n_4771), .b(n_4310), .o(n_4811) );
na02f80 g761008 ( .a(n_19219), .b(n_19170), .o(n_19430) );
na02f80 g770494 ( .a(n_10474), .b(n_10433), .o(n_10475) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_31_ ( .ck(newNet_3491), .d(n_22897), .o(delay_add_ln22_unr14_stage6_stallmux_q_31_) );
no02f80 g776907 ( .a(n_3718), .b(n_3029), .o(n_3739) );
ao22s80 FE_RC_3791_0 ( .a(n_44365), .b(n_16891), .c(delay_xor_ln22_unr12_stage5_stallmux_q_2_), .d(FE_OCP_RBN3206_n_44365), .o(n_16970) );
in01f80 g747338 ( .a(n_32551), .o(n_32552) );
no02f80 g754203 ( .a(n_25968), .b(n_25991), .o(n_26118) );
in01f80 g751710 ( .a(n_28415), .o(n_28416) );
na02f80 FE_RC_4034_0 ( .a(n_45026), .b(n_22251), .o(FE_RN_1752_0) );
in01f80 fopt783256 ( .a(n_6720), .o(n_44823) );
na02f80 g740325 ( .a(n_40270), .b(n_39915), .o(n_40396) );
in01f80 g779575 ( .a(n_1467), .o(n_1421) );
na02f80 g780581 ( .a(n_745), .b(n_744), .o(n_814) );
in01f80 g743728 ( .a(n_36343), .o(n_36344) );
na02f80 g758516 ( .a(n_21940), .b(n_21954), .o(n_21971) );
na02f80 g775588 ( .a(n_5783), .b(n_5728), .o(n_5791) );
in01f80 g762234 ( .a(n_18187), .o(n_18214) );
in01f80 newInst_3707 ( .a(newNet_2942), .o(newNet_3707) );
in01f80 g754425 ( .a(n_25731), .o(n_25757) );
na02f80 g775450 ( .a(n_5642), .b(n_5719), .o(n_5730) );
in01f80 g750628 ( .a(n_29441), .o(n_31045) );
no02f80 g740142 ( .a(n_39816), .b(n_39817), .o(n_39818) );
in01f80 g757831 ( .a(n_22553), .o(n_22569) );
no02f80 g760376 ( .a(n_20150), .b(n_20063), .o(n_20207) );
in01f80 FE_RC_1739_0 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(FE_RN_486_0) );
ao12f80 g760670 ( .a(n_19743), .b(n_19742), .c(FE_OCP_RBN3842_n_19555), .o(n_21434) );
in01f80 g775845 ( .a(n_4907), .o(n_4964) );
in01f80 g769624 ( .a(n_11349), .o(n_11350) );
in01f80 FE_OCPC1757_n_33213 ( .a(n_33213), .o(FE_OCPN1757_n_33213) );
in01f80 FE_OCP_RBC2306_n_24288 ( .a(n_24288), .o(FE_OCP_RBN2306_n_24288) );
in01f80 g747808 ( .a(n_33624), .o(n_33625) );
in01f80 newInst_808 ( .a(newNet_396), .o(newNet_808) );
ao22s80 g757079 ( .a(n_23523), .b(n_23148), .c(n_23524), .d(n_23149), .o(n_23810) );
na02f80 g736956 ( .a(n_43242), .b(n_42714), .o(n_43518) );
no02f80 g779606 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .o(n_1832) );
in01f80 FE_OCPC1012_n_41478 ( .a(n_41478), .o(FE_OCPN1012_n_41478) );
oa12f80 g751025 ( .a(n_30097), .b(n_30096), .c(n_30095), .o(n_30208) );
na02f80 g766286 ( .a(n_14200), .b(n_14117), .o(n_14285) );
oa12f80 g769983 ( .a(n_10082), .b(n_11057), .c(FE_OCPN1388_n_11041), .o(n_11042) );
na02f80 g738264 ( .a(n_41919), .b(n_41918), .o(n_41920) );
in01f80 newInst_3099 ( .a(newNet_3098), .o(newNet_3099) );
in01f80 g758565 ( .a(n_22604), .o(n_22605) );
in01f80 FE_OCP_RBC2459_n_13765 ( .a(FE_OCP_RBN2456_n_13765), .o(FE_OCP_RBN2459_n_13765) );
ao12f80 g742938 ( .a(n_36999), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n_37061) );
na02f80 g776483 ( .a(n_4253), .b(n_3082), .o(n_4457) );
in01f80 fopt782836 ( .a(n_34890), .o(n_44262) );
ao12f80 g746513 ( .a(n_34443), .b(n_34442), .c(n_34441), .o(n_34891) );
ao22s80 FE_RC_4140_0 ( .a(n_45224), .b(n_11696), .c(FE_RN_1798_0), .d(delay_xor_ln22_unr9_stage4_stallmux_q_2_), .o(n_11734) );
na02f80 FE_RC_2927_0 ( .a(n_27210), .b(n_27211), .o(FE_RN_1275_0) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_0_ ( .ck(newNet_682), .d(n_46381), .o(delay_xor_ln21_unr9_stage4_stallmux_q_0_) );
ao12f80 g746499 ( .a(n_33082), .b(n_33306), .c(n_33106), .o(n_33330) );
in01f80 FE_OCP_RBC3655_n_15097 ( .a(n_15097), .o(FE_OCP_RBN3655_n_15097) );
ao12f80 g766305 ( .a(n_14214), .b(n_14703), .c(n_14136), .o(n_14731) );
na02f80 g777055 ( .a(n_3750), .b(n_4905), .o(n_3804) );
in01f80 newInst_1385 ( .a(newNet_1384), .o(newNet_1385) );
ao12f80 g772486 ( .a(n_8650), .b(n_8649), .c(n_8648), .o(n_9631) );
na02f80 g778364 ( .a(n_2787), .b(n_2115), .o(n_2910) );
na02f80 g744492 ( .a(n_35456), .b(n_35467), .o(n_35457) );
na02f80 g737893 ( .a(n_42201), .b(n_42350), .o(n_42384) );
no02f80 g771590 ( .a(n_8953), .b(n_8309), .o(n_8989) );
no02f80 g760925 ( .a(n_19446), .b(FE_OCPN1800_FE_OFN780_n_17093), .o(n_19552) );
in01f80 g775982 ( .a(n_5274), .o(n_5275) );
na02f80 g763338 ( .a(n_17185), .b(n_17223), .o(n_17380) );
in01f80 g758864 ( .a(n_21679), .o(n_21612) );
na02f80 FE_RC_3683_0 ( .a(FE_RN_1616_0), .b(FE_RN_1617_0), .o(FE_RN_1618_0) );
no02f80 FE_RC_1402_0 ( .a(FE_RN_408_0), .b(FE_RN_409_0), .o(FE_RN_410_0) );
no02f80 g772602 ( .a(n_8390), .b(n_8389), .o(n_8423) );
no02f80 g740585 ( .a(n_39595), .b(n_39606), .o(n_39629) );
in01f80 g751122 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30588) );
in01f80 g765939 ( .a(n_14794), .o(n_14815) );
ao12f80 g767234 ( .a(n_13157), .b(n_13716), .c(n_13284), .o(n_13767) );
na02f80 g749592 ( .a(n_30374), .b(n_30020), .o(n_30489) );
na02f80 g750562 ( .a(n_29381), .b(n_29270), .o(n_29451) );
no02f80 g759366 ( .a(n_20918), .b(n_20956), .o(n_21042) );
oa12f80 g756441 ( .a(n_23599), .b(n_23740), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n_23741) );
no02f80 g759709 ( .a(n_20418), .b(n_45060), .o(n_20480) );
no02f80 g740942 ( .a(n_39110), .b(n_39015), .o(n_39145) );
no02f80 g753098 ( .a(FE_OCPN1750_n_27223), .b(n_27178), .o(n_27398) );
no02f80 g770156 ( .a(n_10903), .b(n_10871), .o(n_10920) );
no02f80 g747791 ( .a(n_33372), .b(n_33336), .o(n_33884) );
in01f80 g766408 ( .a(n_14273), .o(n_14317) );
no02f80 g770031 ( .a(n_10797), .b(n_44464), .o(n_10826) );
oa22f80 FE_RC_1223_0 ( .a(n_6489), .b(n_6398), .c(n_6399), .d(n_6499), .o(n_6643) );
no02f80 g771218 ( .a(n_9535), .b(FE_OCP_RBN3572_n_44563), .o(n_9556) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_0_ ( .ck(newNet_425), .d(n_32431), .o(delay_xor_ln22_unr21_stage8_stallmux_q_0_) );
in01f80 FE_OFC5_n_43918 ( .a(FE_OFN0_n_43918), .o(FE_OFN5_n_43918) );
oa22f80 FE_RC_388_0 ( .a(n_1018), .b(n_44652), .c(n_975), .d(n_44637), .o(n_1345) );
na02f80 g776864 ( .a(n_3684), .b(n_2894), .o(n_3736) );
na02f80 g760812 ( .a(n_20121), .b(n_20120), .o(n_20122) );
in01f80 g772662 ( .a(n_46418), .o(n_8367) );
no02f80 g762350 ( .a(n_45002), .b(n_18521), .o(n_18835) );
no02f80 g767350 ( .a(n_13446), .b(n_13453), .o(n_13482) );
oa12f80 g764349 ( .a(n_16314), .b(n_16361), .c(n_16422), .o(n_16452) );
in01f80 newInst_415 ( .a(newNet_3), .o(newNet_415) );
in01f80 FE_OCP_RBC2120_n_45224 ( .a(FE_OCP_RBN2118_n_45224), .o(FE_OCP_RBN2120_n_45224) );
oa22f80 g764124 ( .a(n_16601), .b(n_17584), .c(n_16578), .d(n_16338), .o(n_16636) );
no02f80 g745952 ( .a(n_34064), .b(n_33961), .o(n_34078) );
no02f80 g750979 ( .a(n_29856), .b(n_30129), .o(n_30130) );
no02f80 g776791 ( .a(n_47010), .b(n_4231), .o(n_4331) );
in01f80 g784792 ( .a(n_47332), .o(n_47333) );
ao12f80 g770913 ( .a(n_9481), .b(n_10131), .c(n_9548), .o(n_10255) );
in01f80 newInst_1170 ( .a(newNet_1169), .o(newNet_1170) );
na02f80 FE_RC_2161_0 ( .a(n_14452), .b(FE_OCP_RBN2810_n_15433), .o(FE_RN_766_0) );
no02f80 g766489 ( .a(n_13995), .b(n_13029), .o(n_14030) );
no02f80 g742993 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .b(delay_add_ln22_unr23_stage9_stallmux_q_7_), .o(n_36966) );
na02f80 g760963 ( .a(n_19223), .b(n_19222), .o(n_19286) );
in01f80 g779778 ( .a(n_1423), .o(n_1471) );
in01f80 newInst_2196 ( .a(newNet_2195), .o(newNet_2196) );
oa12f80 g745204 ( .a(n_34208), .b(n_34415), .c(n_34188), .o(n_34440) );
in01f80 FE_OCPC984_n_25210 ( .a(n_25210), .o(FE_OCPN984_n_25210) );
in01f80 g755998 ( .a(n_25521), .o(n_25522) );
ao12f80 g758874 ( .a(n_21518), .b(n_22030), .c(n_21483), .o(n_22117) );
na02f80 g740153 ( .a(n_39781), .b(n_39841), .o(n_39918) );
in01f80 newInst_1839 ( .a(newNet_252), .o(newNet_1839) );
na02f80 g742084 ( .a(n_37945), .b(n_37309), .o(n_38283) );
oa22f80 g757616 ( .a(n_22709), .b(n_22801), .c(n_22666), .d(n_22793), .o(n_22766) );
in01f80 newInst_2125 ( .a(newNet_851), .o(newNet_2125) );
oa22f80 g784377 ( .a(n_6500), .b(FE_OFN806_n_46196), .c(n_6490), .d(FE_OFN84_n_46137), .o(n_46183) );
no02f80 g778588 ( .a(n_2661), .b(n_2660), .o(n_2662) );
in01f80 newInst_874 ( .a(newNet_313), .o(newNet_874) );
na02f80 g784757 ( .a(n_8889), .b(n_47239), .o(n_47243) );
no02f80 g747193 ( .a(n_32758), .b(FE_OCP_RBN1339_n_32653), .o(n_32759) );
in01f80 FE_OCP_RBC2651_n_9030 ( .a(n_9030), .o(FE_OCP_RBN2651_n_9030) );
in01f80 g778405 ( .a(n_3217), .o(n_3178) );
in01f80 g736473 ( .a(n_43726), .o(n_43727) );
in01f80 newInst_314 ( .a(newNet_313), .o(newNet_314) );
na02f80 g746385 ( .a(n_33486), .b(n_33485), .o(n_33487) );
ao12f80 g739254 ( .a(n_40786), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_21_), .o(n_41079) );
oa12f80 g749342 ( .a(n_31122), .b(n_30693), .c(n_29229), .o(n_30813) );
na02f80 FE_RC_268_0 ( .a(FE_OCP_RBN1369_n_20763), .b(FE_OCP_RBN3853_n_20848), .o(FE_RN_80_0) );
ao22s80 g737211 ( .a(n_42938), .b(n_42354), .c(n_42927), .d(n_42353), .o(n_42992) );
na02f80 g771032 ( .a(n_9887), .b(n_9922), .o(n_10040) );
in01f80 g763918 ( .a(n_17297), .o(n_17298) );
in01f80 g736810 ( .a(n_43089), .o(n_43090) );
in01f80 g750024 ( .a(n_30401), .o(n_30402) );
na02f80 g779076 ( .a(n_2060), .b(n_2081), .o(n_2427) );
no02f80 g771760 ( .a(FE_OCP_RBN3547_n_44575), .b(n_9001), .o(n_9168) );
in01f80 g754844 ( .a(n_25487), .o(n_25488) );
na02f80 g749298 ( .a(n_30626), .b(FE_OCPN1410_n_27014), .o(n_30656) );
no02f80 g746117 ( .a(n_33847), .b(FE_RN_1821_0), .o(n_33875) );
in01f80 g766480 ( .a(n_14069), .o(n_14070) );
no02f80 g764796 ( .a(n_15756), .b(n_13880), .o(n_15937) );
na02f80 g762310 ( .a(n_18090), .b(n_17944), .o(n_18094) );
in01f80 FE_OCP_RBC3586_n_25295 ( .a(n_25295), .o(FE_OCP_RBN3586_n_25295) );
oa22f80 g763779 ( .a(n_16686), .b(FE_OFN767_n_15670), .c(n_16658), .d(n_16339), .o(n_16730) );
oa22f80 g739806 ( .a(n_40429), .b(n_40358), .c(n_40430), .d(n_40357), .o(n_40469) );
in01f80 g743760 ( .a(n_36309), .o(n_36372) );
in01f80 g757407 ( .a(n_22992), .o(n_22993) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_27_ ( .ck(newNet_3212), .d(n_36632), .o(delay_add_ln22_unr23_stage9_stallmux_q_27_) );
in01f80 g772282 ( .a(n_8733), .o(n_8734) );
in01f80 FE_OCP_RBC2158_n_1614 ( .a(n_1614), .o(FE_OCP_RBN2158_n_1614) );
no03m80 FE_RC_3685_0 ( .a(n_1542), .b(n_1547), .c(n_1380), .o(n_1602) );
in01f80 FE_OCPC1792_n_25044 ( .a(FE_OCPN1791_n_25044), .o(FE_OCPN1792_n_25044) );
oa22f80 FE_RC_385_0 ( .a(n_928), .b(FE_OCPN874_n_44672), .c(n_875), .d(n_44637), .o(n_1316) );
no03m80 g766806 ( .a(n_14455), .b(n_14421), .c(n_14491), .o(n_14492) );
no02f80 g748035 ( .a(n_44347), .b(n_32502), .o(n_33000) );
na02f80 g744734 ( .a(n_35177), .b(n_35148), .o(n_35201) );
no02f80 g774777 ( .a(n_6415), .b(n_6330), .o(n_6442) );
in01f80 FE_OCP_RBC2422_n_24501 ( .a(n_24501), .o(FE_OCP_RBN2422_n_24501) );
no02f80 g739157 ( .a(n_40914), .b(n_40748), .o(n_40943) );
in01f80 g736545 ( .a(n_43639), .o(n_43640) );
oa22f80 g779879 ( .a(n_44652), .b(n_1152), .c(n_44623), .d(n_1138), .o(n_1311) );
no02f80 g755417 ( .a(n_24700), .b(n_24728), .o(n_24839) );
ao12f80 g773824 ( .a(n_7114), .b(n_7118), .c(n_7113), .o(n_7182) );
no02f80 g764934 ( .a(n_15542), .b(n_15501), .o(n_15687) );
ao12f80 g744856 ( .a(n_36419), .b(n_36420), .c(n_35797), .o(n_36464) );
no02f80 g768839 ( .a(n_12036), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n_11996) );
in01f80 newInst_94 ( .a(newNet_93), .o(newNet_94) );
na02f80 g741580 ( .a(n_38669), .b(n_37636), .o(n_38766) );
ao12f80 g784662 ( .a(n_7490), .b(n_7462), .c(n_7292), .o(n_46992) );
in01f80 g743279 ( .a(n_36789), .o(n_36798) );
na02f80 g775234 ( .a(n_5944), .b(n_4973), .o(n_5994) );
in01f80 g755907 ( .a(n_25710), .o(n_25711) );
ao12f80 g778152 ( .a(n_2716), .b(n_2715), .c(n_2714), .o(n_4136) );
na02f80 g773588 ( .a(n_7425), .b(n_7424), .o(n_7472) );
in01f80 g771048 ( .a(n_9456), .o(n_9472) );
in01f80 fopt783566 ( .a(n_34768), .o(n_45185) );
ao12f80 g765958 ( .a(n_15064), .b(n_15090), .c(n_15063), .o(n_15712) );
in01f80 FE_OCP_RBC2111_n_11548 ( .a(n_11548), .o(FE_OCP_RBN2111_n_11548) );
ao22s80 g751506 ( .a(n_28597), .b(n_28541), .c(n_28458), .d(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n_28674) );
in01f80 g769361 ( .a(n_11892), .o(n_12014) );
in01f80 FE_OCP_RBC2137_n_11907 ( .a(n_11907), .o(FE_OCP_RBN2137_n_11907) );
na02f80 g744793 ( .a(n_35116), .b(n_30545), .o(n_35174) );
in01f80 newInst_3295 ( .a(newNet_3294), .o(newNet_3295) );
in01f80 g775461 ( .a(n_5897), .o(n_5898) );
ao12f80 g766258 ( .a(n_14757), .b(n_14780), .c(n_14756), .o(n_15747) );
no02f80 g767499 ( .a(n_13143), .b(n_13227), .o(n_13296) );
in01f80 g755943 ( .a(n_24274), .o(n_24268) );
in01f80 g753737 ( .a(n_26524), .o(n_26555) );
no02f80 g763061 ( .a(n_17620), .b(delay_add_ln22_unr11_stage5_stallmux_q_5_), .o(n_17639) );
na02f80 g743702 ( .a(n_36343), .b(n_35831), .o(n_36375) );
ao12f80 g751319 ( .a(n_28659), .b(n_28684), .c(n_28658), .o(n_29860) );
no02f80 g767654 ( .a(n_12865), .b(n_12801), .o(n_12879) );
na02f80 g776222 ( .a(n_4666), .b(n_4665), .o(n_4741) );
in01f80 newInst_2493 ( .a(newNet_2492), .o(newNet_2493) );
in01f80 FE_OCP_DRV_C1539_n_35427 ( .a(n_35427), .o(FE_OCP_DRV_N1539_n_35427) );
in01f80 g741223 ( .a(n_39320), .o(n_39321) );
na02f80 g759949 ( .a(n_21374), .b(n_21593), .o(n_21692) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_0_ ( .ck(newNet_2130), .d(n_4157), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_) );
no02f80 g758043 ( .a(n_22692), .b(n_22695), .o(n_22696) );
oa22f80 g772216 ( .a(n_8654), .b(n_8536), .c(n_8653), .d(n_8570), .o(n_8781) );
in01f80 g774066 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_30_), .o(n_6681) );
na02f80 g757692 ( .a(FE_OCP_RBN3817_n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_1_), .o(n_22615) );
in01f80 g768341 ( .a(n_12592), .o(n_12593) );
na02f80 g775429 ( .a(n_5730), .b(n_5771), .o(n_5909) );
no02f80 g760247 ( .a(FE_OCP_RBN3617_n_20249), .b(n_19454), .o(n_20605) );
na02f80 g766095 ( .a(n_14517), .b(n_14557), .o(n_14638) );
in01f80 newInst_2031 ( .a(newNet_1058), .o(newNet_2031) );
na02f80 g742117 ( .a(n_38135), .b(n_38134), .o(n_38158) );
no02f80 g746923 ( .a(FE_OCP_RBN3390_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(n_33449) );
in01f80 g762352 ( .a(n_18449), .o(n_18450) );
ao12f80 g765020 ( .a(n_15380), .b(n_15460), .c(n_15532), .o(n_15498) );
na02f80 g751569 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .o(n_28784) );
in01f80 g754379 ( .a(FE_OCP_RBN2814_n_25817), .o(n_25873) );
na02f80 g762404 ( .a(FE_OFN751_n_45003), .b(n_18103), .o(n_18729) );
in01f80 g780497 ( .a(n_1043), .o(n_1044) );
in01f80 g747385 ( .a(n_32547), .o(n_32548) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_22_ ( .ck(newNet_3415), .d(n_27727), .o(delay_add_ln22_unr17_stage7_stallmux_q_22_) );
no02f80 g741519 ( .a(n_38707), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38708) );
in01f80 g744204 ( .a(n_36258), .o(n_36259) );
oa22f80 FE_RC_3888_0 ( .a(n_32575), .b(n_32523), .c(n_32601), .d(n_32576), .o(n_32655) );
na02f80 g761072 ( .a(n_19064), .b(n_17881), .o(n_19089) );
in01f80 g750631 ( .a(n_29399), .o(n_29400) );
in01f80 g744474 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_23_), .o(n_36762) );
na02f80 g740172 ( .a(FE_OCP_RBN3056_n_39913), .b(n_46948), .o(n_40037) );
in01f80 FE_RC_3639_0 ( .a(FE_RN_1596_0), .o(FE_RN_1594_0) );
no02f80 g778034 ( .a(n_3085), .b(n_3084), .o(n_3140) );
na03f80 FE_RC_1148_0 ( .a(n_37353), .b(n_37366), .c(n_37357), .o(n_37373) );
oa22f80 FE_RC_3290_0 ( .a(n_31827), .b(n_32220), .c(n_31828), .d(n_32219), .o(n_32310) );
in01f80 g764626 ( .a(n_15818), .o(n_15819) );
no02f80 g760728 ( .a(n_19597), .b(FE_OCP_RBN1349_n_19270), .o(n_19659) );
in01f80 g780771 ( .a(n_490), .o(n_558) );
in01f80 newInst_740 ( .a(newNet_285), .o(newNet_740) );
in01f80 newInst_3120 ( .a(newNet_85), .o(newNet_3120) );
na02f80 FE_RC_4149_0 ( .a(FE_RN_1800_0), .b(FE_RN_1804_0), .o(n_17194) );
na02f80 g758107 ( .a(n_44267), .b(FE_OCP_RBN1338_n_20941), .o(n_22300) );
ao12f80 g755550 ( .a(n_24716), .b(n_24715), .c(n_24714), .o(n_26428) );
no02f80 g773910 ( .a(n_6883), .b(n_6882), .o(n_6884) );
oa12f80 g764329 ( .a(n_16206), .b(n_16234), .c(n_16233), .o(n_16291) );
na02f80 g778082 ( .a(n_3007), .b(n_2979), .o(n_3085) );
no02f80 g775254 ( .a(n_5944), .b(n_5113), .o(n_5945) );
no02f80 g778541 ( .a(n_2321), .b(n_2717), .o(n_2373) );
na02f80 g743138 ( .a(n_36475), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_36983) );
no02f80 g768594 ( .a(n_45659), .b(delay_xor_ln21_unr9_stage4_stallmux_q_15_), .o(n_12323) );
no02f80 g774371 ( .a(n_6641), .b(n_6541), .o(n_7012) );
ao12f80 g771809 ( .a(n_8869), .b(n_8868), .c(n_8867), .o(n_10073) );
in01f80 g767446 ( .a(n_13235), .o(n_13266) );
no02f80 FE_RC_2823_0 ( .a(FE_RN_1211_0), .b(n_34572), .o(FE_RN_1212_0) );
na02f80 g754321 ( .a(FE_OCP_RBN2813_n_25817), .b(n_23354), .o(n_25879) );
no02f80 g742964 ( .a(n_37139), .b(n_37172), .o(n_37821) );
na02f80 g738570 ( .a(n_41616), .b(n_41557), .o(n_41617) );
in01f80 newInst_3545 ( .a(newNet_3544), .o(newNet_3545) );
in01f80 g770104 ( .a(n_10874), .o(n_10889) );
no02f80 g760872 ( .a(n_19438), .b(n_19377), .o(n_19439) );
in01f80 FE_OCP_RBC3496_n_13818 ( .a(FE_OCP_RBN2358_n_13818), .o(FE_OCP_RBN3496_n_13818) );
na02f80 g766058 ( .a(n_14736), .b(n_14681), .o(n_14760) );
no02f80 g778577 ( .a(n_2420), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_), .o(n_2546) );
no02f80 g777691 ( .a(FE_OCP_RBN2560_n_3437), .b(FE_OCP_RBN2464_n_4336), .o(n_3512) );
no02f80 g739946 ( .a(n_40089), .b(n_39957), .o(n_40090) );
in01f80 g742703 ( .a(n_37373), .o(n_37374) );
no02f80 FE_RC_2159_0 ( .a(FE_RN_763_0), .b(FE_RN_764_0), .o(n_15552) );
in01f80 g736650 ( .a(n_43442), .o(n_43412) );
in01f80 newInst_706 ( .a(newNet_705), .o(newNet_706) );
no02f80 g773015 ( .a(n_7713), .b(n_7684), .o(n_7756) );
in01f80 g737561 ( .a(n_42492), .o(n_42529) );
ao12f80 g756827 ( .a(n_23811), .b(n_23724), .c(n_23671), .o(n_23838) );
na02f80 g738593 ( .a(n_41804), .b(n_41850), .o(n_41957) );
in01f80 g776552 ( .a(n_4317), .o(n_4318) );
in01f80 FE_RC_3170_0 ( .a(n_22347), .o(FE_RN_1404_0) );
no02f80 FE_RC_2639_0 ( .a(FE_RN_1100_0), .b(n_2392), .o(n_2433) );
oa12f80 g756070 ( .a(n_24905), .b(n_24904), .c(n_24903), .o(n_24979) );
oa12f80 g736886 ( .a(n_43192), .b(FE_OCP_RBN3074_n_43230), .c(n_43052), .o(n_43595) );
in01f80 g769203 ( .a(n_12048), .o(n_12049) );
na03f80 g761834 ( .a(n_18477), .b(n_47246), .c(n_18440), .o(n_18478) );
oa12f80 g764478 ( .a(n_16574), .b(n_16573), .c(n_16572), .o(n_16616) );
no02f80 g747803 ( .a(n_33191), .b(n_32584), .o(n_33242) );
in01f80 g749744 ( .a(n_31633), .o(n_31634) );
in01f80 FE_OCP_RBC1728_FE_RN_1583_0 ( .a(FE_RN_1583_0), .o(FE_OCP_RBN1728_FE_RN_1583_0) );
no02f80 g749529 ( .a(n_30593), .b(n_30592), .o(n_30594) );
in01f80 g775635 ( .a(FE_OCP_RBN3696_n_5284), .o(n_5320) );
no02f80 FE_RC_273_0 ( .a(FE_RN_81_0), .b(FE_OCP_RBN3064_n_22170), .o(FE_RN_83_0) );
na02f80 g761888 ( .a(n_18440), .b(n_18400), .o(n_18509) );
no02f80 g747212 ( .a(n_32671), .b(n_32670), .o(n_32697) );
in01f80 g778074 ( .a(n_3035), .o(n_3036) );
no02f80 g743306 ( .a(n_36675), .b(n_36750), .o(n_36743) );
no02f80 g748010 ( .a(n_32981), .b(n_33028), .o(n_33070) );
no02f80 g774283 ( .a(n_6684), .b(n_6585), .o(n_6695) );
no02f80 FE_RC_2222_0 ( .a(n_32920), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(FE_RN_805_0) );
in01f80 newInst_758 ( .a(newNet_757), .o(newNet_758) );
in01f80 g762120 ( .a(n_18777), .o(n_18778) );
no02f80 g766555 ( .a(n_14115), .b(n_12868), .o(n_14089) );
in01f80 FE_RC_2386_0 ( .a(n_42423), .o(FE_RN_933_0) );
oa12f80 g758741 ( .a(n_21451), .b(n_22210), .c(n_21697), .o(n_22286) );
na02f80 g773755 ( .a(n_7186), .b(n_7160), .o(n_7244) );
in01f80 g761736 ( .a(n_18746), .o(n_18803) );
na02f80 g746030 ( .a(n_33957), .b(n_33872), .o(n_33960) );
no02f80 g760898 ( .a(n_19459), .b(n_19424), .o(n_20265) );
in01f80 FE_OCP_RBC2815_n_25986 ( .a(n_25986), .o(FE_OCP_RBN2815_n_25986) );
in01f80 FE_OCP_RBC2870_n_10480 ( .a(n_10480), .o(FE_OCP_RBN2870_n_10480) );
no02f80 g763505 ( .a(FE_OCP_RBN3079_n_16977), .b(n_16940), .o(n_17454) );
na02f80 g765671 ( .a(n_15066), .b(n_13478), .o(n_15132) );
no02f80 g775863 ( .a(n_4922), .b(FE_OCP_RBN2728_n_4219), .o(n_5030) );
in01f80 FE_RC_4190_0 ( .a(FE_RN_1835_0), .o(FE_RN_1831_0) );
no02f80 g747261 ( .a(n_33722), .b(n_33394), .o(n_33795) );
in01f80 FE_RC_466_0 ( .a(n_28385), .o(FE_RN_136_0) );
na02f80 g755140 ( .a(n_25551), .b(FE_OCP_RBN2423_n_24501), .o(n_25612) );
na02f80 g761692 ( .a(n_18600), .b(FE_OFN778_n_17093), .o(n_18649) );
oa22f80 FE_RC_3905_0 ( .a(n_45091), .b(FE_OCP_RBN3851_n_20848), .c(n_45013), .d(n_20848), .o(n_21006) );
na02f80 g746612 ( .a(n_34390), .b(n_34389), .o(n_34417) );
na02f80 FE_RC_1143_0 ( .a(FE_OCPN1241_n_7721), .b(n_8077), .o(FE_RN_345_0) );
ao12f80 g743152 ( .a(n_36911), .b(n_36910), .c(n_36909), .o(n_36947) );
in01f80 g769224 ( .a(n_11587), .o(n_11588) );
in01f80 g755336 ( .a(n_24967), .o(n_24968) );
in01f80 g767601 ( .a(n_14153), .o(n_13048) );
in01f80 g765096 ( .a(n_15530), .o(n_15606) );
in01f80 newInst_2600 ( .a(newNet_2599), .o(newNet_2600) );
na02f80 g773229 ( .a(n_7569), .b(n_7557), .o(n_7570) );
in01f80 FE_OCP_RBC2764_n_25732 ( .a(n_25732), .o(FE_OCP_RBN2764_n_25732) );
no02f80 g737173 ( .a(FE_OCP_RBN3032_n_43000), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_43020) );
oa12f80 g760439 ( .a(n_20600), .b(n_20624), .c(n_20599), .o(n_21251) );
no02f80 FE_RC_3594_0 ( .a(FE_RN_1568_0), .b(n_25098), .o(n_25154) );
in01f80 g779019 ( .a(n_2858), .o(n_2102) );
no02f80 g769011 ( .a(n_11530), .b(FE_OCP_RBN3093_n_11475), .o(n_11646) );
oa12f80 g773441 ( .a(n_7584), .b(n_7595), .c(n_7651), .o(n_7678) );
na02f80 g770703 ( .a(n_10220), .b(FE_OCP_RBN2855_n_10112), .o(n_10260) );
no02f80 g737369 ( .a(n_42838), .b(n_42468), .o(n_42854) );
ao12f80 g756178 ( .a(n_22089), .b(n_24157), .c(n_24121), .o(n_24246) );
oa22f80 g784422 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_8_), .c(n_36785), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46234) );
oa12f80 g772973 ( .a(n_7305), .b(n_7662), .c(n_7262), .o(n_7731) );
in01f80 g740631 ( .a(n_39635), .o(n_39636) );
na02f80 g742032 ( .a(n_38000), .b(n_44875), .o(n_38053) );
in01f80 g746004 ( .a(n_34030), .o(n_34031) );
no02f80 g773980 ( .a(n_7172), .b(delay_xor_ln21_unr6_stage3_stallmux_q_23_), .o(n_7254) );
in01f80 g753127 ( .a(n_27500), .o(n_27501) );
oa12f80 g754071 ( .a(n_26092), .b(n_26091), .c(FE_OCPN1530_n_26090), .o(n_26150) );
no02f80 g774350 ( .a(n_6512), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6544) );
in01f80 g773846 ( .a(n_7090), .o(n_7091) );
no02f80 g771893 ( .a(n_8857), .b(n_8805), .o(n_8969) );
na02f80 g745796 ( .a(n_34113), .b(n_34026), .o(n_34147) );
na02f80 g759752 ( .a(n_20636), .b(n_20635), .o(n_20637) );
oa22f80 FE_RC_843_0 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .b(n_42155), .c(n_42196), .d(n_42154), .o(n_42182) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_1_ ( .ck(newNet_2392), .d(n_35378), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_) );
in01f80 g745089 ( .a(n_34795), .o(n_34769) );
in01f80 g743017 ( .a(n_36996), .o(n_36957) );
in01f80 g768510 ( .a(n_12387), .o(n_12388) );
na02f80 g770076 ( .a(n_10940), .b(n_10914), .o(n_10941) );
na02f80 g748936 ( .a(n_31102), .b(n_27315), .o(n_31178) );
no02f80 g751304 ( .a(n_29651), .b(n_29650), .o(n_29652) );
in01f80 g777275 ( .a(n_5111), .o(n_5112) );
in01f80 FE_OCP_RBC3375_n_6822 ( .a(n_6822), .o(FE_OCP_RBN3375_n_6822) );
no02f80 g756754 ( .a(n_24035), .b(n_24032), .o(n_24065) );
ao12f80 g780788 ( .a(n_425), .b(n_420), .c(n_501), .o(n_519) );
ao12f80 g755351 ( .a(n_24788), .b(n_24699), .c(FE_OCPN1482_n_22207), .o(n_24810) );
in01f80 g773163 ( .a(n_7889), .o(n_7829) );
in01f80 newInst_1408 ( .a(newNet_1407), .o(newNet_1408) );
ao12f80 g780849 ( .a(n_463), .b(n_521), .c(n_479), .o(n_652) );
na02f80 g779031 ( .a(n_2119), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_16_), .o(n_2175) );
no02f80 g767000 ( .a(n_13559), .b(FE_OCPN860_n_12880), .o(n_13572) );
in01f80 FE_RC_1135_0 ( .a(FE_OCPN871_n_2737), .o(FE_RN_343_0) );
in01f80 g746545 ( .a(n_34962), .o(n_34963) );
na02f80 g773687 ( .a(n_7336), .b(n_7086), .o(n_7389) );
no02f80 g763005 ( .a(n_17937), .b(n_17359), .o(n_17938) );
na02f80 g771429 ( .a(n_9134), .b(n_8309), .o(n_9253) );
na02f80 g776106 ( .a(n_5007), .b(n_4966), .o(n_5105) );
na02f80 g757649 ( .a(n_22769), .b(n_22634), .o(n_22677) );
no02f80 g751274 ( .a(n_29724), .b(n_29723), .o(n_29725) );
na02f80 g774944 ( .a(n_6194), .b(n_6207), .o(n_6301) );
ao12f80 g780761 ( .a(n_524), .b(n_523), .c(n_522), .o(n_695) );
in01f80 newInst_2868 ( .a(newNet_2867), .o(newNet_2868) );
no02f80 FE_RC_3798_0 ( .a(FE_RN_1658_0), .b(FE_RN_1659_0), .o(FE_RN_1660_0) );
in01f80 g749367 ( .a(n_30758), .o(n_31122) );
in01f80 g761517 ( .a(n_18944), .o(n_18975) );
na02f80 g776068 ( .a(n_5046), .b(n_5064), .o(n_5243) );
na02f80 g750785 ( .a(n_29313), .b(n_29290), .o(n_29291) );
in01f80 g757825 ( .a(n_23698), .o(n_23061) );
ao12f80 g746143 ( .a(n_34670), .b(n_35089), .c(n_34638), .o(n_35163) );
in01f80 FE_OCP_RBC2473_n_8664 ( .a(FE_OCP_RBN2472_n_8664), .o(FE_OCP_RBN2473_n_8664) );
no04s80 g742883 ( .a(n_37293), .b(n_37543), .c(n_45897), .d(n_37247), .o(n_38372) );
in01f80 FE_RC_3771_0 ( .a(n_13418), .o(FE_RN_1655_0) );
oa12f80 g760501 ( .a(n_20000), .b(n_19999), .c(n_20007), .o(n_20059) );
no02f80 g759619 ( .a(n_20759), .b(n_20789), .o(n_20872) );
na02f80 g737037 ( .a(n_43082), .b(n_43130), .o(n_43530) );
no02f80 g736632 ( .a(n_43156), .b(n_43045), .o(n_43157) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_8_ ( .ck(newNet_2800), .d(n_10530), .o(delay_add_ln22_unr8_stage4_stallmux_q_8_) );
na02f80 g751437 ( .a(n_28719), .b(n_28721), .o(n_28725) );
in01f80 g750741 ( .a(n_29340), .o(n_29341) );
na02f80 g738229 ( .a(n_41924), .b(n_41941), .o(n_41942) );
in01f80 g753500 ( .a(n_26848), .o(n_26849) );
oa22f80 FE_RC_3918_0 ( .a(n_22460), .b(n_22743), .c(n_22501), .d(n_22703), .o(n_22903) );
no02f80 FE_RC_2034_0 ( .a(FE_RN_678_0), .b(n_25893), .o(FE_RN_679_0) );
na02f80 g774956 ( .a(n_6118), .b(n_5981), .o(n_6166) );
no02f80 FE_RC_2910_0 ( .a(FE_RN_1264_0), .b(FE_RN_1263_0), .o(FE_RN_1265_0) );
in01f80 FE_RC_4253_0 ( .a(FE_RN_1872_0), .o(n_22065) );
no02f80 g776726 ( .a(n_3894), .b(n_3792), .o(n_3942) );
na02f80 g781053 ( .a(cos_out_23), .b(FE_OFN1_n_43918), .o(n_298) );
na02f80 g742390 ( .a(n_37721), .b(n_37697), .o(n_37746) );
in01f80 FE_OCP_DRV_C1607_n_31473 ( .a(n_31473), .o(FE_OCP_DRV_N1607_n_31473) );
na02f80 g778134 ( .a(n_3494), .b(FE_OCP_RBN2297_n_2438), .o(n_2866) );
in01f80 g770662 ( .a(n_10225), .o(n_11380) );
ao12f80 g767368 ( .a(n_13417), .b(n_13397), .c(n_13383), .o(n_13468) );
na02f80 g780446 ( .a(n_855), .b(n_7), .o(n_784) );
in01f80 FE_OCP_RBC3038_n_47269 ( .a(n_47269), .o(FE_OCP_RBN3038_n_47269) );
in01f80 g768928 ( .a(n_11776), .o(n_11847) );
in01f80 newInst_2467 ( .a(newNet_2466), .o(newNet_2467) );
no02f80 g746711 ( .a(n_33270), .b(n_33202), .o(n_33290) );
na02f80 g758989 ( .a(n_21288), .b(n_21287), .o(n_21326) );
no02f80 g766294 ( .a(n_14281), .b(n_14330), .o(n_14441) );
in01f80 g781247 ( .a(n_133), .o(n_134) );
na02f80 g744255 ( .a(FE_OCPN1510_n_44174), .b(n_36091), .o(n_36242) );
no02f80 g740224 ( .a(n_40031), .b(FE_OCP_RBN3022_n_39942), .o(n_40104) );
no02f80 g740418 ( .a(FE_OCP_RBN3027_n_39942), .b(FE_OCP_RBN2871_n_39542), .o(n_40128) );
in01f80 g741488 ( .a(n_38746), .o(n_38750) );
no02f80 g756007 ( .a(n_25188), .b(n_25285), .o(n_25340) );
no02f80 FE_RC_2286_0 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_), .b(FE_RN_855_0), .o(FE_RN_856_0) );
na02f80 g742441 ( .a(n_37693), .b(FE_OCP_RBN3398_n_37624), .o(n_37696) );
na02f80 g775613 ( .a(n_5552), .b(n_5517), .o(n_5518) );
no02f80 g775397 ( .a(n_5796), .b(n_5654), .o(n_5888) );
na02f80 g758029 ( .a(n_22229), .b(n_22267), .o(n_22381) );
in01f80 g740809 ( .a(n_39352), .o(n_39353) );
no02f80 g768521 ( .a(n_12339), .b(n_12345), .o(n_12419) );
na02f80 g757994 ( .a(n_22923), .b(n_22847), .o(n_22978) );
in01f80 newInst_615 ( .a(newNet_197), .o(newNet_615) );
no02f80 g742078 ( .a(FE_OCP_RBN3441_n_37945), .b(n_37548), .o(n_38333) );
ao12f80 g760638 ( .a(n_20257), .b(n_20277), .c(n_20256), .o(n_21246) );
na02f80 g774007 ( .a(n_6860), .b(n_4948), .o(n_6968) );
ao12f80 g772419 ( .a(n_8495), .b(n_8503), .c(n_8494), .o(n_9681) );
no02f80 g742799 ( .a(n_37331), .b(n_37330), .o(n_37332) );
in01f80 newInst_1941 ( .a(newNet_1940), .o(newNet_1941) );
no02f80 g750648 ( .a(n_29440), .b(FE_OCP_DRV_N3739_n_29439), .o(n_29466) );
na02f80 g769641 ( .a(n_11310), .b(n_11259), .o(n_11326) );
in01f80 g772289 ( .a(n_8732), .o(n_10409) );
oa12f80 g767920 ( .a(n_12708), .b(n_12707), .c(n_12706), .o(n_12763) );
na03f80 g767362 ( .a(n_13077), .b(n_13638), .c(n_13621), .o(n_13675) );
no02f80 g774787 ( .a(n_45479), .b(n_6263), .o(n_6321) );
na02f80 g776740 ( .a(n_3946), .b(n_3868), .o(n_4081) );
ao12f80 g756351 ( .a(n_23594), .b(n_23948), .c(n_23635), .o(n_24002) );
in01f80 g768542 ( .a(n_12299), .o(n_12300) );
oa12f80 g775560 ( .a(n_5394), .b(n_5590), .c(n_5288), .o(n_5622) );
in01f80 newInst_3676 ( .a(newNet_3675), .o(newNet_3676) );
na02f80 g741525 ( .a(n_38691), .b(n_38721), .o(n_38722) );
in01f80 g764775 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .o(n_17158) );
no02f80 g737664 ( .a(FE_OCPN887_n_42367), .b(n_41884), .o(n_42589) );
no02f80 g770651 ( .a(n_9946), .b(n_9936), .o(n_10106) );
in01f80 FE_OCP_RBC2617_n_44561 ( .a(FE_OCP_RBN3573_n_44563), .o(FE_OCP_RBN2617_n_44561) );
in01f80 g759780 ( .a(n_21627), .o(n_21628) );
in01f80 g751321 ( .a(n_29600), .o(n_29992) );
in01f80 g754715 ( .a(n_26547), .o(n_26608) );
in01f80 g775306 ( .a(n_5561), .o(n_5562) );
oa12f80 g761622 ( .a(n_18843), .b(n_19526), .c(n_18932), .o(n_19578) );
in01f80 FE_OFC759_n_45813 ( .a(FE_OFN757_n_45813), .o(FE_OFN759_n_45813) );
no02f80 g754228 ( .a(n_25898), .b(n_23254), .o(n_25922) );
ao12f80 g778301 ( .a(n_2600), .b(n_2599), .c(FE_OCP_RBN2274_n_2457), .o(n_4231) );
in01f80 FE_OCP_RBC2568_n_8904 ( .a(n_8904), .o(FE_OCP_RBN2568_n_8904) );
in01f80 FE_OCP_RBC2118_n_45224 ( .a(FE_OCP_RBN2116_n_45224), .o(FE_OCP_RBN2118_n_45224) );
in01f80 g766389 ( .a(n_14199), .o(n_14187) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_10_ ( .ck(newNet_3175), .d(n_40419), .o(delay_add_ln22_unr27_stage10_stallmux_q_10_) );
oa12f80 g784439 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .b(n_37138), .c(n_46197), .o(n_46251) );
na02f80 g742506 ( .a(n_37580), .b(n_37560), .o(n_37667) );
ao12f80 g770601 ( .a(n_10429), .b(n_10428), .c(n_8687), .o(n_10637) );
in01f80 g758441 ( .a(FE_OCPN1440_n_23339), .o(n_23353) );
oa22f80 g744623 ( .a(n_36575), .b(n_35965), .c(n_36576), .d(n_35964), .o(n_36640) );
na02f80 g736878 ( .a(n_43355), .b(n_43501), .o(n_43603) );
na02f80 g736759 ( .a(n_43110), .b(n_43183), .o(n_43220) );
no02f80 g751917 ( .a(n_29170), .b(n_29200), .o(n_29336) );
na02f80 g751013 ( .a(n_29855), .b(n_29854), .o(n_29947) );
ao12f80 g772557 ( .a(n_8234), .b(n_8276), .c(n_8208), .o(n_8403) );
in01f80 newInst_3132 ( .a(newNet_43), .o(newNet_3132) );
oa12f80 g778298 ( .a(n_2901), .b(n_2910), .c(delay_add_ln22_unr2_stage2_stallmux_q_31_), .o(n_2973) );
oa22f80 g784552 ( .a(FE_OFN800_n_46285), .b(n_10885), .c(FE_OCP_RBN3709_n_46337), .d(n_10799), .o(n_46373) );
in01f80 g739894 ( .a(n_40343), .o(n_40344) );
no02f80 g761534 ( .a(FE_OCP_RBN1837_FE_RN_1542_0), .b(n_18320), .o(n_18801) );
no02f80 g774336 ( .a(n_6504), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6550) );
in01f80 g763801 ( .a(n_17465), .o(n_17466) );
na02f80 g743851 ( .a(n_36013), .b(n_35913), .o(n_36071) );
no02f80 g756715 ( .a(n_23432), .b(n_23329), .o(n_23507) );
in01f80 g774048 ( .a(n_6889), .o(n_6845) );
na02f80 g772668 ( .a(n_8275), .b(n_8251), .o(n_8252) );
na02f80 FE_RC_2107_0 ( .a(FE_RN_728_0), .b(FE_OCP_RBN1215_n_20595), .o(n_20694) );
no02f80 g748813 ( .a(n_32410), .b(n_32499), .o(n_32765) );
ao12f80 g740983 ( .a(n_39026), .b(FE_OCP_RBN2638_n_38806), .c(n_39055), .o(n_39161) );
ao12f80 g776814 ( .a(n_3880), .b(n_3987), .c(n_3943), .o(n_4075) );
in01f80 FE_RC_1122_0 ( .a(n_23229), .o(FE_RN_339_0) );
no02f80 g752434 ( .a(n_28401), .b(n_28379), .o(n_28380) );
no02f80 g739365 ( .a(n_40727), .b(n_40802), .o(n_41057) );
na02f80 g763524 ( .a(FE_OCP_RBN3079_n_16977), .b(n_16050), .o(n_17115) );
na02f80 g769923 ( .a(n_10974), .b(n_44463), .o(n_11026) );
no02f80 FE_RC_2174_0 ( .a(FE_RN_774_0), .b(n_26378), .o(n_26445) );
in01f80 g746333 ( .a(n_34160), .o(n_33632) );
no02f80 g754700 ( .a(n_26160), .b(n_26192), .o(n_26193) );
oa22f80 g780120 ( .a(n_1194), .b(n_1203), .c(n_1185), .d(FE_OFN761_n_45813), .o(n_1211) );
ao12f80 g749578 ( .a(n_31186), .b(n_31672), .c(n_31257), .o(n_31709) );
in01f80 g760419 ( .a(n_20098), .o(n_20099) );
in01f80 g764406 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n_16618) );
ao12f80 g768818 ( .a(n_11966), .b(n_12005), .c(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n_12125) );
na02f80 g776453 ( .a(n_4542), .b(FE_OCP_RBN2538_n_3645), .o(n_4591) );
no02f80 g755070 ( .a(n_25351), .b(n_25377), .o(n_25477) );
in01f80 g780270 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_8_), .o(n_1047) );
no02f80 g755347 ( .a(n_24910), .b(n_24620), .o(n_24937) );
na02f80 g763772 ( .a(n_17160), .b(n_17015), .o(n_17367) );
in01f80 g768287 ( .a(n_12656), .o(n_12657) );
in01f80 FE_OCPC1472_n_13434 ( .a(FE_OCPN1471_n_13434), .o(FE_OCPN1472_n_13434) );
na02f80 g748113 ( .a(n_31562), .b(n_31548), .o(n_31746) );
in01f80 newInst_1460 ( .a(newNet_1459), .o(newNet_1460) );
in01f80 g760451 ( .a(n_20064), .o(n_20065) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_17_ ( .ck(newNet_2481), .d(n_32263), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_) );
oa12f80 g738220 ( .a(n_41934), .b(n_41946), .c(n_41933), .o(n_41960) );
in01f80 FE_OFC834_n_2285 ( .a(n_2285), .o(FE_OFN834_n_2285) );
oa12f80 g739854 ( .a(n_40194), .b(n_40402), .c(n_40273), .o(n_40429) );
no02f80 g765138 ( .a(n_15083), .b(n_14210), .o(n_15125) );
na02f80 g766828 ( .a(n_13908), .b(n_14452), .o(n_14562) );
no02f80 g774294 ( .a(FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .o(n_6600) );
no02f80 g753203 ( .a(n_27087), .b(n_27117), .o(n_27118) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_3_ ( .ck(newNet_1803), .d(n_16410), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_) );
in01f80 g765227 ( .a(n_15637), .o(n_15638) );
oa12f80 g751283 ( .a(n_29694), .b(n_29693), .c(n_29692), .o(n_30086) );
ao12f80 g750268 ( .a(n_30253), .b(n_30812), .c(n_30125), .o(n_30925) );
in01f80 newInst_2417 ( .a(newNet_2416), .o(newNet_2417) );
na02f80 g775323 ( .a(n_5826), .b(n_5880), .o(n_5971) );
in01f80 g757052 ( .a(n_24007), .o(n_23899) );
no02f80 g749571 ( .a(n_45631), .b(n_30356), .o(n_30357) );
na02f80 g743421 ( .a(n_36647), .b(n_36750), .o(n_36688) );
no02f80 g757865 ( .a(n_22420), .b(n_22473), .o(n_22474) );
na02f80 g757853 ( .a(n_22421), .b(n_22064), .o(n_22444) );
no02f80 FE_RC_2409_0 ( .a(FE_RN_949_0), .b(n_6641), .o(n_7031) );
in01f80 newInst_3694 ( .a(newNet_3693), .o(newNet_3694) );
in01f80 newInst_2667 ( .a(newNet_2666), .o(newNet_2667) );
in01f80 g771799 ( .a(n_8872), .o(n_8906) );
na02f80 g765512 ( .a(FE_OFN765_n_15670), .b(n_15663), .o(n_15749) );
no02f80 g776808 ( .a(n_3738), .b(n_2989), .o(n_3834) );
oa22f80 g771312 ( .a(n_9780), .b(n_9435), .c(n_9654), .d(n_9436), .o(n_9832) );
na02f80 g737610 ( .a(n_42463), .b(n_42441), .o(n_42442) );
no02f80 g756936 ( .a(n_23806), .b(n_23700), .o(n_23990) );
no02f80 g774033 ( .a(n_6775), .b(n_6595), .o(n_6791) );
no02f80 g773075 ( .a(n_7988), .b(n_7909), .o(n_7989) );
oa12f80 g751215 ( .a(FE_OCPN962_n_28506), .b(n_28790), .c(n_28471), .o(n_28852) );
na02f80 g741241 ( .a(FE_OCP_RBN2638_n_38806), .b(n_38485), .o(n_38879) );
na02f80 g749484 ( .a(n_30471), .b(n_30239), .o(n_30469) );
na02f80 g778649 ( .a(n_2387), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_), .o(n_2422) );
in01f80 FE_OCPC976_n_31594 ( .a(n_31594), .o(FE_OCPN976_n_31594) );
in01f80 g741232 ( .a(n_39201), .o(n_39202) );
in01f80 FE_OCP_RBC2308_n_29298 ( .a(n_29298), .o(FE_OCP_RBN2308_n_29298) );
na02f80 g746249 ( .a(n_33644), .b(n_33620), .o(n_33660) );
no02f80 g742314 ( .a(n_37832), .b(n_37811), .o(n_37864) );
in01f80 newInst_3324 ( .a(newNet_3323), .o(newNet_3324) );
no02f80 g778126 ( .a(n_2888), .b(n_3378), .o(n_2928) );
in01f80 g759554 ( .a(n_20930), .o(n_20931) );
na02f80 g750732 ( .a(n_46960), .b(FE_OFN788_n_25834), .o(n_29239) );
no02f80 g750879 ( .a(n_29020), .b(n_28605), .o(n_29063) );
ao22s80 FE_RC_3878_0 ( .a(n_24620), .b(n_24798), .c(n_22280), .d(n_24799), .o(n_24891) );
no02f80 g772849 ( .a(n_7976), .b(n_7783), .o(n_8041) );
na02f80 g763679 ( .a(n_17306), .b(n_17055), .o(n_17370) );
no02f80 g774358 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .o(n_6868) );
na02f80 g744072 ( .a(n_44222), .b(FE_OCP_RBN2563_n_34905), .o(n_35948) );
no02f80 g768661 ( .a(n_12104), .b(n_11825), .o(n_12242) );
na02f80 FE_RC_2894_0 ( .a(n_39816), .b(FE_RN_1253_0), .o(FE_RN_1254_0) );
in01f80 g741314 ( .a(n_38901), .o(n_38990) );
in01f80 g765065 ( .a(n_15321), .o(n_15284) );
no02f80 g770758 ( .a(n_10175), .b(n_10257), .o(n_10461) );
no02f80 g765319 ( .a(FE_OCP_RBN3507_n_13860), .b(FE_OCP_RBN2681_n_15048), .o(n_15269) );
in01f80 newInst_3475 ( .a(newNet_1698), .o(newNet_3475) );
in01f80 g741775 ( .a(n_38512), .o(n_38513) );
no02f80 g759044 ( .a(n_21084), .b(n_45070), .o(n_21202) );
in01f80 FE_RC_3105_0 ( .a(n_31770), .o(FE_RN_1373_0) );
in01f80 newInst_3344 ( .a(newNet_3343), .o(newNet_3344) );
in01f80 FE_OCP_RBC3268_n_45224 ( .a(FE_OCP_RBN3269_n_45224), .o(FE_OCP_RBN3268_n_45224) );
no02f80 g741664 ( .a(n_38524), .b(n_38218), .o(n_38570) );
in01f80 g746965 ( .a(n_33136), .o(n_33137) );
in01f80 g775517 ( .a(n_5741), .o(n_5742) );
no02f80 g778556 ( .a(n_2456), .b(n_2350), .o(n_2501) );
na02f80 g754937 ( .a(n_25270), .b(n_24633), .o(n_25506) );
in01f80 g774088 ( .a(n_6824), .o(n_6825) );
oa12f80 g765118 ( .a(n_15417), .b(n_15416), .c(n_15415), .o(n_15489) );
na02f80 FE_RC_3554_0 ( .a(FE_RN_1541_0), .b(n_18650), .o(FE_RN_1542_0) );
no02f80 g743956 ( .a(n_35751), .b(n_35754), .o(n_35787) );
no02f80 g774317 ( .a(FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .o(n_6708) );
in01f80 newInst_838 ( .a(newNet_837), .o(newNet_838) );
na02f80 g746236 ( .a(n_33706), .b(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33752) );
in01f80 FE_RC_42_0 ( .a(n_2538), .o(FE_RN_10_0) );
in01f80 FE_OCP_RBC3366_n_44722 ( .a(FE_OCP_RBN3365_n_44722), .o(FE_OCP_RBN3366_n_44722) );
oa22f80 g751526 ( .a(FE_OCP_RBN3408_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_), .c(FE_OCP_RBN3406_n_28597), .d(n_27803), .o(n_28845) );
na02f80 g776297 ( .a(n_4604), .b(n_4464), .o(n_4638) );
in01f80 FE_OCP_RBC1727_FE_RN_1583_0 ( .a(FE_RN_1583_0), .o(FE_OCP_RBN1727_FE_RN_1583_0) );
in01f80 newInst_608 ( .a(newNet_607), .o(newNet_608) );
in01f80 g750340 ( .a(n_30756), .o(n_30783) );
na02f80 g749842 ( .a(FE_OCP_RBN3009_n_31117), .b(n_31145), .o(n_31460) );
in01f80 FE_OCP_RBC2529_n_9044 ( .a(n_9044), .o(FE_OCP_RBN2529_n_9044) );
oa22f80 g747770 ( .a(n_33372), .b(n_33114), .c(n_33571), .d(n_33552), .o(n_33999) );
in01f80 g748118 ( .a(n_32021), .o(n_32022) );
ao12f80 g781010 ( .a(n_268), .b(n_267), .c(n_266), .o(n_465) );
ao12f80 g746412 ( .a(n_33483), .b(n_33484), .c(n_33482), .o(n_33534) );
in01f80 FE_OCP_RBC2890_n_10568 ( .a(n_10568), .o(FE_OCP_RBN2890_n_10568) );
na02f80 g740183 ( .a(FE_OCP_RBN3719_n_39913), .b(n_40007), .o(n_40178) );
oa12f80 g741802 ( .a(n_38442), .b(n_38441), .c(n_38440), .o(n_38562) );
na02f80 g737779 ( .a(n_42580), .b(n_42515), .o(n_42625) );
in01f80 newInst_3566 ( .a(newNet_3565), .o(newNet_3566) );
in01f80 newInst_3377 ( .a(newNet_3376), .o(newNet_3377) );
no02f80 g750426 ( .a(n_29545), .b(n_29630), .o(n_29580) );
in01f80 g753715 ( .a(n_27198), .o(n_27199) );
ao22s80 FE_RC_3427_0 ( .a(FE_RN_1643_0), .b(n_25928), .c(n_23317), .d(n_26113), .o(n_26039) );
ao12f80 g747605 ( .a(n_34072), .b(n_34071), .c(n_34070), .o(n_35655) );
no02f80 g747741 ( .a(n_33317), .b(n_33316), .o(n_33318) );
in01f80 g751456 ( .a(n_28572), .o(n_28573) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_0_ ( .ck(newNet_987), .d(n_22449), .o(delay_xor_ln21_unr15_stage6_stallmux_q_0_) );
ao12f80 g742407 ( .a(n_37740), .b(n_37762), .c(n_37739), .o(n_37797) );
na02f80 g755319 ( .a(n_25577), .b(n_25576), .o(n_25578) );
in01f80 g774129 ( .a(n_7286), .o(n_6730) );
in01f80 g772711 ( .a(n_8239), .o(n_8240) );
na02f80 g760981 ( .a(n_19323), .b(n_19253), .o(n_19380) );
oa22f80 FE_RC_389_0 ( .a(n_1004), .b(n_44652), .c(n_967), .d(n_44637), .o(n_1328) );
in01f80 newInst_1928 ( .a(newNet_263), .o(newNet_1928) );
na02f80 g746432 ( .a(n_33468), .b(n_33467), .o(n_33469) );
na02f80 g764259 ( .a(n_16723), .b(n_16384), .o(n_16772) );
oa12f80 g778928 ( .a(n_1663), .b(n_2148), .c(n_1783), .o(n_2184) );
in01f80 FE_OCPC1395_n_7881 ( .a(n_7881), .o(FE_OCPN1395_n_7881) );
in01f80 newInst_3464 ( .a(newNet_3463), .o(newNet_3464) );
ao22s80 g770016 ( .a(n_10808), .b(n_10416), .c(n_10798), .d(n_10415), .o(n_10944) );
in01f80 newInst_2558 ( .a(newNet_2550), .o(newNet_2558) );
no02f80 g770236 ( .a(n_10629), .b(FE_OFN756_n_44461), .o(n_10669) );
in01f80 g775186 ( .a(n_5766), .o(n_5787) );
in01f80 g764111 ( .a(n_16603), .o(n_16604) );
na02f80 g737702 ( .a(n_42285), .b(n_42312), .o(n_42402) );
in01f80 g768057 ( .a(n_12963), .o(n_13034) );
na03f80 g743249 ( .a(n_37878), .b(n_38019), .c(n_38021), .o(n_38076) );
in01f80 g756407 ( .a(n_23792), .o(n_23793) );
in01f80 newInst_2571 ( .a(newNet_2094), .o(newNet_2571) );
in01f80 newInst_1112 ( .a(newNet_458), .o(newNet_1112) );
in01f80 g772019 ( .a(n_9733), .o(n_9734) );
no02f80 g748108 ( .a(n_32804), .b(n_32803), .o(n_32805) );
in01f80 g774939 ( .a(n_6267), .o(n_6245) );
na02f80 g770507 ( .a(n_10324), .b(n_47263), .o(n_10365) );
ao12f80 g764744 ( .a(n_15495), .b(n_45135), .c(n_15493), .o(n_15661) );
in01f80 FE_OCP_RBC1704_n_22740 ( .a(n_22740), .o(FE_OCP_RBN1704_n_22740) );
in01f80 g760787 ( .a(n_19594), .o(n_19595) );
in01f80 newInst_2848 ( .a(newNet_2097), .o(newNet_2848) );
no02f80 g773052 ( .a(n_7645), .b(n_7703), .o(n_7752) );
no02f80 g740523 ( .a(n_39665), .b(n_39677), .o(n_39702) );
na02f80 g779182 ( .a(n_1938), .b(n_1011), .o(n_2007) );
oa22f80 FE_RC_644_0 ( .a(n_29426), .b(n_28845), .c(n_29425), .d(n_28846), .o(n_29553) );
na02f80 g756601 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_22_), .o(n_23761) );
ao12f80 g773033 ( .a(n_7235), .b(n_7636), .c(n_7252), .o(n_7662) );
in01f80 FE_OCP_RBC3659_n_15314 ( .a(FE_OCP_RBN3658_n_15314), .o(FE_OCP_RBN3659_n_15314) );
no02f80 g742245 ( .a(n_37848), .b(n_37847), .o(n_37905) );
oa12f80 g745469 ( .a(n_34154), .b(n_34167), .c(n_34153), .o(n_35594) );
no02f80 g756527 ( .a(FE_OCP_RBN2276_n_24077), .b(n_23809), .o(n_24109) );
na02f80 g752330 ( .a(n_27868), .b(n_27802), .o(n_27831) );
na02f80 g746552 ( .a(n_34757), .b(n_34775), .o(n_34803) );
oa22f80 FE_RC_1439_0 ( .a(n_32287), .b(n_32311), .c(n_28336), .d(n_32286), .o(n_32352) );
in01f80 g738161 ( .a(n_42029), .o(n_42016) );
no02f80 g751393 ( .a(n_29838), .b(n_29359), .o(n_29360) );
ao22s80 FE_RC_3787_0 ( .a(n_31046), .b(n_30799), .c(n_31045), .d(n_31122), .o(n_31148) );
in01f80 g753785 ( .a(n_26465), .o(n_26466) );
in01f80 g762064 ( .a(n_18669), .o(n_18670) );
in01f80 g781166 ( .a(FE_OCPN1386_n_470), .o(n_193) );
in01f80 newInst_2245 ( .a(newNet_2244), .o(newNet_2245) );
na02f80 g777022 ( .a(n_3770), .b(n_3802), .o(n_3973) );
na02f80 g739716 ( .a(n_40542), .b(n_40438), .o(n_40563) );
no02f80 g777984 ( .a(n_3079), .b(n_3037), .o(n_3142) );
in01f80 g765173 ( .a(n_15160), .o(n_15161) );
na02f80 g744158 ( .a(n_35551), .b(n_35556), .o(n_35552) );
in01f80 g757314 ( .a(n_23191), .o(n_23042) );
in01f80 FE_OCP_RBC3661_n_15429 ( .a(n_15429), .o(FE_OCP_RBN3661_n_15429) );
in01f80 g736678 ( .a(n_43095), .o(n_43096) );
oa12f80 g737428 ( .a(n_42723), .b(n_42722), .c(n_42721), .o(n_42772) );
in01f80 g738484 ( .a(n_41391), .o(n_41769) );
no02f80 g757901 ( .a(n_22885), .b(n_24105), .o(n_22886) );
no02f80 g774090 ( .a(n_7172), .b(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .o(n_7195) );
in01f80 g768655 ( .a(n_12228), .o(n_12293) );
in01f80 FE_OFC764_n_15670 ( .a(FE_OFN762_n_15670), .o(FE_OFN764_n_15670) );
na02f80 g756810 ( .a(n_23452), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .o(n_23512) );
in01f80 newInst_1891 ( .a(newNet_1890), .o(newNet_1891) );
na02f80 g770946 ( .a(n_9806), .b(n_9820), .o(n_9893) );
ao12f80 g778073 ( .a(n_2375), .b(n_2924), .c(n_2331), .o(n_3008) );
in01f80 fopt783583 ( .a(n_8405), .o(n_45213) );
na02f80 g755440 ( .a(n_24874), .b(FE_OCPN1512_n_22280), .o(n_24828) );
in01f80 newInst_715 ( .a(newNet_576), .o(newNet_715) );
in01f80 g740794 ( .a(n_39355), .o(n_39448) );
na02f80 g742470 ( .a(n_37626), .b(n_37598), .o(n_37665) );
in01f80 FE_RC_2248_0 ( .a(n_37279), .o(FE_RN_827_0) );
na02f80 g770029 ( .a(n_10958), .b(n_10957), .o(n_10989) );
na02f80 g742906 ( .a(n_37006), .b(n_36465), .o(n_37007) );
oa12f80 g754503 ( .a(n_26934), .b(n_26933), .c(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_26997) );
oa12f80 g759815 ( .a(n_21668), .b(n_21691), .c(n_21595), .o(n_21821) );
oa12f80 g750387 ( .a(n_30591), .b(n_30590), .c(n_30589), .o(n_31251) );
na02f80 g739574 ( .a(n_40653), .b(n_40654), .o(n_40646) );
in01f80 newInst_1702 ( .a(newNet_1701), .o(newNet_1702) );
no02f80 g741986 ( .a(n_38057), .b(n_37974), .o(n_38013) );
in01f80 fopt783659 ( .a(n_10742), .o(n_45304) );
in01f80 g770437 ( .a(n_10631), .o(n_10680) );
na02f80 g748872 ( .a(n_32375), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32555) );
no02f80 g776213 ( .a(n_4913), .b(n_4866), .o(n_5015) );
in01f80 newInst_1101 ( .a(newNet_1100), .o(newNet_1101) );
in01f80 g750460 ( .a(n_29620), .o(n_29621) );
in01f80 g744319 ( .a(n_35565), .o(n_35566) );
na02f80 g766962 ( .a(n_13519), .b(n_12954), .o(n_13633) );
in01f80 g775917 ( .a(n_5013), .o(n_5014) );
no02f80 g740432 ( .a(FE_OCP_RBN3031_n_39942), .b(n_40202), .o(n_40238) );
na02f80 g750092 ( .a(n_29831), .b(FE_OCP_DRV_N1576_n_28829), .o(n_29864) );
ao12f80 g777754 ( .a(n_3307), .b(n_3306), .c(n_3305), .o(n_4797) );
in01f80 g744265 ( .a(n_35619), .o(n_35588) );
in01f80 fopt783289 ( .a(n_44869), .o(n_44867) );
in01f80 g749292 ( .a(n_30657), .o(n_30658) );
oa12f80 g755461 ( .a(n_24713), .b(n_24779), .c(n_24636), .o(n_24834) );
na02f80 g759359 ( .a(n_20997), .b(n_20666), .o(n_21120) );
in01f80 FE_OCP_RBC3213_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3213_n_44365) );
ao12f80 g741843 ( .a(n_38063), .b(n_38363), .c(n_37940), .o(n_38397) );
ao12f80 g739193 ( .a(n_45153), .b(n_40831), .c(n_40575), .o(n_40832) );
ao12f80 g780231 ( .a(n_1081), .b(n_1080), .c(n_1079), .o(n_1138) );
na02f80 g754016 ( .a(n_26141), .b(n_26124), .o(n_26210) );
na02f80 g755603 ( .a(n_24597), .b(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24719) );
oa22f80 FE_RC_3339_0 ( .a(n_14755), .b(n_14803), .c(n_14773), .d(n_14802), .o(n_14911) );
no02f80 FE_RC_2641_0 ( .a(n_2759), .b(n_3421), .o(FE_RN_1101_0) );
in01f80 g769425 ( .a(n_11455), .o(n_11440) );
no02f80 g746899 ( .a(FE_OCP_RBN3384_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n_33323) );
no02f80 g747663 ( .a(n_32300), .b(n_31869), .o(n_32301) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_5_ ( .ck(newNet_1901), .d(n_36845), .o(delay_sub_ln22_unr24_stage9_stallmux_q_5_) );
no02f80 g739422 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .o(n_40811) );
in01f80 g775196 ( .a(n_5927), .o(n_5941) );
na02f80 g738535 ( .a(n_41390), .b(n_41389), .o(n_41408) );
in01f80 g748718 ( .a(n_31419), .o(n_31420) );
no02f80 g738274 ( .a(n_41823), .b(n_41733), .o(n_41919) );
na02f80 g740209 ( .a(n_39895), .b(n_39803), .o(n_39975) );
no02f80 g744850 ( .a(n_35134), .b(n_35096), .o(n_35135) );
oa22f80 g740352 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39470), .c(FE_OCP_RBN3028_n_39942), .d(n_39894), .o(n_40386) );
in01f80 g772478 ( .a(n_10137), .o(n_8539) );
na02f80 FE_RC_2701_0 ( .a(n_8302), .b(n_8231), .o(FE_RN_1134_0) );
in01f80 g764990 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_5_), .o(n_17589) );
no02f80 g740090 ( .a(n_40107), .b(n_40034), .o(n_40136) );
no02f80 g779415 ( .a(n_1494), .b(n_1427), .o(n_1509) );
oa22f80 g741095 ( .a(FE_OCP_RBN2687_n_38870), .b(n_38484), .c(FE_OCPN957_n_39096), .d(n_38508), .o(n_39364) );
no02f80 g781324 ( .a(n_7), .b(beta_26), .o(n_119) );
ao12f80 g774122 ( .a(n_7143), .b(n_6872), .c(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .o(n_7322) );
na02f80 g767826 ( .a(n_12799), .b(n_12747), .o(n_13221) );
in01f80 newInst_630 ( .a(newNet_629), .o(newNet_630) );
no02f80 g775430 ( .a(n_5576), .b(n_5544), .o(n_5700) );
na02f80 g756195 ( .a(n_24816), .b(n_24815), .o(n_24817) );
na02f80 g763745 ( .a(n_16661), .b(n_16670), .o(n_16710) );
na02f80 g776983 ( .a(n_3943), .b(n_3879), .o(n_3966) );
na02f80 g771622 ( .a(n_9392), .b(FE_OFN361_n_9391), .o(n_9393) );
in01f80 g738204 ( .a(n_41989), .o(n_41990) );
no02f80 g777188 ( .a(n_5006), .b(n_4863), .o(n_5949) );
na02f80 FE_RC_2998_0 ( .a(FE_RN_1310_0), .b(FE_RN_1311_0), .o(FE_RN_1312_0) );
na02f80 g767647 ( .a(FE_OCP_RBN2201_n_12808), .b(n_12849), .o(n_12866) );
no02f80 g771364 ( .a(n_9089), .b(n_9112), .o(n_9255) );
in01f80 FE_RC_646_0 ( .a(n_37471), .o(FE_RN_204_0) );
no02f80 g746506 ( .a(n_34527), .b(n_35542), .o(n_34528) );
na02f80 g760126 ( .a(n_20395), .b(n_47258), .o(n_20495) );
in01f80 newInst_1646 ( .a(newNet_1645), .o(newNet_1646) );
in01f80 newInst_1375 ( .a(newNet_1374), .o(newNet_1375) );
no02f80 g770553 ( .a(n_10354), .b(n_10338), .o(n_10372) );
oa22f80 FE_RC_3033_0 ( .a(n_11701), .b(n_11954), .c(n_11700), .d(n_11982), .o(n_12158) );
in01f80 FE_RC_2792_0 ( .a(n_13017), .o(FE_RN_1193_0) );
no02f80 g749887 ( .a(n_30117), .b(FE_OCP_RBN3567_n_29857), .o(n_30175) );
na02f80 g760187 ( .a(n_20603), .b(n_20626), .o(n_20744) );
oa12f80 g766155 ( .a(n_14837), .b(n_14836), .c(n_14835), .o(n_15865) );
in01f80 FE_RC_850_0 ( .a(FE_RN_254_0), .o(n_29533) );
na02f80 g781076 ( .a(n_273), .b(n_270), .o(n_271) );
no02f80 g753199 ( .a(n_25957), .b(n_27103), .o(n_27119) );
ao22s80 FE_RC_1499_0 ( .a(FE_OCP_RBN3835_n_19241), .b(n_19781), .c(FE_OCP_RBN3834_n_19241), .d(FE_OCP_RBN3217_n_19781), .o(n_19891) );
no02f80 g779738 ( .a(n_1379), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .o(n_1456) );
na02f80 g777159 ( .a(n_5112), .b(n_5247), .o(n_5258) );
in01f80 newInst_408 ( .a(newNet_407), .o(newNet_408) );
no02f80 g752791 ( .a(n_28107), .b(n_28106), .o(n_28130) );
no02f80 FE_RC_4254_0 ( .a(FE_RN_1871_0), .b(n_21983), .o(FE_RN_1872_0) );
no02f80 g741143 ( .a(n_38853), .b(n_38892), .o(n_38893) );
in01f80 FE_RC_3775_0 ( .a(n_23919), .o(FE_RN_1657_0) );
no02f80 g740241 ( .a(n_40274), .b(n_40152), .o(n_40316) );
in01f80 FE_OCP_RBC3055_n_39913 ( .a(FE_OCP_RBN3053_n_39913), .o(FE_OCP_RBN3055_n_39913) );
in01f80 newInst_243 ( .a(newNet_114), .o(newNet_243) );
no02f80 g744896 ( .a(n_34999), .b(n_30546), .o(n_35030) );
na02f80 g764922 ( .a(n_15434), .b(n_15187), .o(n_15475) );
oa12f80 g758825 ( .a(n_21603), .b(n_21705), .c(n_21529), .o(n_21794) );
in01f80 newInst_902 ( .a(newNet_901), .o(newNet_902) );
in01f80 FE_OCP_RBC3591_n_14704 ( .a(n_14704), .o(FE_OCP_RBN3591_n_14704) );
na02f80 g737905 ( .a(n_42189), .b(n_42188), .o(n_42193) );
in01f80 newInst_3329 ( .a(newNet_184), .o(newNet_3329) );
oa12f80 g762958 ( .a(n_17982), .b(n_17981), .c(n_17980), .o(n_18531) );
in01f80 g755052 ( .a(n_25537), .o(n_25538) );
no02f80 g758724 ( .a(n_21897), .b(n_21896), .o(n_21910) );
in01f80 newInst_2938 ( .a(newNet_2937), .o(newNet_2938) );
in01f80 g777350 ( .a(n_3990), .o(n_3991) );
in01f80 g776442 ( .a(n_4689), .o(n_4644) );
in01f80 g739629 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_), .o(n_40582) );
in01f80 g770932 ( .a(n_9853), .o(n_9854) );
in01f80 newInst_3239 ( .a(newNet_2772), .o(newNet_3239) );
in01f80 g783839 ( .a(n_45528), .o(n_45529) );
no02f80 g776477 ( .a(n_4234), .b(n_3837), .o(n_4422) );
ao12f80 g736683 ( .a(n_43033), .b(n_43039), .c(n_43051), .o(n_43094) );
na02f80 g738955 ( .a(n_41238), .b(n_41237), .o(n_41239) );
na02f80 g747621 ( .a(n_32190), .b(n_31840), .o(n_32221) );
in01f80 g764442 ( .a(n_16273), .o(n_16368) );
in01f80 g768126 ( .a(n_12647), .o(n_12648) );
na02f80 g750728 ( .a(n_29169), .b(n_28768), .o(n_29219) );
oa12f80 g756284 ( .a(n_23663), .b(n_23949), .c(n_23609), .o(n_24056) );
no02f80 g774749 ( .a(n_6272), .b(FE_OCP_RBN2979_n_5656), .o(n_6294) );
in01f80 g743502 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_23_), .o(n_36992) );
in01f80 g756056 ( .a(n_24307), .o(n_24308) );
in01f80 g758032 ( .a(n_22377), .o(n_22378) );
na02f80 g740724 ( .a(n_39414), .b(n_38983), .o(n_39484) );
in01f80 g748372 ( .a(n_31823), .o(n_31824) );
in01f80 g755517 ( .a(n_26307), .o(n_26855) );
in01f80 g742204 ( .a(n_38296), .o(n_38297) );
na02f80 g776771 ( .a(n_4026), .b(n_4000), .o(n_4095) );
in01f80 g760822 ( .a(n_19535), .o(n_19536) );
in01f80 g779751 ( .a(n_1508), .o(n_1516) );
oa22f80 g757701 ( .a(n_22540), .b(n_22801), .c(n_22514), .d(n_22580), .o(n_22581) );
in01f80 g780985 ( .a(n_377), .o(n_403) );
no02f80 g766543 ( .a(n_14059), .b(FE_OCP_RBN2245_n_13017), .o(n_14121) );
in01f80 g742152 ( .a(n_38153), .o(n_38154) );
no02f80 g754113 ( .a(n_26818), .b(n_26578), .o(n_26911) );
in01f80 newInst_676 ( .a(newNet_675), .o(newNet_676) );
na02f80 g781019 ( .a(cos_out_4), .b(FE_OFN2_n_43918), .o(n_345) );
no02f80 g754408 ( .a(n_25754), .b(n_25509), .o(n_25807) );
oa12f80 g736599 ( .a(n_343), .b(n_43236), .c(FE_OFN2_n_43918), .o(n_43381) );
no02f80 g744832 ( .a(n_34982), .b(n_30588), .o(n_35015) );
oa12f80 g736265 ( .a(n_331), .b(n_43902), .c(FE_OFN4_n_43918), .o(n_43913) );
in01f80 g749179 ( .a(n_32205), .o(n_32203) );
ao12f80 g752726 ( .a(n_27787), .b(n_27909), .c(n_27882), .o(n_27997) );
oa12f80 g743714 ( .a(n_37359), .b(n_37405), .c(n_46233), .o(n_37540) );
no02f80 g742429 ( .a(n_37650), .b(n_37630), .o(n_37707) );
ms00f80 sin_out_reg_29_ ( .ck(newNet_36), .d(n_43920), .o(sin_out_29) );
oa12f80 g749085 ( .a(n_30751), .b(n_30750), .c(n_27014), .o(n_30834) );
in01f80 g740068 ( .a(n_40113), .o(n_40141) );
na02f80 g772236 ( .a(n_8608), .b(n_8104), .o(n_8633) );
na02f80 g773027 ( .a(n_8047), .b(n_8110), .o(n_8166) );
no02f80 g767494 ( .a(n_13393), .b(n_12788), .o(n_13444) );
no02f80 g777606 ( .a(n_3480), .b(n_3451), .o(n_4528) );
na02f80 g744545 ( .a(n_35334), .b(n_35234), .o(n_35369) );
oa12f80 g780153 ( .a(n_1149), .b(n_1170), .c(n_1148), .o(n_1190) );
na02f80 g780751 ( .a(n_584), .b(n_578), .o(n_579) );
in01f80 FE_OCPC1486_n_27315 ( .a(FE_OCPN1485_n_27315), .o(FE_OCPN1486_n_27315) );
ao12f80 g759957 ( .a(n_20090), .b(n_20195), .c(n_20144), .o(n_20251) );
na02f80 g745800 ( .a(n_44100), .b(n_33342), .o(n_34117) );
in01f80 FE_OCPC1450_n_20443 ( .a(FE_OCPN1449_n_20443), .o(FE_OCPN1450_n_20443) );
na02f80 g748443 ( .a(n_31699), .b(n_31756), .o(n_31784) );
in01f80 FE_RC_835_0 ( .a(n_8309), .o(FE_RN_249_0) );
oa12f80 g780999 ( .a(n_280), .b(n_279), .c(n_278), .o(n_493) );
in01f80 g749304 ( .a(n_30706), .o(n_30707) );
no02f80 g761318 ( .a(n_19827), .b(n_20178), .o(n_19934) );
in01f80 FE_OCP_RBC2127_n_6745 ( .a(n_6745), .o(FE_OCP_RBN2127_n_6745) );
ao22s80 g773892 ( .a(n_7007), .b(n_6856), .c(n_6996), .d(n_6855), .o(n_7071) );
no02f80 g750509 ( .a(n_30480), .b(n_30479), .o(n_30481) );
in01f80 g738453 ( .a(n_41853), .o(n_41854) );
in01f80 g756650 ( .a(n_23581), .o(n_23574) );
no02f80 FE_RC_2588_0 ( .a(n_12105), .b(n_12106), .o(FE_RN_1070_0) );
na02f80 g765384 ( .a(FE_OCP_RBN3622_n_15135), .b(n_14277), .o(n_15578) );
na02f80 g741589 ( .a(n_38639), .b(n_38636), .o(n_38664) );
in01f80 g781281 ( .a(n_123), .o(n_124) );
in01f80 g751576 ( .a(n_28489), .o(n_28490) );
na02f80 g759449 ( .a(n_21885), .b(n_21884), .o(n_21886) );
in01f80 newInst_2174 ( .a(newNet_2173), .o(newNet_2174) );
in01f80 newInst_266 ( .a(newNet_265), .o(newNet_266) );
in01f80 g763017 ( .a(n_17737), .o(n_17738) );
na02f80 g741036 ( .a(n_38864), .b(n_38836), .o(n_38895) );
no02f80 g759112 ( .a(n_21462), .b(n_21463), .o(n_21491) );
in01f80 g779842 ( .a(n_1377), .o(n_1416) );
na02f80 g770733 ( .a(n_10146), .b(FE_OFN755_n_44461), .o(n_10242) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_24_ ( .ck(newNet_1103), .d(n_11261), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_) );
no02f80 g760083 ( .a(n_21099), .b(n_21098), .o(n_21100) );
ao22s80 g739016 ( .a(n_41119), .b(n_41071), .c(n_41085), .d(n_41070), .o(n_41198) );
na02f80 g754358 ( .a(n_26941), .b(n_26940), .o(n_26942) );
in01f80 g751153 ( .a(n_30059), .o(n_30060) );
in01f80 g745290 ( .a(n_36172), .o(n_36173) );
oa12f80 g780083 ( .a(n_1196), .b(n_1198), .c(n_1195), .o(n_1207) );
na02f80 g777319 ( .a(n_5494), .b(n_4760), .o(n_5001) );
ao12f80 g738074 ( .a(n_42063), .b(n_42062), .c(n_42061), .o(n_42459) );
in01f80 g756480 ( .a(n_23923), .o(n_23924) );
na02f80 g775079 ( .a(n_5968), .b(n_5962), .o(n_5979) );
no02f80 g737301 ( .a(n_42909), .b(n_42891), .o(n_43250) );
in01f80 g739658 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_), .o(n_40558) );
in01f80 newInst_240 ( .a(newNet_239), .o(newNet_240) );
na02f80 g737001 ( .a(n_43230), .b(n_42994), .o(n_43501) );
in01f80 newInst_819 ( .a(newNet_818), .o(newNet_819) );
na02f80 g766694 ( .a(n_14217), .b(n_13977), .o(n_14308) );
oa12f80 g756347 ( .a(n_24031), .b(n_24453), .c(n_23981), .o(n_24514) );
no02f80 g742807 ( .a(n_37311), .b(n_37111), .o(n_37312) );
in01f80 newInst_2620 ( .a(newNet_2619), .o(newNet_2620) );
in01f80 FE_OCP_DRV_C1587_n_31012 ( .a(n_31012), .o(FE_OCP_DRV_N1587_n_31012) );
in01f80 FE_OCP_RBC2330_n_9003 ( .a(n_9003), .o(FE_OCP_RBN2330_n_9003) );
na02f80 g767938 ( .a(n_12627), .b(n_12448), .o(n_12654) );
na02f80 g769330 ( .a(n_11784), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11960) );
no02f80 g746216 ( .a(n_33711), .b(n_33689), .o(n_33690) );
na02f80 g756774 ( .a(n_23411), .b(n_23080), .o(n_23426) );
ao12f80 g752736 ( .a(n_27908), .b(n_27909), .c(n_27907), .o(n_27994) );
in01f80 newInst_1765 ( .a(newNet_1316), .o(newNet_1765) );
in01f80 g743888 ( .a(n_36011), .o(n_36041) );
oa12f80 g747976 ( .a(n_33071), .b(n_33070), .c(n_33069), .o(n_33573) );
ao12f80 g779464 ( .a(n_1759), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_14_), .o(n_1773) );
ao22s80 FE_RC_1252_0 ( .a(FE_OCP_RBN2410_n_13960), .b(n_13437), .c(FE_OCP_RBN2250_n_13017), .d(n_13960), .o(n_14127) );
na02f80 g755475 ( .a(n_24623), .b(FE_OCPN1474_n_24624), .o(n_24655) );
na02f80 g758318 ( .a(FE_OCPN992_n_22249), .b(n_21281), .o(n_22368) );
oa22f80 g778455 ( .a(n_2629), .b(n_2145), .c(n_2556), .d(n_2146), .o(n_2685) );
no02f80 g764986 ( .a(n_15499), .b(n_15535), .o(n_15679) );
in01f80 g771133 ( .a(n_9706), .o(n_9707) );
na02f80 g744112 ( .a(n_35547), .b(n_35590), .o(n_35591) );
no02f80 g752922 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .o(n_27992) );
na02f80 g767019 ( .a(n_13760), .b(n_13795), .o(n_13864) );
in01f80 FE_OCPC1463_n_29630 ( .a(n_29630), .o(FE_OCPN1463_n_29630) );
in01f80 g758842 ( .a(n_21509), .o(n_21554) );
no02f80 g766953 ( .a(n_14338), .b(n_14291), .o(n_14995) );
na02f80 g780407 ( .a(n_881), .b(n_806), .o(n_851) );
na02f80 g754269 ( .a(n_26944), .b(n_26943), .o(n_26945) );
no02f80 g775933 ( .a(n_5321), .b(n_3819), .o(n_5534) );
ao22s80 FE_RC_770_0 ( .a(n_9982), .b(n_10062), .c(n_9983), .d(n_10095), .o(n_10274) );
na02f80 g765502 ( .a(FE_OFN765_n_15670), .b(n_15669), .o(n_15783) );
in01f80 g739383 ( .a(n_40969), .o(n_40970) );
in01f80 newInst_3667 ( .a(newNet_3666), .o(newNet_3667) );
na02f80 g741788 ( .a(n_38344), .b(n_38113), .o(n_38369) );
in01f80 newInst_3089 ( .a(newNet_3088), .o(newNet_3089) );
no02f80 g766323 ( .a(n_14533), .b(FE_OCP_RBN2506_n_13896), .o(n_14534) );
na02f80 g754461 ( .a(n_26831), .b(n_26816), .o(n_26869) );
in01f80 g742642 ( .a(n_37446), .o(n_37447) );
in01f80 newInst_2991 ( .a(newNet_150), .o(newNet_2991) );
in01f80 newInst_2236 ( .a(newNet_2235), .o(newNet_2236) );
na02f80 g768757 ( .a(n_12065), .b(n_11758), .o(n_12108) );
na02f80 g751889 ( .a(n_29201), .b(n_29105), .o(n_29251) );
no02f80 g737507 ( .a(n_42475), .b(n_42474), .o(n_42541) );
in01f80 g766505 ( .a(n_14154), .o(n_14243) );
oa12f80 g751072 ( .a(n_30060), .b(n_30156), .c(n_29781), .o(n_30897) );
no02f80 g757360 ( .a(FE_OCPN1020_n_23078), .b(n_22912), .o(n_23000) );
oa12f80 g766769 ( .a(n_12836), .b(n_13601), .c(n_12766), .o(n_13694) );
na02f80 g758188 ( .a(n_22404), .b(n_22253), .o(n_22459) );
na02f80 g771865 ( .a(n_10077), .b(n_9952), .o(n_10942) );
no02f80 g744057 ( .a(n_44222), .b(n_35742), .o(n_35911) );
in01f80 g761798 ( .a(n_18676), .o(n_18677) );
na02f80 g775415 ( .a(n_5640), .b(n_4675), .o(n_5668) );
in01f80 newInst_130 ( .a(newNet_129), .o(newNet_130) );
no03m80 FE_RC_138_0 ( .a(beta_31), .b(n_65), .c(n_169), .o(n_170) );
na02f80 g745543 ( .a(n_35496), .b(n_34914), .o(n_35511) );
no02f80 g751367 ( .a(n_28745), .b(n_28626), .o(n_29017) );
in01f80 g773422 ( .a(n_7586), .o(n_7587) );
in01f80 FE_OCP_RBC3531_n_13765 ( .a(FE_OCP_RBN3527_n_13765), .o(FE_OCP_RBN3531_n_13765) );
in01f80 g748894 ( .a(n_32411), .o(n_32484) );
in01f80 newInst_3537 ( .a(newNet_2938), .o(newNet_3537) );
in01f80 FE_OCP_RBC2396_n_24451 ( .a(n_24451), .o(FE_OCP_RBN2396_n_24451) );
no02f80 g765185 ( .a(FE_OCP_RBN2786_n_15079), .b(FE_OCP_RBN2507_n_13896), .o(n_15159) );
ao22s80 FE_RC_3338_0 ( .a(n_24137), .b(FE_OCP_RBN2277_n_24173), .c(n_24121), .d(n_24173), .o(n_24306) );
in01f80 g752000 ( .a(n_29002), .o(n_29003) );
na02f80 FE_RC_4151_0 ( .a(FE_RN_1805_0), .b(n_22632), .o(n_22674) );
no02f80 g747348 ( .a(n_33575), .b(n_33392), .o(n_33628) );
oa22f80 g749820 ( .a(n_31311), .b(n_31294), .c(n_31530), .d(n_30392), .o(n_31637) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_6_ ( .ck(newNet_2511), .d(n_26807), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_) );
in01f80 g756316 ( .a(n_25129), .o(n_24627) );
na02f80 g752431 ( .a(n_44696), .b(FE_OCP_RBN3306_n_44722), .o(n_27893) );
no02f80 g777840 ( .a(n_3193), .b(n_3177), .o(n_4953) );
no02f80 g743124 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .o(n_37040) );
in01f80 g768731 ( .a(n_12100), .o(n_12101) );
na02f80 g774011 ( .a(n_6861), .b(delay_add_ln22_unr5_stage3_stallmux_q_4_), .o(n_6969) );
no02f80 g741189 ( .a(n_38847), .b(n_38512), .o(n_39004) );
no02f80 g747106 ( .a(n_32799), .b(n_32797), .o(n_32798) );
na02f80 g747681 ( .a(n_32089), .b(n_31879), .o(n_32223) );
no02f80 g738038 ( .a(n_42122), .b(n_42196), .o(n_42123) );
no02f80 g753559 ( .a(n_26722), .b(n_25101), .o(n_26846) );
na02f80 g768497 ( .a(n_12347), .b(n_12389), .o(n_12408) );
in01f80 g769109 ( .a(n_11749), .o(n_11750) );
na02f80 g778718 ( .a(n_2235), .b(n_2494), .o(n_2245) );
in01f80 g752297 ( .a(n_27964), .o(n_27965) );
ao12f80 g756783 ( .a(n_23251), .b(n_23348), .c(n_23252), .o(n_23397) );
na02f80 FE_RC_2418_0 ( .a(FE_RN_955_0), .b(n_7470), .o(FE_RN_956_0) );
no02f80 g750307 ( .a(n_29733), .b(n_29735), .o(n_29734) );
oa22f80 g753411 ( .a(n_26786), .b(n_26750), .c(n_26787), .d(n_26751), .o(n_26853) );
na03f80 FE_RC_1085_0 ( .a(n_29634), .b(n_29528), .c(n_29616), .o(n_29648) );
ao12f80 g765233 ( .a(n_15664), .b(n_15830), .c(n_15666), .o(n_15832) );
in01f80 newInst_2045 ( .a(newNet_2044), .o(newNet_2045) );
na02f80 g757035 ( .a(n_23803), .b(n_23985), .o(n_24025) );
in01f80 newInst_1695 ( .a(newNet_1694), .o(newNet_1695) );
in01f80 FE_OCP_RBC3486_n_2438 ( .a(FE_OCP_RBN2293_n_2438), .o(FE_OCP_RBN3486_n_2438) );
oa22f80 FE_RC_739_0 ( .a(n_45625), .b(n_36186), .c(n_36508), .d(n_36187), .o(n_36592) );
in01f80 FE_OCP_DRV_C1542_n_26125 ( .a(FE_OCP_DRV_N1541_n_26125), .o(FE_OCP_DRV_N1542_n_26125) );
no02f80 g752025 ( .a(n_28168), .b(n_28144), .o(n_28248) );
in01f80 g738284 ( .a(n_41867), .o(n_41868) );
na02f80 g751557 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_18_), .o(n_28508) );
oa12f80 g754129 ( .a(n_26051), .b(n_25984), .c(n_24219), .o(n_26111) );
oa12f80 g772266 ( .a(n_8590), .b(n_8585), .c(n_8642), .o(n_8692) );
na02f80 g759918 ( .a(FE_OCP_RBN3677_n_21051), .b(n_21134), .o(n_21136) );
ao12f80 g761084 ( .a(n_19787), .b(n_19766), .c(n_19991), .o(n_19992) );
ao12f80 g763258 ( .a(n_16782), .b(n_17083), .c(n_16832), .o(n_17237) );
oa12f80 g753696 ( .a(n_26480), .b(n_26479), .c(n_26506), .o(n_26536) );
in01f80 newInst_2505 ( .a(newNet_2050), .o(newNet_2505) );
in01f80 g749455 ( .a(n_30621), .o(n_30640) );
in01f80 g769668 ( .a(n_11362), .o(n_11363) );
in01f80 FE_OCP_RBC2828_n_30731 ( .a(n_30731), .o(FE_OCP_RBN2828_n_30731) );
na02f80 g748228 ( .a(n_31765), .b(n_31773), .o(n_31851) );
in01f80 FE_OCP_RBC2494_n_8641 ( .a(n_8641), .o(FE_OCP_RBN2494_n_8641) );
oa22f80 FE_RC_1309_0 ( .a(n_34622), .b(n_34875), .c(n_34623), .d(n_34901), .o(n_34999) );
in01f80 FE_OCP_RBC3406_n_28597 ( .a(FE_OCP_RBN3404_n_28597), .o(FE_OCP_RBN3406_n_28597) );
in01f80 FE_OFC40_n_45813 ( .a(FE_OFN757_n_45813), .o(FE_OFN40_n_45813) );
in01f80 g780902 ( .a(n_461), .o(n_451) );
na02f80 g751770 ( .a(n_28930), .b(n_28841), .o(n_29246) );
na02f80 g773947 ( .a(n_7011), .b(n_7010), .o(n_7126) );
in01f80 g753601 ( .a(n_26694), .o(n_26695) );
in01f80 g754637 ( .a(n_27246), .o(n_27366) );
no02f80 g760111 ( .a(n_20404), .b(n_20343), .o(n_20406) );
in01f80 newInst_3714 ( .a(newNet_723), .o(newNet_3714) );
no02f80 g742022 ( .a(n_37908), .b(n_44866), .o(n_37976) );
in01f80 newInst_2741 ( .a(newNet_2740), .o(newNet_2741) );
no02f80 g770081 ( .a(n_10950), .b(FE_OCP_RBN2661_n_9292), .o(n_10984) );
no02f80 g776030 ( .a(n_4726), .b(FE_OCP_RBN2723_n_4219), .o(n_4800) );
in01f80 g740110 ( .a(n_40277), .o(n_40278) );
in01f80 g750776 ( .a(n_29196), .o(n_29169) );
in01f80 g755662 ( .a(n_24556), .o(n_24714) );
in01f80 FE_OCPC1741_n_19138 ( .a(n_19138), .o(FE_OCPN1741_n_19138) );
in01f80 FE_RC_1035_0 ( .a(n_23043), .o(FE_RN_297_0) );
no02f80 g737621 ( .a(n_42330), .b(n_42372), .o(n_42428) );
in01f80 newInst_1771 ( .a(newNet_221), .o(newNet_1771) );
in01f80 drc784094 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_45840) );
in01f80 g754483 ( .a(n_25675), .o(n_25653) );
in01f80 g773141 ( .a(n_7667), .o(n_7668) );
oa22f80 g754603 ( .a(FE_OCP_RBN2957_n_26231), .b(n_25686), .c(FE_OCP_RBN2960_n_26231), .d(n_26417), .o(n_26886) );
in01f80 g756608 ( .a(n_23656), .o(n_24067) );
na02f80 g768086 ( .a(FE_OCPN860_n_12880), .b(n_12840), .o(n_13196) );
in01f80 FE_OCP_DRV_C1552_n_19010 ( .a(FE_OCP_DRV_N1551_n_19010), .o(FE_OCP_DRV_N1552_n_19010) );
in01f80 g767893 ( .a(n_13064), .o(n_12996) );
na02f80 g778701 ( .a(n_2365), .b(n_2364), .o(n_2423) );
ao12f80 g737380 ( .a(n_42370), .b(n_42796), .c(n_42359), .o(n_42812) );
in01f80 FE_OCPC1791_n_25044 ( .a(n_25044), .o(FE_OCPN1791_n_25044) );
na02f80 g771127 ( .a(n_9758), .b(n_9617), .o(n_9844) );
ao12f80 g775649 ( .a(n_5035), .b(n_45319), .c(n_5007), .o(n_5236) );
na02f80 g776041 ( .a(n_4837), .b(n_4517), .o(n_4853) );
no02f80 g780610 ( .a(n_713), .b(n_731), .o(n_746) );
na02f80 g781029 ( .a(cos_out_21), .b(FE_OFN1_n_43918), .o(n_342) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_4_ ( .ck(newNet_2059), .d(n_4857), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_) );
in01f80 g781154 ( .a(n_384), .o(n_376) );
in01f80 g771391 ( .a(n_9142), .o(n_9366) );
no02f80 g759629 ( .a(n_20761), .b(n_20760), .o(n_20790) );
na02f80 g764913 ( .a(FE_OCPN994_n_15552), .b(n_14524), .o(n_15648) );
na02f80 FE_RC_2269_0 ( .a(n_25197), .b(n_25162), .o(FE_RN_844_0) );
na02f80 g784395 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46206) );
in01f80 FE_OCPC885_n_42216 ( .a(FE_OCPN884_n_42216), .o(FE_OCPN885_n_42216) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_24_ ( .ck(newNet_3219), .d(n_36544), .o(delay_add_ln22_unr23_stage9_stallmux_q_24_) );
in01f80 newInst_2544 ( .a(newNet_1016), .o(newNet_2544) );
no02f80 g777672 ( .a(n_3462), .b(n_3512), .o(n_3598) );
oa12f80 g742822 ( .a(n_37145), .b(n_37286), .c(n_37036), .o(n_37314) );
na02f80 g767940 ( .a(n_12848), .b(n_12847), .o(n_12890) );
in01f80 g740883 ( .a(n_39844), .o(n_39459) );
no02f80 g770066 ( .a(n_10809), .b(n_10762), .o(n_10884) );
oa12f80 g759480 ( .a(n_20469), .b(n_20595), .c(n_20407), .o(n_20620) );
oa22f80 g748857 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_15_), .c(n_32422), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32881) );
na02f80 g753280 ( .a(n_27110), .b(n_27210), .o(n_27298) );
in01f80 g759175 ( .a(n_21386), .o(n_21387) );
in01f80 FE_OCP_RBC2731_n_4219 ( .a(FE_OCP_RBN2726_n_4219), .o(FE_OCP_RBN2731_n_4219) );
na02f80 g769075 ( .a(n_12157), .b(n_12081), .o(n_12279) );
oa12f80 g773546 ( .a(n_7406), .b(n_7405), .c(n_7404), .o(n_7445) );
na02f80 g771653 ( .a(n_8885), .b(n_7548), .o(n_8886) );
in01f80 g763210 ( .a(n_17433), .o(n_17545) );
na02f80 g759591 ( .a(n_21881), .b(n_21880), .o(n_21882) );
na02f80 g760879 ( .a(n_19365), .b(n_18706), .o(n_19366) );
na02f80 g779615 ( .a(n_1596), .b(n_1613), .o(n_2092) );
no02f80 g764166 ( .a(n_16474), .b(FE_OCP_RBN2679_n_14768), .o(n_16475) );
in01f80 FE_OCP_DRV_C1581_n_35500 ( .a(n_35500), .o(FE_OCP_DRV_N1581_n_35500) );
in01f80 FE_OCP_RBC2990_n_35539 ( .a(FE_OCP_RBN2986_n_35539), .o(FE_OCP_RBN2990_n_35539) );
in01f80 FE_OCP_RBC1144_n_29292 ( .a(n_29292), .o(FE_OCP_RBN1144_n_29292) );
in01f80 g772332 ( .a(n_8755), .o(n_8756) );
in01f80 fopt784716 ( .a(n_17835), .o(n_47195) );
na02f80 g754027 ( .a(n_26952), .b(n_26951), .o(n_26953) );
no02f80 g766599 ( .a(n_14435), .b(n_14392), .o(n_14393) );
in01f80 g739565 ( .a(n_40631), .o(n_40632) );
in01f80 g758405 ( .a(FE_RN_1667_0), .o(n_26663) );
na02f80 g748136 ( .a(n_31805), .b(n_31851), .o(n_31852) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_22_ ( .ck(newNet_815), .d(n_1312), .o(delay_xor_ln21_unr3_stage2_stallmux_q_22_) );
na02f80 g736409 ( .a(n_43800), .b(n_43420), .o(n_43801) );
no02f80 g768453 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .o(n_12396) );
in01f80 newInst_1331 ( .a(newNet_1330), .o(newNet_1331) );
in01f80 newInst_2369 ( .a(newNet_2368), .o(newNet_2369) );
ao12f80 g779479 ( .a(n_2021), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_23_), .o(n_2028) );
in01f80 newInst_2497 ( .a(newNet_2496), .o(newNet_2497) );
in01f80 newInst_324 ( .a(newNet_323), .o(newNet_324) );
ao12f80 g779046 ( .a(n_2041), .b(n_2043), .c(n_2040), .o(n_2346) );
ao22s80 FE_RC_3884_0 ( .a(n_30869), .b(n_30868), .c(n_30867), .d(n_30870), .o(n_30978) );
oa12f80 g763209 ( .a(n_17159), .b(n_17736), .c(n_17462), .o(n_17789) );
na02f80 g761554 ( .a(n_18895), .b(n_18894), .o(n_18896) );
in01f80 newInst_3052 ( .a(newNet_2521), .o(newNet_3052) );
in01f80 g770093 ( .a(n_11057), .o(n_10972) );
in01f80 g771646 ( .a(n_9074), .o(n_9132) );
no02f80 FE_RC_3756_0 ( .a(FE_RN_1650_0), .b(n_40992), .o(n_41030) );
in01f80 newInst_1573 ( .a(newNet_1572), .o(newNet_1573) );
ao12f80 g746844 ( .a(n_32943), .b(n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_19_), .o(n_33505) );
in01f80 g780066 ( .a(n_1225), .o(n_1226) );
oa12f80 g738611 ( .a(n_41616), .b(n_41713), .c(n_41263), .o(n_42132) );
in01f80 FE_OCP_DRV_C3742_n_25400 ( .a(n_25400), .o(FE_OCP_DRV_N3742_n_25400) );
ao12f80 g740028 ( .a(n_39776), .b(n_39861), .c(n_39806), .o(n_39955) );
no02f80 g769864 ( .a(n_11048), .b(n_44453), .o(n_11136) );
na02f80 g741907 ( .a(n_38320), .b(n_38012), .o(n_38356) );
na02f80 g744328 ( .a(n_44211), .b(n_34948), .o(n_35683) );
in01f80 g779371 ( .a(n_1625), .o(n_1707) );
in01f80 FE_OCP_RBC2974_n_5531 ( .a(FE_OCP_RBN2973_n_5531), .o(FE_OCP_RBN2974_n_5531) );
oa22f80 g779858 ( .a(n_44659), .b(n_938), .c(n_44637), .d(n_916), .o(n_1337) );
na02f80 g777311 ( .a(FE_OCP_RBN2692_FE_OCPN843_n_3912), .b(n_4018), .o(n_4106) );
in01f80 newInst_1416 ( .a(newNet_710), .o(newNet_1416) );
no02f80 g756236 ( .a(n_24707), .b(n_24706), .o(n_24708) );
ao12f80 g757279 ( .a(n_23073), .b(n_23072), .c(n_23071), .o(n_24361) );
in01f80 FE_OCP_RBC3629_n_38870 ( .a(FE_OCP_RBN3627_n_38870), .o(FE_OCP_RBN3629_n_38870) );
na02f80 g784119 ( .a(n_7212), .b(n_7211), .o(n_45866) );
in01f80 g752818 ( .a(n_27437), .o(n_27403) );
no02f80 g743965 ( .a(n_35827), .b(n_35826), .o(n_35865) );
oa22f80 g751087 ( .a(n_30303), .b(n_29490), .c(n_30156), .d(n_29935), .o(n_30476) );
oa12f80 g739481 ( .a(n_44769), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n_40893) );
in01f80 g765786 ( .a(n_15005), .o(n_15006) );
no02f80 g761247 ( .a(n_19009), .b(n_19036), .o(n_19101) );
no02f80 g768357 ( .a(n_12542), .b(n_12541), .o(n_12543) );
oa22f80 g754001 ( .a(n_26978), .b(n_26901), .c(n_26950), .d(n_26902), .o(n_27015) );
in01f80 g754691 ( .a(n_26548), .o(n_26639) );
no02f80 g762698 ( .a(n_18235), .b(n_18234), .o(n_18236) );
in01f80 FE_RC_4202_0 ( .a(n_19561), .o(n_19588) );
ao12f80 g755556 ( .a(n_24569), .b(n_24568), .c(n_24567), .o(n_26360) );
na03f80 FE_RC_1013_0 ( .a(n_29018), .b(n_29017), .c(n_28699), .o(n_29038) );
in01f80 g742368 ( .a(n_37916), .o(n_37831) );
na02f80 g771528 ( .a(n_9333), .b(n_9158), .o(n_9377) );
na02f80 g765142 ( .a(n_15971), .b(n_15969), .o(n_16022) );
in01f80 g760357 ( .a(n_20236), .o(n_20237) );
in01f80 FE_OCP_RBC2928_n_39614 ( .a(n_39614), .o(FE_OCP_RBN2928_n_39614) );
no02f80 FE_RC_2967_0 ( .a(FE_OCP_RBN2720_n_9494), .b(n_11017), .o(FE_RN_1296_0) );
no02f80 g777681 ( .a(n_3327), .b(n_3304), .o(n_5109) );
in01f80 g758852 ( .a(n_21730), .o(n_21731) );
no02f80 g779636 ( .a(n_1444), .b(n_1443), .o(n_2128) );
na02f80 FE_RC_6_0 ( .a(FE_RN_0_0), .b(n_1402), .o(FE_RN_2_0) );
ao22s80 g771167 ( .a(n_9374), .b(n_9291), .c(n_9375), .d(n_9290), .o(n_9584) );
no02f80 g770747 ( .a(FE_OCPN3771_n_8669), .b(n_10100), .o(n_10116) );
in01f80 g750914 ( .a(n_31294), .o(n_30392) );
in01f80 newInst_3517 ( .a(newNet_1338), .o(newNet_3517) );
in01f80 g749135 ( .a(n_30956), .o(n_30957) );
no02f80 g780688 ( .a(n_650), .b(n_649), .o(n_651) );
na02f80 g765399 ( .a(n_15022), .b(n_15052), .o(n_15198) );
in01f80 FE_OCP_RBC3532_n_13765 ( .a(FE_OCP_RBN3527_n_13765), .o(FE_OCP_RBN3532_n_13765) );
na02f80 FE_RC_3312_0 ( .a(FE_RN_1456_0), .b(FE_RN_1457_0), .o(FE_RN_1458_0) );
in01f80 g771086 ( .a(n_10070), .o(n_10125) );
na02f80 g767903 ( .a(n_12921), .b(n_46985), .o(n_13025) );
na02f80 g737200 ( .a(n_42971), .b(n_42825), .o(n_42995) );
na02f80 g759234 ( .a(n_21260), .b(n_21342), .o(n_21416) );
na02f80 g751732 ( .a(n_28347), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_), .o(n_28404) );
in01f80 g751481 ( .a(n_28768), .o(n_28769) );
no02f80 g764330 ( .a(n_16235), .b(n_16236), .o(n_16325) );
na02f80 g766518 ( .a(n_14172), .b(n_14222), .o(n_16143) );
in01f80 g771723 ( .a(n_8992), .o(n_9041) );
in01f80 g751477 ( .a(n_28643), .o(n_28644) );
no02f80 g748905 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .o(n_32498) );
in01f80 FE_OCPC3770_n_8669 ( .a(n_8669), .o(FE_OCPN3770_n_8669) );
na02f80 g766372 ( .a(n_14653), .b(n_14040), .o(n_14701) );
na02f80 g744881 ( .a(n_35001), .b(n_30504), .o(n_35034) );
in01f80 FE_RC_1942_0 ( .a(n_12956), .o(FE_RN_619_0) );
oa22f80 g739829 ( .a(n_40417), .b(n_40315), .c(n_40418), .d(n_40314), .o(n_40458) );
in01f80 FE_OCP_RBC2236_n_29055 ( .a(n_29055), .o(FE_OCP_RBN2236_n_29055) );
oa22f80 g737267 ( .a(n_42871), .b(n_42525), .c(n_42857), .d(n_42524), .o(n_43299) );
na02f80 g738942 ( .a(n_41171), .b(n_40943), .o(n_41202) );
in01f80 g774378 ( .a(n_6920), .o(n_6921) );
oa22f80 FE_RC_584_0 ( .a(n_42086), .b(n_41766), .c(n_41767), .d(n_42085), .o(n_42144) );
no02f80 g745105 ( .a(n_34661), .b(n_34375), .o(n_34711) );
in01f80 fopt782791 ( .a(n_44211), .o(n_44180) );
in01f80 FE_OCP_RBC3827_n_18951 ( .a(n_18951), .o(FE_OCP_RBN3827_n_18951) );
in01f80 g739760 ( .a(n_40526), .o(n_40527) );
ao12f80 g761752 ( .a(n_19294), .b(n_19293), .c(n_19292), .o(n_19790) );
no02f80 g778618 ( .a(n_2592), .b(n_2545), .o(n_3071) );
na02f80 g761067 ( .a(n_20115), .b(n_20114), .o(n_20116) );
in01f80 g752713 ( .a(n_27362), .o(n_27358) );
na02f80 g772928 ( .a(n_8091), .b(n_7730), .o(n_8094) );
ao12f80 g780692 ( .a(n_645), .b(n_647), .c(n_497), .o(n_650) );
in01f80 g766597 ( .a(n_13922), .o(n_13923) );
ao12f80 g772029 ( .a(n_8081), .b(n_8852), .c(n_8110), .o(n_8932) );
in01f80 g772327 ( .a(n_8719), .o(n_8720) );
oa12f80 g742582 ( .a(n_37573), .b(n_37572), .c(n_37571), .o(n_37637) );
no02f80 g747670 ( .a(n_33243), .b(n_33258), .o(n_33297) );
ao12f80 g765107 ( .a(n_16101), .b(n_16100), .c(n_16245), .o(n_16259) );
na02f80 g773702 ( .a(n_7263), .b(n_7305), .o(n_7309) );
in01f80 g775113 ( .a(n_5946), .o(n_5976) );
ao12f80 g763026 ( .a(n_17641), .b(n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_8_), .o(n_17741) );
in01f80 newInst_1867 ( .a(newNet_1866), .o(newNet_1867) );
in01f80 g766140 ( .a(n_14600), .o(n_14601) );
in01f80 g757923 ( .a(n_23083), .o(n_23084) );
no02f80 g746077 ( .a(n_44842), .b(FE_OCP_RBN2284_n_33846), .o(n_33921) );
in01f80 g749697 ( .a(n_31578), .o(n_31579) );
na02f80 g759294 ( .a(n_20858), .b(n_45010), .o(n_20980) );
na02f80 g743415 ( .a(n_37787), .b(n_46248), .o(n_37788) );
in01f80 g771602 ( .a(n_9333), .o(n_9396) );
no02f80 g738435 ( .a(n_41452), .b(n_41409), .o(n_41518) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_3_ ( .ck(newNet_1372), .d(n_36282), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_) );
na02f80 g775907 ( .a(n_5217), .b(n_4868), .o(n_5351) );
no04s80 g756912 ( .a(n_23308), .b(FE_OCPN1017_n_23307), .c(FE_OCPN1022_n_23195), .d(n_23077), .o(n_23328) );
no02f80 FE_RC_1121_0 ( .a(n_2438), .b(FE_RN_338_0), .o(n_44059) );
oa12f80 g738269 ( .a(n_41512), .b(n_41776), .c(n_41548), .o(n_41931) );
in01f80 g753930 ( .a(n_26265), .o(n_26266) );
in01f80 fopt782912 ( .a(n_22705), .o(n_44364) );
na02f80 g762269 ( .a(n_18810), .b(n_18809), .o(n_19292) );
no02f80 g776844 ( .a(n_3850), .b(n_3809), .o(n_3978) );
oa12f80 g752765 ( .a(n_27812), .b(n_27763), .c(n_179), .o(n_27909) );
ao12f80 g754394 ( .a(n_25782), .b(n_25704), .c(n_25504), .o(n_25812) );
na02f80 g759286 ( .a(n_20995), .b(n_21077), .o(n_21078) );
na02f80 g743167 ( .a(n_36888), .b(n_36936), .o(n_36919) );
in01f80 g745892 ( .a(n_35391), .o(n_35371) );
in01f80 g776120 ( .a(n_4837), .o(n_4838) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_3_ ( .ck(newNet_412), .d(n_32511), .o(delay_xor_ln22_unr21_stage8_stallmux_q_3_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_25_ ( .ck(newNet_1599), .d(n_27539), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_) );
no02f80 g742486 ( .a(n_37516), .b(n_37119), .o(n_37564) );
na02f80 g758942 ( .a(n_21281), .b(FE_OCPN1524_n_45072), .o(n_21328) );
in01f80 g750471 ( .a(n_29590), .o(n_29602) );
in01f80 g755447 ( .a(n_24851), .o(n_24852) );
no02f80 g750854 ( .a(n_30235), .b(n_30233), .o(n_30267) );
in01f80 g771589 ( .a(n_8989), .o(n_9189) );
in01f80 FE_OCP_RBC1156_n_18375 ( .a(FE_OCP_RBN1155_n_18375), .o(FE_OCP_RBN1156_n_18375) );
in01f80 g738311 ( .a(n_42191), .o(n_41886) );
na02f80 g753443 ( .a(n_26961), .b(n_26879), .o(n_26962) );
in01f80 newInst_1425 ( .a(newNet_242), .o(newNet_1425) );
in01f80 FE_OCP_RBC3724_n_16975 ( .a(n_16975), .o(FE_OCP_RBN3724_n_16975) );
no02f80 g766441 ( .a(n_14181), .b(n_14154), .o(n_14182) );
in01f80 g781395 ( .a(beta_11), .o(n_51) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_11_ ( .ck(newNet_1347), .d(n_1136), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_) );
oa12f80 g746633 ( .a(n_34473), .b(n_34580), .c(n_34579), .o(n_34581) );
na02f80 g770054 ( .a(n_10850), .b(n_10831), .o(n_10876) );
ao22s80 FE_RC_701_0 ( .a(n_40646), .b(n_40652), .c(n_40651), .d(n_40650), .o(n_40686) );
no02f80 g743977 ( .a(n_36148), .b(n_36147), .o(n_36196) );
no02f80 g747472 ( .a(FE_OCP_RBN3332_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .o(n_32522) );
no02f80 g769347 ( .a(FE_OCP_RBN2002_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_12003) );
in01f80 newInst_3745 ( .a(newNet_3744), .o(newNet_3745) );
in01f80 FE_OCP_RBC2715_n_14982 ( .a(FE_OCP_RBN2714_n_14982), .o(FE_OCP_RBN2715_n_14982) );
ao12f80 g768931 ( .a(n_12043), .b(FE_OCPN867_n_45697), .c(delay_xor_ln21_unr9_stage4_stallmux_q_11_), .o(n_12110) );
na02f80 g779315 ( .a(n_1787), .b(n_1741), .o(n_1697) );
na02f80 g758086 ( .a(n_44268), .b(FE_OCPN1502_n_20723), .o(n_22229) );
in01f80 FE_OCP_RBC3518_n_8498 ( .a(FE_OCP_RBN3517_n_8498), .o(FE_OCP_RBN3518_n_8498) );
na02f80 g767801 ( .a(n_13252), .b(n_13251), .o(n_13253) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_22_ ( .ck(newNet_3046), .d(n_1189), .o(delay_add_ln22_unr2_stage2_stallmux_q_22_) );
oa12f80 g765580 ( .a(n_14488), .b(n_15446), .c(n_14456), .o(n_15521) );
in01f80 FE_OCP_RBC3671_FE_RN_470_0 ( .a(FE_RN_470_0), .o(FE_OCP_RBN3671_FE_RN_470_0) );
no02f80 g741495 ( .a(n_38765), .b(n_38764), .o(n_38772) );
in01f80 g768255 ( .a(n_12714), .o(n_12715) );
na02f80 g745705 ( .a(n_34189), .b(n_34191), .o(n_34190) );
na02f80 g740610 ( .a(n_39640), .b(n_39639), .o(n_39743) );
na02f80 g780617 ( .a(n_679), .b(n_701), .o(n_697) );
no02f80 g740239 ( .a(n_39973), .b(n_39940), .o(n_39971) );
in01f80 g762383 ( .a(n_18664), .o(n_18490) );
in01f80 FE_OCPC1746_n_29420 ( .a(FE_OCPN1745_n_29420), .o(FE_OCPN1746_n_29420) );
in01f80 g741615 ( .a(n_38627), .o(n_38641) );
ao12f80 g760492 ( .a(n_19772), .b(n_19976), .c(n_19975), .o(n_20003) );
na02f80 g773851 ( .a(n_7022), .b(n_5619), .o(n_7092) );
in01f80 g773013 ( .a(n_7784), .o(n_7785) );
ao12f80 g754584 ( .a(n_26716), .b(FE_OCP_RBN2960_n_26231), .c(n_26348), .o(n_26908) );
in01f80 g760304 ( .a(n_20244), .o(n_20262) );
in01f80 FE_OCP_RBC2538_n_3645 ( .a(n_3645), .o(FE_OCP_RBN2538_n_3645) );
na02f80 FE_RC_2446_0 ( .a(FE_RN_976_0), .b(n_13393), .o(n_13462) );
in01f80 g760516 ( .a(n_19997), .o(n_19998) );
no02f80 g739236 ( .a(n_40692), .b(n_41008), .o(n_41089) );
oa12f80 g749819 ( .a(n_30977), .b(n_30976), .c(n_30975), .o(n_31410) );
in01f80 newInst_1322 ( .a(newNet_1321), .o(newNet_1322) );
na02f80 g775331 ( .a(n_5752), .b(n_5744), .o(n_5816) );
in01f80 g778868 ( .a(n_2741), .o(n_2759) );
no02f80 g774752 ( .a(n_6319), .b(n_6322), .o(n_6320) );
na02f80 FE_RC_3643_0 ( .a(n_31273), .b(FE_RN_1598_0), .o(n_31305) );
na02f80 g750117 ( .a(FE_OCP_RBN2573_n_29922), .b(n_45758), .o(n_30371) );
no02f80 g764835 ( .a(n_15792), .b(FE_OFN823_n_15791), .o(n_15843) );
no02f80 g766943 ( .a(n_14758), .b(n_14257), .o(n_14350) );
na02f80 g753882 ( .a(n_27034), .b(n_26885), .o(n_27066) );
na02f80 g772652 ( .a(n_8229), .b(FE_OCPN891_n_7802), .o(n_8250) );
oa12f80 g741347 ( .a(n_38798), .b(n_38801), .c(n_38797), .o(n_39745) );
in01f80 g774770 ( .a(n_6347), .o(n_6348) );
na02f80 g761935 ( .a(n_18268), .b(n_17556), .o(n_18366) );
in01f80 g746298 ( .a(n_34200), .o(n_33686) );
no02f80 g751355 ( .a(n_29410), .b(n_29409), .o(n_29411) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_0_ ( .ck(newNet_2034), .d(n_9428), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_0_) );
na02f80 g744016 ( .a(n_36190), .b(n_36143), .o(n_36299) );
na02f80 g754283 ( .a(n_25832), .b(n_45532), .o(n_25916) );
in01f80 g764867 ( .a(n_15591), .o(n_15592) );
no02f80 g772780 ( .a(n_7943), .b(n_7415), .o(n_7972) );
na02f80 FE_RC_4083_0 ( .a(FE_RN_1784_0), .b(n_16912), .o(FE_RN_1783_0) );
in01f80 newInst_1879 ( .a(newNet_1878), .o(newNet_1879) );
no02f80 g741978 ( .a(n_37946), .b(n_37939), .o(n_37986) );
in01f80 newInst_489 ( .a(newNet_337), .o(newNet_489) );
in01f80 g781341 ( .a(n_86), .o(n_87) );
na02f80 g764502 ( .a(n_16269), .b(n_16268), .o(n_16270) );
in01f80 FE_RC_1899_0 ( .a(n_11813), .o(FE_RN_594_0) );
no02f80 g739412 ( .a(FE_OCPN897_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n_40981) );
no02f80 g737448 ( .a(n_42654), .b(n_42306), .o(n_42703) );
oa22f80 g744558 ( .a(n_36623), .b(n_36169), .c(n_36642), .d(n_36170), .o(n_36698) );
oa12f80 g768722 ( .a(n_11613), .b(n_12024), .c(n_11656), .o(n_12023) );
ao22s80 FE_RC_1464_0 ( .a(n_27501), .b(n_27648), .c(n_27500), .d(n_27649), .o(n_27729) );
no02f80 g769085 ( .a(n_11497), .b(n_11517), .o(n_11700) );
oa12f80 g744501 ( .a(n_35317), .b(n_35414), .c(n_35351), .o(n_35460) );
no02f80 g758371 ( .a(n_22187), .b(n_21166), .o(n_22383) );
in01f80 g754364 ( .a(n_25819), .o(n_25820) );
in01f80 newInst_1861 ( .a(newNet_338), .o(newNet_1861) );
no02f80 g763937 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n_17462) );
na02f80 g766785 ( .a(n_13691), .b(n_13706), .o(n_13836) );
no02f80 g769195 ( .a(n_12077), .b(n_12076), .o(n_12678) );
no02f80 g748157 ( .a(n_31869), .b(n_31864), .o(n_31906) );
in01f80 FE_OCP_RBC2197_n_12830 ( .a(n_12830), .o(FE_OCP_RBN2197_n_12830) );
na02f80 g749853 ( .a(FE_OCP_RBN3012_n_31117), .b(n_30615), .o(n_31285) );
na02f80 g763928 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .o(n_17155) );
oa12f80 g775784 ( .a(n_4612), .b(n_5339), .c(n_4685), .o(n_5432) );
no02f80 g738187 ( .a(n_42009), .b(n_42008), .o(n_42010) );
no02f80 g737043 ( .a(n_43171), .b(n_43104), .o(n_43223) );
na02f80 g752347 ( .a(n_28435), .b(n_28434), .o(n_28436) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_21_ ( .ck(newNet_3048), .d(n_1168), .o(delay_add_ln22_unr2_stage2_stallmux_q_21_) );
in01f80 fopt783050 ( .a(n_44490), .o(n_44498) );
no02f80 g744991 ( .a(n_34971), .b(n_34652), .o(n_34972) );
in01f80 newInst_1930 ( .a(newNet_1929), .o(newNet_1930) );
na02f80 g749874 ( .a(FE_OCP_RBN3010_n_31117), .b(n_31039), .o(n_31394) );
no02f80 g763923 ( .a(FE_OCP_RBN3294_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_), .o(n_17096) );
no02f80 g750326 ( .a(n_29673), .b(n_45760), .o(n_29705) );
na02f80 g756579 ( .a(n_23606), .b(n_22754), .o(n_23762) );
ao22s80 g775468 ( .a(n_5695), .b(n_5466), .c(n_5696), .d(n_5465), .o(n_5820) );
in01f80 newInst_3113 ( .a(newNet_3112), .o(newNet_3113) );
in01f80 g754217 ( .a(n_26136), .o(n_26076) );
ao12f80 g772054 ( .a(n_8531), .b(n_8471), .c(n_7594), .o(n_8532) );
na02f80 g745622 ( .a(n_34286), .b(n_34560), .o(n_34650) );
in01f80 FE_OCP_DRV_C1600_n_21493 ( .a(FE_OCP_DRV_N1599_n_21493), .o(FE_OCP_DRV_N1600_n_21493) );
in01f80 newInst_440 ( .a(newNet_433), .o(newNet_440) );
na02f80 g737253 ( .a(n_42936), .b(n_42956), .o(n_42957) );
in01f80 g740400 ( .a(n_39964), .o(n_40033) );
in01f80 g737234 ( .a(n_42962), .o(n_43300) );
in01f80 g776569 ( .a(n_4350), .o(n_4351) );
na02f80 g767656 ( .a(n_13259), .b(n_13084), .o(n_13326) );
na02f80 g759974 ( .a(n_20435), .b(n_45101), .o(n_20500) );
no02f80 g739924 ( .a(n_40436), .b(n_40097), .o(n_40438) );
na02f80 g774051 ( .a(n_6957), .b(n_6956), .o(n_6958) );
na02f80 g753110 ( .a(n_27455), .b(n_27527), .o(n_27546) );
no02f80 g774857 ( .a(n_6266), .b(n_6250), .o(n_6315) );
in01f80 FE_RC_2878_0 ( .a(FE_RN_1244_0), .o(n_14472) );
no02f80 g759924 ( .a(FE_OCP_RBN3677_n_21051), .b(n_21294), .o(n_21247) );
na02f80 g775590 ( .a(n_5551), .b(n_5520), .o(n_5521) );
oa12f80 g780144 ( .a(n_1111), .b(n_1170), .c(n_936), .o(n_1181) );
na02f80 g751312 ( .a(n_29636), .b(n_29130), .o(n_29675) );
oa12f80 g745350 ( .a(n_35723), .b(FE_OCP_RBN2995_n_35539), .c(n_35653), .o(n_36157) );
na02f80 g756274 ( .a(n_24668), .b(n_24667), .o(n_24669) );
in01f80 g778561 ( .a(n_3058), .o(n_3125) );
in01f80 newInst_1199 ( .a(newNet_913), .o(newNet_1199) );
oa12f80 g747692 ( .a(n_33699), .b(n_33571), .c(n_33684), .o(n_34419) );
in01f80 g773593 ( .a(n_7399), .o(n_7400) );
na02f80 g778098 ( .a(n_2987), .b(n_2865), .o(n_3016) );
na02f80 g771347 ( .a(n_9549), .b(n_9610), .o(n_9791) );
no03m80 FE_RC_1722_0 ( .a(n_28145), .b(n_28226), .c(FE_RN_476_0), .o(n_28271) );
na02f80 g737338 ( .a(n_42833), .b(n_42388), .o(n_42860) );
ao12f80 g762601 ( .a(n_17709), .b(n_45524), .c(n_17531), .o(n_18383) );
in01f80 g749509 ( .a(n_30598), .o(n_30597) );
na02f80 g773238 ( .a(n_8635), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n_8699) );
in01f80 g737655 ( .a(n_42815), .o(n_42816) );
oa22f80 g757874 ( .a(n_22169), .b(n_21971), .c(n_22140), .d(n_21972), .o(n_22359) );
na02f80 g761295 ( .a(n_19030), .b(n_19004), .o(n_19139) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_7_ ( .ck(newNet_3187), .d(n_35791), .o(delay_add_ln22_unr23_stage9_stallmux_q_7_) );
na02f80 g772791 ( .a(n_8175), .b(n_8174), .o(n_8208) );
in01f80 g749081 ( .a(n_32249), .o(n_32250) );
in01f80 g759251 ( .a(n_21305), .o(n_21384) );
in01f80 FE_RC_2414_0 ( .a(n_7095), .o(FE_RN_953_0) );
no03m80 FE_RC_1047_0 ( .a(n_1435), .b(n_1494), .c(n_1427), .o(n_1513) );
in01f80 g745535 ( .a(n_34562), .o(n_34563) );
ao12f80 g742364 ( .a(n_37807), .b(n_37806), .c(n_37817), .o(n_38752) );
oa12f80 g746125 ( .a(n_33450), .b(n_33772), .c(n_33379), .o(n_33898) );
in01f80 newInst_3104 ( .a(newNet_3103), .o(newNet_3104) );
no02f80 g779543 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_13_), .o(n_1706) );
no02f80 g767896 ( .a(n_12990), .b(FE_OCPN860_n_12880), .o(n_13040) );
na02f80 g783832 ( .a(n_32090), .b(n_31880), .o(n_45517) );
in01f80 g748727 ( .a(n_31329), .o(n_31358) );
ao12f80 g756888 ( .a(n_23803), .b(n_24086), .c(n_24088), .o(n_24151) );
na02f80 g759595 ( .a(n_20793), .b(n_20761), .o(n_20794) );
in01f80 g765762 ( .a(n_15103), .o(n_15142) );
no02f80 g775226 ( .a(n_5905), .b(n_5707), .o(n_5970) );
no02f80 g738378 ( .a(n_41770), .b(n_41727), .o(n_41789) );
in01f80 g744359 ( .a(n_46222), .o(n_36822) );
oa22f80 g737878 ( .a(n_42270), .b(n_42107), .c(FE_OCPN1231_n_42201), .d(n_42081), .o(n_42610) );
in01f80 g775337 ( .a(n_5735), .o(n_5809) );
in01f80 FE_RC_2914_0 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(FE_RN_1268_0) );
in01f80 FE_OCP_RBC2972_n_31239 ( .a(n_31239), .o(FE_OCP_RBN2972_n_31239) );
in01f80 newInst_88 ( .a(newNet_87), .o(newNet_88) );
in01f80 g778066 ( .a(n_3061), .o(n_3062) );
in01f80 g743373 ( .a(n_36720), .o(n_36721) );
oa12f80 g750256 ( .a(n_29615), .b(n_29808), .c(FE_OCP_RBN3526_n_29624), .o(n_29831) );
na02f80 g759624 ( .a(n_20598), .b(n_20317), .o(n_20648) );
no02f80 g738120 ( .a(n_42105), .b(n_41617), .o(n_42082) );
in01f80 g736867 ( .a(n_43539), .o(n_43540) );
in01f80 newInst_3664 ( .a(newNet_3248), .o(newNet_3664) );
oa22f80 g738460 ( .a(n_41660), .b(n_41275), .c(FE_OCPN952_n_41540), .d(n_41631), .o(n_41851) );
in01f80 newInst_1543 ( .a(newNet_1542), .o(newNet_1543) );
oa22f80 FE_RC_1307_0 ( .a(n_14659), .b(n_14560), .c(n_14485), .d(n_14660), .o(n_14763) );
na02f80 g754040 ( .a(n_26117), .b(n_26175), .o(n_26202) );
na03f80 FE_RC_3678_0 ( .a(n_6236), .b(n_6354), .c(n_6386), .o(n_6416) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_3_ ( .ck(newNet_2445), .d(n_31326), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_) );
no02f80 g758812 ( .a(n_21731), .b(n_21538), .o(n_21787) );
na02f80 g775836 ( .a(n_5373), .b(n_5431), .o(n_5463) );
na02f80 g773766 ( .a(n_7202), .b(n_5999), .o(n_7252) );
in01f80 g762346 ( .a(n_18725), .o(n_18808) );
na02f80 g737951 ( .a(n_42201), .b(n_41954), .o(n_42359) );
no02f80 g738983 ( .a(n_41205), .b(n_41206), .o(n_41238) );
no02f80 g759676 ( .a(n_20349), .b(n_20281), .o(n_20383) );
na02f80 g760208 ( .a(FE_OCP_RBN1332_n_20249), .b(FE_OCPN1044_n_20307), .o(n_20333) );
in01f80 g764187 ( .a(n_16499), .o(n_16472) );
na02f80 g761334 ( .a(n_19848), .b(n_19845), .o(n_19906) );
oa22f80 g765996 ( .a(FE_OCPN971_n_14716), .b(n_13563), .c(n_14707), .d(n_13562), .o(n_14809) );
in01f80 g775209 ( .a(n_6062), .o(n_6024) );
in01f80 FE_OCPC1235_n_32791 ( .a(n_32791), .o(FE_OCPN1235_n_32791) );
na02f80 g739141 ( .a(n_41041), .b(n_41040), .o(n_41042) );
in01f80 FE_OCP_RBC2847_n_39479 ( .a(n_39479), .o(FE_OCP_RBN2847_n_39479) );
na02f80 g745074 ( .a(n_34754), .b(n_34481), .o(n_34792) );
in01f80 g751565 ( .a(n_28631), .o(n_28565) );
no02f80 g784729 ( .a(n_11962), .b(n_11643), .o(n_47212) );
na02f80 g740857 ( .a(n_39347), .b(n_39254), .o(n_39381) );
in01f80 g761729 ( .a(n_18824), .o(n_18791) );
in01f80 g767842 ( .a(n_13015), .o(n_12928) );
no02f80 g773024 ( .a(n_7761), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n_7762) );
in01f80 newInst_2823 ( .a(newNet_2822), .o(newNet_2823) );
na02f80 g742846 ( .a(n_37165), .b(n_36975), .o(n_37196) );
in01f80 g770026 ( .a(n_10917), .o(n_10918) );
ao22s80 g762304 ( .a(n_18087), .b(n_18036), .c(n_18130), .d(n_18037), .o(n_19751) );
in01f80 newInst_787 ( .a(newNet_786), .o(newNet_787) );
no02f80 g748525 ( .a(n_31677), .b(n_31676), .o(n_31698) );
no02f80 g740383 ( .a(n_39803), .b(n_39513), .o(n_39939) );
no02f80 g762745 ( .a(FE_OCP_RBN2148_FE_OCPN861_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .o(n_17872) );
in01f80 g750571 ( .a(n_30214), .o(n_29472) );
na02f80 FE_RC_2002_0 ( .a(FE_RN_657_0), .b(n_20062), .o(n_20075) );
na02f80 FE_RC_492_0 ( .a(FE_RN_146_0), .b(n_28458), .o(n_28632) );
na03f80 FE_RC_2438_0 ( .a(n_32709), .b(FE_RN_972_0), .c(n_46413), .o(n_32713) );
ao12f80 FE_RC_2645_0 ( .a(FE_RN_1103_0), .b(n_23172), .c(n_23173), .o(n_23248) );
no02f80 g758789 ( .a(n_21510), .b(n_21509), .o(n_21619) );
in01f80 fopt783569 ( .a(n_3161), .o(n_45190) );
oa12f80 g743556 ( .a(n_46206), .b(n_37586), .c(n_46213), .o(n_37634) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_22_ ( .ck(newNet_1608), .d(n_27448), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_) );
in01f80 newInst_1217 ( .a(newNet_56), .o(newNet_1217) );
no02f80 g777216 ( .a(n_3599), .b(n_3646), .o(n_3784) );
in01f80 g747876 ( .a(n_32214), .o(n_32215) );
ao12f80 g748447 ( .a(n_32587), .b(n_32677), .c(n_32482), .o(n_32766) );
in01f80 newInst_2756 ( .a(newNet_2755), .o(newNet_2756) );
no02f80 g769097 ( .a(n_11482), .b(n_11313), .o(n_11484) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_23_ ( .ck(newNet_3308), .d(n_32311), .o(delay_add_ln22_unr20_stage8_stallmux_q_23_) );
oa22f80 FE_RC_1169_0 ( .a(n_12117), .b(FE_OFN802_n_46285), .c(FE_OFN771_n_46337), .d(n_12113), .o(n_46352) );
ao12f80 g757913 ( .a(n_22186), .b(n_22388), .c(n_22269), .o(n_22448) );
na02f80 g766279 ( .a(n_14165), .b(n_14203), .o(n_14204) );
no02f80 FE_RC_1958_0 ( .a(FE_RN_1654_0), .b(FE_RN_630_0), .o(FE_RN_631_0) );
no02f80 g744040 ( .a(n_44223), .b(n_34724), .o(n_36297) );
oa22f80 FE_RC_3449_0 ( .a(n_29704), .b(n_29788), .c(n_29763), .d(n_29717), .o(n_29845) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_6_ ( .ck(newNet_2705), .d(n_15722), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_) );
no02f80 g743051 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_37019) );
in01f80 newInst_1517 ( .a(newNet_1516), .o(newNet_1517) );
na02f80 g746493 ( .a(n_34500), .b(n_34526), .o(n_34587) );
na02f80 g751417 ( .a(n_28477), .b(n_28454), .o(n_28455) );
in01f80 newInst_2651 ( .a(newNet_2650), .o(newNet_2651) );
no02f80 g764698 ( .a(n_15808), .b(n_15806), .o(n_15807) );
no02f80 g741727 ( .a(n_38502), .b(n_38501), .o(n_38503) );
in01f80 newInst_3077 ( .a(newNet_3076), .o(newNet_3077) );
oa22f80 g780037 ( .a(n_1243), .b(n_1059), .c(n_1242), .d(n_1060), .o(n_1249) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_7_ ( .ck(newNet_2509), .d(n_26853), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_) );
in01f80 g742626 ( .a(n_37467), .o(n_37488) );
in01f80 newInst_2161 ( .a(newNet_990), .o(newNet_2161) );
ao12f80 g746848 ( .a(n_32949), .b(FE_OCP_RBN2169_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(n_33301) );
in01f80 newInst_125 ( .a(newNet_124), .o(newNet_125) );
na02f80 g771943 ( .a(n_8696), .b(FE_OCP_RBN3467_n_7886), .o(n_8698) );
na02f80 FE_RC_462_0 ( .a(FE_RN_141_0), .b(FE_RN_133_0), .o(FE_RN_134_0) );
in01f80 g777904 ( .a(n_3220), .o(n_3221) );
oa12f80 g750682 ( .a(n_30360), .b(n_30359), .c(n_30358), .o(n_30416) );
na02f80 g775257 ( .a(n_5667), .b(n_5655), .o(n_5707) );
na02f80 g766023 ( .a(n_14971), .b(n_14742), .o(n_14744) );
no02f80 g742126 ( .a(n_37868), .b(n_37905), .o(n_37989) );
no02f80 g763080 ( .a(n_17483), .b(n_17515), .o(n_17484) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_16_ ( .ck(newNet_739), .d(n_46149), .o(delay_xor_ln21_unr6_stage3_stallmux_q_16_) );
oa22f80 g749287 ( .a(n_32063), .b(n_31629), .c(n_32035), .d(n_31630), .o(n_32173) );
no02f80 g768797 ( .a(n_12020), .b(n_12091), .o(n_12174) );
in01f80 newInst_328 ( .a(newNet_327), .o(newNet_328) );
oa22f80 g779896 ( .a(n_44652), .b(n_1017), .c(n_44661), .d(n_972), .o(n_1335) );
in01f80 g755498 ( .a(n_24820), .o(n_24821) );
in01f80 g776698 ( .a(n_4273), .o(n_4274) );
na02f80 g744308 ( .a(FE_OCP_RBN2903_n_44174), .b(n_35092), .o(n_36088) );
in01f80 FE_OCPC1775_n_18263 ( .a(n_18263), .o(FE_OCPN1775_n_18263) );
no02f80 FE_RC_154_0 ( .a(FE_RN_47_0), .b(n_17890), .o(n_17996) );
na02f80 g769776 ( .a(n_11235), .b(n_11152), .o(n_11262) );
in01f80 FE_OCP_RBC1200_n_25763 ( .a(n_25763), .o(FE_OCP_RBN1200_n_25763) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_1_ ( .ck(newNet_639), .d(n_46384), .o(delay_xor_ln21_unr9_stage4_stallmux_q_1_) );
in01f80 FE_RC_2709_0 ( .a(n_12547), .o(FE_RN_1140_0) );
na02f80 g769704 ( .a(n_11374), .b(n_11306), .o(n_11359) );
in01f80 newInst_2866 ( .a(newNet_2865), .o(newNet_2866) );
no02f80 g776055 ( .a(n_5110), .b(n_5109), .o(n_5153) );
ao12f80 g757270 ( .a(n_23023), .b(n_44066), .c(delay_xor_ln22_unr15_stage6_stallmux_q_8_), .o(n_23047) );
in01f80 FE_OCPC1005_n_13962 ( .a(FE_OCP_RBN2507_n_13896), .o(FE_OCPN1005_n_13962) );
na02f80 g738469 ( .a(n_41387), .b(n_41415), .o(n_41825) );
in01f80 FE_OCP_RBC3421_n_12879 ( .a(n_12879), .o(FE_OCP_RBN3421_n_12879) );
in01f80 FE_OCP_DRV_C1577_n_33904 ( .a(n_33904), .o(FE_OCP_DRV_N1577_n_33904) );
in01f80 g774508 ( .a(n_6703), .o(n_6664) );
na02f80 g769038 ( .a(n_11696), .b(n_45224), .o(n_11697) );
oa22f80 g778748 ( .a(n_2338), .b(n_2029), .c(n_2381), .d(n_2028), .o(n_2476) );
na02f80 g771979 ( .a(FE_OCP_RBN3644_n_44490), .b(n_9767), .o(n_9873) );
in01f80 FE_RC_557_0 ( .a(n_30281), .o(FE_RN_168_0) );
in01f80 g757807 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_16_), .o(n_23560) );
no02f80 g779607 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .o(n_2073) );
no02f80 g745171 ( .a(n_34493), .b(n_34204), .o(n_34574) );
in01f80 g778778 ( .a(n_45903), .o(n_2235) );
no02f80 g763068 ( .a(n_17863), .b(n_17426), .o(n_17905) );
ao12f80 g772297 ( .a(n_8604), .b(n_8620), .c(FE_OCP_RBN3465_n_7886), .o(n_8730) );
no02f80 g766067 ( .a(n_14993), .b(n_14992), .o(n_14994) );
oa22f80 FE_RC_3127_0 ( .a(n_27536), .b(n_31239), .c(n_27366), .d(FE_OCP_RBN2971_n_31239), .o(n_31360) );
na02f80 g771887 ( .a(n_8860), .b(n_8770), .o(n_8861) );
no02f80 g758982 ( .a(n_21202), .b(n_21126), .o(n_21240) );
na02f80 g773979 ( .a(FE_OCP_RBN3376_n_6822), .b(n_6831), .o(n_6908) );
in01f80 FE_OCPC860_n_12880 ( .a(FE_OCPN859_n_12880), .o(FE_OCPN860_n_12880) );
in01f80 g778908 ( .a(n_2338), .o(n_2381) );
no02f80 g773109 ( .a(n_7682), .b(n_7727), .o(n_7786) );
na02f80 g780429 ( .a(n_943), .b(n_926), .o(n_1020) );
na02f80 g778548 ( .a(n_2712), .b(n_2662), .o(n_2713) );
oa22f80 g758637 ( .a(n_22397), .b(n_21861), .c(n_22430), .d(n_21862), .o(n_22545) );
no02f80 g755865 ( .a(n_25056), .b(n_25029), .o(n_25057) );
in01f80 FE_OCP_RBC2361_n_13818 ( .a(FE_OCP_RBN3496_n_13818), .o(FE_OCP_RBN2361_n_13818) );
oa12f80 g750963 ( .a(n_30231), .b(n_30182), .c(n_30156), .o(n_30975) );
in01f80 FE_OCP_RBC2837_FE_RN_745_0 ( .a(FE_RN_745_0), .o(FE_OCP_RBN2837_FE_RN_745_0) );
oa12f80 g773572 ( .a(n_7418), .b(n_7417), .c(n_7416), .o(n_8444) );
in01f80 g771190 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .o(n_11542) );
oa12f80 g775555 ( .a(n_5521), .b(n_5551), .c(n_5520), .o(n_5645) );
no02f80 g761472 ( .a(n_19647), .b(n_19677), .o(n_19761) );
in01f80 g750800 ( .a(FE_OCP_RBN3436_n_29163), .o(n_30136) );
in01f80 g770888 ( .a(n_10050), .o(n_10051) );
na02f80 FE_RC_2872_0 ( .a(n_29059), .b(n_30399), .o(FE_RN_1240_0) );
no02f80 g753091 ( .a(n_27188), .b(n_27146), .o(n_27274) );
in01f80 g764766 ( .a(n_15768), .o(n_15812) );
no02f80 g765188 ( .a(n_15198), .b(n_14210), .o(n_15233) );
na02f80 g754983 ( .a(n_25619), .b(n_25551), .o(n_25667) );
na02f80 g736820 ( .a(n_43144), .b(n_43130), .o(n_43143) );
no02f80 g756013 ( .a(n_25160), .b(n_25258), .o(n_25735) );
no02f80 g772001 ( .a(FE_OCPN955_n_44460), .b(n_9767), .o(n_9825) );
in01f80 newInst_2069 ( .a(newNet_1124), .o(newNet_2069) );
na02f80 g774763 ( .a(n_6253), .b(n_6230), .o(n_6373) );
no02f80 g755134 ( .a(n_25374), .b(n_24528), .o(n_25554) );
no02f80 g775665 ( .a(n_47000), .b(n_5629), .o(n_5661) );
no02f80 g772924 ( .a(n_7863), .b(n_7900), .o(n_7901) );
in01f80 g738847 ( .a(n_41312), .o(n_41324) );
in01f80 g742761 ( .a(n_37894), .o(n_37406) );
oa22f80 g781201 ( .a(n_164), .b(n_136), .c(n_169), .d(n_137), .o(n_362) );
in01f80 g775281 ( .a(n_5836), .o(n_5837) );
in01f80 FE_OCP_RBC2195_n_2103 ( .a(n_2103), .o(FE_OCP_RBN2195_n_2103) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_6_ ( .ck(newNet_1680), .d(n_21802), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_) );
no02f80 g752204 ( .a(n_28586), .b(n_28585), .o(n_28587) );
na02f80 g775920 ( .a(n_5023), .b(n_4727), .o(n_5240) );
na02f80 g773643 ( .a(n_7306), .b(n_7169), .o(n_7347) );
no02f80 g742103 ( .a(n_37872), .b(n_37882), .o(n_37908) );
in01f80 FE_RC_313_0 ( .a(n_20991), .o(FE_RN_94_0) );
in01f80 newInst_3457 ( .a(newNet_3380), .o(newNet_3457) );
na02f80 g776388 ( .a(n_4593), .b(n_4539), .o(n_4762) );
na02f80 FE_RC_2001_0 ( .a(FE_OCPN1790_n_18119), .b(FE_RN_656_0), .o(FE_RN_657_0) );
no02f80 g769978 ( .a(n_10993), .b(n_10927), .o(n_10994) );
na02f80 g762183 ( .a(n_18162), .b(n_16921), .o(n_18243) );
in01f80 g742556 ( .a(n_37509), .o(n_37510) );
na02f80 g776157 ( .a(n_4851), .b(n_4217), .o(n_4927) );
na02f80 g758952 ( .a(n_22058), .b(n_22057), .o(n_22059) );
na02f80 g759997 ( .a(n_20674), .b(n_20533), .o(n_20710) );
oa12f80 g754835 ( .a(n_25951), .b(n_25977), .c(n_25950), .o(n_26679) );
in01f80 g758716 ( .a(n_21766), .o(n_21767) );
no02f80 g736691 ( .a(n_43435), .b(n_43387), .o(n_43436) );
na02f80 g762208 ( .a(n_18695), .b(n_18816), .o(n_18837) );
in01f80 g781357 ( .a(beta_31), .o(n_29) );
no02f80 g771370 ( .a(n_9567), .b(n_9338), .o(n_9611) );
in01f80 g770542 ( .a(n_10469), .o(n_10470) );
in01f80 g778001 ( .a(n_3172), .o(n_3173) );
no02f80 g740113 ( .a(n_40110), .b(n_40135), .o(n_40249) );
in01f80 g744577 ( .a(n_35393), .o(n_35394) );
oa12f80 g748647 ( .a(n_32645), .b(n_32424), .c(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_33028) );
in01f80 newInst_3256 ( .a(newNet_3255), .o(newNet_3256) );
no02f80 g778055 ( .a(n_2995), .b(n_2953), .o(n_3056) );
na02f80 g751839 ( .a(n_29334), .b(n_29309), .o(n_29769) );
no02f80 g780817 ( .a(n_449), .b(n_420), .o(n_466) );
in01f80 g773412 ( .a(n_7669), .o(n_7670) );
no02f80 g778642 ( .a(n_2293), .b(n_2219), .o(n_2335) );
ao12f80 g745236 ( .a(n_34439), .b(n_34465), .c(n_34438), .o(n_34516) );
in01f80 FE_OCP_RBC2984_n_35539 ( .a(FE_OCP_RBN3697_n_35543), .o(FE_OCP_RBN2984_n_35539) );
na02f80 g758076 ( .a(n_44267), .b(n_20717), .o(n_22267) );
no02f80 g766121 ( .a(n_14628), .b(FE_OCP_RBN3529_n_13765), .o(n_14629) );
in01f80 g772877 ( .a(n_8006), .o(n_8007) );
na02f80 g771281 ( .a(n_9531), .b(n_9586), .o(n_9617) );
no02f80 g776893 ( .a(n_3789), .b(n_3821), .o(n_5629) );
oa22f80 FE_RC_1151_0 ( .a(n_38258), .b(n_38571), .c(n_38570), .d(n_38259), .o(n_38615) );
in01f80 FE_OCPC1485_n_27315 ( .a(n_27315), .o(FE_OCPN1485_n_27315) );
in01f80 g763483 ( .a(n_17734), .o(n_17708) );
no02f80 g778544 ( .a(n_2273), .b(n_2267), .o(n_2332) );
in01f80 newInst_195 ( .a(newNet_159), .o(newNet_195) );
ao12f80 g779109 ( .a(n_1669), .b(n_1964), .c(n_1646), .o(n_2023) );
no02f80 g772734 ( .a(n_8254), .b(n_45827), .o(n_8291) );
in01f80 FE_OCP_RBC3561_n_29857 ( .a(n_29857), .o(FE_OCP_RBN3561_n_29857) );
oa12f80 g783844 ( .a(n_45841), .b(n_39594), .c(n_39579), .o(n_45530) );
na02f80 g743310 ( .a(n_36690), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36756) );
in01f80 FE_OCP_DRV_C3154_n_24425 ( .a(FE_OCP_DRV_N3153_n_24425), .o(FE_OCP_DRV_N3154_n_24425) );
na02f80 g784783 ( .a(n_11089), .b(n_44511), .o(n_47269) );
in01f80 g756792 ( .a(n_23422), .o(n_23423) );
in01f80 g757371 ( .a(n_24142), .o(n_24249) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_17_ ( .ck(newNet_247), .d(n_46180), .o(delay_xor_ln22_unr6_stage3_stallmux_q_17_) );
no02f80 g738339 ( .a(n_41790), .b(n_41813), .o(n_41859) );
in01f80 newInst_1476 ( .a(newNet_1475), .o(newNet_1476) );
in01f80 newInst_2380 ( .a(newNet_722), .o(newNet_2380) );
in01f80 g742755 ( .a(n_37299), .o(n_37317) );
in01f80 g746954 ( .a(n_33032), .o(n_33078) );
no02f80 g756814 ( .a(n_23753), .b(n_23703), .o(n_24171) );
in01f80 g771629 ( .a(n_8817), .o(n_8818) );
oa12f80 g751723 ( .a(n_28312), .b(n_28322), .c(n_28311), .o(n_28349) );
in01f80 g738968 ( .a(n_41211), .o(n_41212) );
in01f80 g741744 ( .a(n_38564), .o(n_38543) );
na02f80 FE_RC_2219_0 ( .a(FE_RN_802_0), .b(n_32750), .o(n_32782) );
no02f80 g741686 ( .a(n_38566), .b(n_38551), .o(n_38591) );
in01f80 FE_OCP_RBC3644_n_44490 ( .a(FE_OCP_RBN3640_n_44490), .o(FE_OCP_RBN3644_n_44490) );
in01f80 FE_OFC777_n_17093 ( .a(n_17093), .o(FE_OFN777_n_17093) );
in01f80 g741663 ( .a(n_38570), .o(n_38571) );
na02f80 g742199 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38209), .o(n_38227) );
na02f80 g752429 ( .a(FE_OCP_RBN3309_n_44722), .b(n_27719), .o(n_27868) );
in01f80 FE_RC_1159_0 ( .a(FE_OCPN1013_n_41478), .o(FE_RN_348_0) );
na02f80 g755691 ( .a(n_25311), .b(n_25368), .o(n_25369) );
ms00f80 delay_sub_ln23_0_unr27_stage9_stallmux_q_reg ( .ck(newNet_1440), .d(FE_OCP_RBN2994_n_35539), .o(delay_sub_ln23_0_unr27_stage10_stallmux_z) );
in01f80 g778372 ( .a(n_2947), .o(n_2791) );
no02f80 g767961 ( .a(n_13032), .b(n_13150), .o(n_13164) );
na02f80 g749351 ( .a(n_30644), .b(n_30281), .o(n_30675) );
na02f80 g758003 ( .a(n_22733), .b(n_22725), .o(n_22852) );
no02f80 g777147 ( .a(n_4818), .b(n_4721), .o(n_4796) );
in01f80 g736624 ( .a(n_43238), .o(n_43239) );
oa12f80 g763705 ( .a(n_17498), .b(n_17497), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n_17537) );
in01f80 g747943 ( .a(n_33191), .o(n_33208) );
no02f80 g752112 ( .a(n_28688), .b(n_28260), .o(n_28749) );
no02f80 g770308 ( .a(n_10520), .b(n_10488), .o(n_10629) );
in01f80 newInst_100 ( .a(newNet_99), .o(newNet_100) );
no02f80 g739478 ( .a(FE_OCPN932_n_40736), .b(n_40523), .o(n_40775) );
na02f80 g751740 ( .a(n_28321), .b(n_28344), .o(n_28514) );
in01f80 newInst_523 ( .a(newNet_522), .o(newNet_523) );
in01f80 g781237 ( .a(n_136), .o(n_137) );
in01f80 FE_OCP_RBC2644_n_34980 ( .a(n_34980), .o(FE_OCP_RBN2644_n_34980) );
in01f80 FE_OCPC1018_n_23078 ( .a(n_23078), .o(FE_OCPN1018_n_23078) );
oa22f80 g763875 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .c(n_17496), .d(FE_OCP_RBN3359_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17526) );
no02f80 g746784 ( .a(n_33855), .b(n_33338), .o(n_33378) );
in01f80 g770486 ( .a(FE_OCP_RBN2874_n_10477), .o(n_11435) );
na02f80 g761277 ( .a(n_19906), .b(n_19931), .o(n_19907) );
na02f80 FE_RC_3752_0 ( .a(FE_RN_1647_0), .b(FE_RN_536_0), .o(n_12137) );
in01f80 g742512 ( .a(n_37606), .o(n_37624) );
na02f80 g773819 ( .a(n_7130), .b(n_5884), .o(n_7207) );
in01f80 FE_OCP_RBC3131_n_43762 ( .a(n_43762), .o(FE_OCP_RBN3131_n_43762) );
no02f80 g739416 ( .a(n_40710), .b(n_40808), .o(n_40876) );
in01f80 g767970 ( .a(n_13198), .o(n_13199) );
na02f80 g745716 ( .a(n_34185), .b(n_44102), .o(n_34221) );
in01f80 g769726 ( .a(n_11394), .o(n_11306) );
in01f80 g780297 ( .a(n_1056), .o(n_1008) );
no02f80 FE_RC_3076_0 ( .a(FE_RN_1353_0), .b(FE_RN_1354_0), .o(FE_RN_1355_0) );
in01f80 FE_RC_2762_0 ( .a(n_8907), .o(FE_RN_1176_0) );
na02f80 g740598 ( .a(n_39592), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39616) );
in01f80 g759930 ( .a(n_21403), .o(n_21404) );
na02f80 g780557 ( .a(n_745), .b(n_748), .o(n_761) );
na02f80 g747129 ( .a(n_32708), .b(n_32775), .o(n_32898) );
na02f80 g755399 ( .a(n_24894), .b(n_24893), .o(n_24961) );
oa12f80 g762627 ( .a(n_17608), .b(n_45529), .c(n_17605), .o(n_18327) );
no02f80 g741014 ( .a(n_39011), .b(n_38987), .o(n_39139) );
in01f80 g762070 ( .a(n_18390), .o(n_18461) );
ao12f80 g784615 ( .a(n_42634), .b(n_42379), .c(n_42587), .o(n_46943) );
no02f80 g755987 ( .a(n_24908), .b(n_24907), .o(n_24909) );
na02f80 g751789 ( .a(n_28271), .b(n_28270), .o(n_28272) );
in01f80 g768062 ( .a(n_12810), .o(n_12776) );
oa12f80 g769888 ( .a(n_10979), .b(n_11003), .c(n_10923), .o(n_11081) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_20_ ( .ck(newNet_2098), .d(n_6248), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_20_) );
in01f80 g757949 ( .a(n_22273), .o(n_22274) );
no02f80 g773529 ( .a(n_7435), .b(n_7271), .o(n_7462) );
in01f80 newInst_3563 ( .a(newNet_1957), .o(newNet_3563) );
na02f80 g737189 ( .a(n_42964), .b(n_42976), .o(n_43003) );
in01f80 g747309 ( .a(n_32729), .o(n_32730) );
in01f80 g752407 ( .a(n_27773), .o(n_27829) );
na02f80 g739059 ( .a(n_41087), .b(n_41086), .o(n_41088) );
no02f80 g768048 ( .a(n_12790), .b(n_12871), .o(n_12918) );
na02f80 g750809 ( .a(n_29037), .b(n_28704), .o(n_29097) );
in01f80 FE_OCP_RBC1362_n_20504 ( .a(n_20504), .o(FE_OCP_RBN1362_n_20504) );
in01f80 g736889 ( .a(n_43591), .o(n_43592) );
in01f80 g777298 ( .a(n_5186), .o(n_5187) );
ms00f80 sin_out_reg_14_ ( .ck(newNet_80), .d(n_43824), .o(sin_out_14) );
in01f80 g755045 ( .a(n_25446), .o(n_25447) );
in01f80 newInst_79 ( .a(newNet_78), .o(newNet_79) );
in01f80 g741490 ( .a(n_38758), .o(n_38759) );
in01f80 newInst_1491 ( .a(newNet_1490), .o(newNet_1491) );
na02f80 g743509 ( .a(n_37634), .b(n_46240), .o(n_37635) );
in01f80 newInst_1975 ( .a(newNet_1974), .o(newNet_1975) );
in01f80 FE_RC_2426_0 ( .a(n_6717), .o(FE_RN_963_0) );
in01f80 g750285 ( .a(n_29755), .o(n_29792) );
oa22f80 g741105 ( .a(FE_OCP_RBN3626_n_38870), .b(FE_OCP_RBN2397_n_38586), .c(FE_OCP_RBN2685_n_38870), .d(n_38608), .o(n_39207) );
in01f80 newInst_2251 ( .a(newNet_2083), .o(newNet_2251) );
in01f80 FE_OCP_RBC3135_n_6567 ( .a(n_6567), .o(FE_OCP_RBN3135_n_6567) );
in01f80 fopt783366 ( .a(n_44955), .o(n_44954) );
ao22s80 FE_RC_1286_0 ( .a(n_38705), .b(FE_OCP_RBN2531_n_38693), .c(n_38693), .d(n_38706), .o(n_38753) );
in01f80 newInst_3373 ( .a(newNet_3372), .o(newNet_3373) );
in01f80 g764247 ( .a(n_16464), .o(n_16465) );
in01f80 g768854 ( .a(n_12058), .o(n_12150) );
na02f80 g752226 ( .a(n_27919), .b(n_27839), .o(n_27920) );
in01f80 FE_OCP_RBC3731_n_31819 ( .a(FE_OCP_RBN3085_n_31819), .o(FE_OCP_RBN3731_n_31819) );
no02f80 g738926 ( .a(n_41172), .b(n_40944), .o(n_41231) );
no02f80 g780477 ( .a(n_845), .b(n_754), .o(n_1098) );
ao12f80 g781199 ( .a(n_93), .b(n_157), .c(n_104), .o(n_172) );
no02f80 g777636 ( .a(n_3474), .b(n_3429), .o(n_3549) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_25_ ( .ck(newNet_1392), .d(n_36700), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_) );
ao12f80 g780737 ( .a(n_560), .b(n_601), .c(n_570), .o(n_605) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_1_ ( .ck(newNet_1749), .d(n_21338), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_) );
na02f80 g751537 ( .a(n_28460), .b(n_28630), .o(n_28734) );
no02f80 g749066 ( .a(n_30888), .b(n_30887), .o(n_30889) );
in01f80 g764412 ( .a(n_16234), .o(n_16228) );
in01f80 g774838 ( .a(n_6362), .o(n_6389) );
no02f80 g765647 ( .a(n_15017), .b(n_15018), .o(n_15038) );
no02f80 g741113 ( .a(n_38995), .b(n_38939), .o(n_38996) );
ao12f80 g767832 ( .a(n_12475), .b(n_12668), .c(n_12507), .o(n_12727) );
oa12f80 g742941 ( .a(n_36996), .b(n_37082), .c(n_36994), .o(n_36997) );
in01f80 newInst_3230 ( .a(newNet_3229), .o(newNet_3230) );
oa12f80 g739774 ( .a(n_40017), .b(n_40406), .c(n_40043), .o(n_40434) );
no02f80 g746379 ( .a(n_33520), .b(n_33519), .o(n_33521) );
ao12f80 g751922 ( .a(n_29024), .b(n_28919), .c(n_28557), .o(n_29536) );
in01f80 g753324 ( .a(n_26991), .o(n_26992) );
na02f80 FE_RC_3614_0 ( .a(FE_RN_1580_0), .b(n_30580), .o(FE_RN_1581_0) );
ao12f80 g782641 ( .a(n_44875), .b(n_37490), .c(n_38268), .o(n_44034) );
in01f80 g770349 ( .a(n_10716), .o(n_10783) );
na02f80 g754905 ( .a(FE_OCP_RBN2593_n_25181), .b(n_24199), .o(n_25275) );
ao12f80 g765240 ( .a(n_14854), .b(n_14944), .c(n_14906), .o(n_15026) );
in01f80 g743897 ( .a(n_46250), .o(n_36980) );
ao12f80 g747706 ( .a(n_33571), .b(n_33684), .c(n_33683), .o(n_33703) );
no02f80 g753262 ( .a(n_27167), .b(n_27170), .o(n_27172) );
no02f80 g759756 ( .a(n_20271), .b(n_20236), .o(n_20298) );
in01f80 g766583 ( .a(FE_OCP_RBN2436_n_14072), .o(n_15299) );
ao22s80 FE_RC_1174_0 ( .a(FE_OCP_RBN2290_n_2438), .b(n_3080), .c(FE_OCP_RBN2295_n_2438), .d(n_3597), .o(n_3116) );
in01f80 FE_OCP_RBC2682_n_35139 ( .a(n_35139), .o(FE_OCP_RBN2682_n_35139) );
in01f80 g751452 ( .a(n_28739), .o(n_28740) );
no02f80 g757998 ( .a(n_22786), .b(n_22785), .o(n_22787) );
na02f80 g762277 ( .a(n_18535), .b(n_18659), .o(n_19228) );
in01f80 g741698 ( .a(n_38519), .o(n_38520) );
no02f80 g773671 ( .a(n_7303), .b(n_7302), .o(n_7304) );
ao12f80 g738283 ( .a(n_41843), .b(n_41842), .c(n_41841), .o(n_42232) );
in01f80 g751031 ( .a(n_29856), .o(n_30182) );
in01f80 newInst_1371 ( .a(newNet_1370), .o(newNet_1371) );
no02f80 g771454 ( .a(n_8977), .b(n_8976), .o(n_9113) );
no02f80 g763199 ( .a(n_17714), .b(n_17305), .o(n_17819) );
na02f80 g740421 ( .a(FE_OCP_RBN3022_n_39942), .b(FE_OCP_RBN2864_n_39523), .o(n_40170) );
in01f80 newInst_2521 ( .a(newNet_2520), .o(newNet_2521) );
in01f80 g773533 ( .a(n_7488), .o(n_7489) );
na02f80 g778041 ( .a(n_3062), .b(n_3109), .o(n_3130) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_16_ ( .ck(newNet_2669), .d(n_22425), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_16_) );
in01f80 g738885 ( .a(n_41263), .o(n_41228) );
no02f80 g775506 ( .a(n_5486), .b(n_5440), .o(n_5441) );
na02f80 g766917 ( .a(n_13967), .b(n_13966), .o(n_14110) );
in01f80 FE_OCP_RBC3662_n_20750 ( .a(n_20750), .o(FE_OCP_RBN3662_n_20750) );
no02f80 g747816 ( .a(n_33238), .b(n_33256), .o(n_33257) );
in01f80 g764320 ( .a(n_16798), .o(n_16770) );
in01f80 newInst_404 ( .a(newNet_403), .o(newNet_404) );
in01f80 newInst_966 ( .a(newNet_965), .o(newNet_966) );
na02f80 g762970 ( .a(n_17739), .b(n_17791), .o(n_17838) );
na02f80 g768643 ( .a(n_12202), .b(n_12201), .o(n_12203) );
oa12f80 g784658 ( .a(n_10900), .b(n_10813), .c(n_10684), .o(n_46988) );
na02f80 g766434 ( .a(n_14101), .b(n_14029), .o(n_14125) );
na02f80 g766025 ( .a(n_14642), .b(n_14601), .o(n_14666) );
no02f80 g752334 ( .a(n_44761), .b(delay_xor_ln22_unr18_stage7_stallmux_q_3_), .o(n_27918) );
no02f80 FE_RC_3295_0 ( .a(FE_RN_1448_0), .b(FE_RN_1449_0), .o(FE_RN_1450_0) );
no02f80 g750182 ( .a(n_29859), .b(n_29787), .o(n_29930) );
no02f80 g777988 ( .a(n_2741), .b(n_47023), .o(n_3037) );
oa12f80 g762672 ( .a(n_18212), .b(n_18237), .c(n_18211), .o(n_18574) );
in01f80 g741620 ( .a(n_38639), .o(n_38640) );
na02f80 g748978 ( .a(n_31127), .b(n_27536), .o(n_31130) );
in01f80 newInst_55 ( .a(newNet_54), .o(newNet_55) );
na02f80 g780590 ( .a(n_890), .b(n_550), .o(n_1006) );
na02f80 g741750 ( .a(n_38474), .b(n_38135), .o(n_38475) );
no02f80 g777788 ( .a(n_3406), .b(n_3556), .o(n_3444) );
in01f80 g762715 ( .a(n_17812), .o(n_17809) );
in01f80 g776451 ( .a(n_4649), .o(n_4650) );
oa12f80 g744589 ( .a(n_36171), .b(n_36577), .c(n_36080), .o(n_36644) );
no02f80 g741992 ( .a(n_38378), .b(n_38329), .o(n_38454) );
in01f80 g771810 ( .a(n_9065), .o(n_9066) );
in01f80 newInst_1584 ( .a(newNet_1069), .o(newNet_1584) );
in01f80 newInst_1755 ( .a(newNet_1754), .o(newNet_1755) );
no02f80 g776371 ( .a(n_47007), .b(n_4662), .o(n_4766) );
no02f80 g741834 ( .a(n_38288), .b(n_38038), .o(n_38321) );
na02f80 g769080 ( .a(n_11715), .b(n_11459), .o(n_11754) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_14_ ( .ck(newNet_1424), .d(n_36527), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_14_) );
ao22s80 g784429 ( .a(n_36744), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .c(n_46197), .d(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n_46241) );
na02f80 g770675 ( .a(n_10191), .b(n_10242), .o(n_10310) );
in01f80 g777855 ( .a(n_3222), .o(n_3238) );
in01f80 g775972 ( .a(n_5171), .o(n_5172) );
in01f80 g753589 ( .a(n_26776), .o(n_26777) );
na02f80 g780187 ( .a(n_1077), .b(n_1159), .o(n_1078) );
in01f80 g767333 ( .a(n_13388), .o(n_13429) );
na02f80 g771539 ( .a(n_9781), .b(n_9605), .o(n_9444) );
na02f80 g744933 ( .a(n_34836), .b(n_30588), .o(n_34864) );
na02f80 g771150 ( .a(n_9458), .b(n_9424), .o(n_9575) );
oa12f80 g738439 ( .a(n_41680), .b(FE_OCPN953_n_41540), .c(n_41590), .o(n_41904) );
no02f80 g745161 ( .a(n_34820), .b(n_34461), .o(n_34767) );
na02f80 g771959 ( .a(n_44463), .b(n_9587), .o(n_9735) );
ao12f80 g759194 ( .a(n_21125), .b(n_21044), .c(n_21074), .o(n_21353) );
na02f80 FE_RC_3703_0 ( .a(FE_RN_1630_0), .b(n_3493), .o(n_47017) );
in01f80 g763075 ( .a(n_17485), .o(n_17486) );
no02f80 g784150 ( .a(n_2168), .b(n_45900), .o(n_45903) );
in01f80 FE_OCP_RBC3492_n_29553 ( .a(n_29553), .o(FE_OCP_RBN3492_n_29553) );
in01f80 fopt783522 ( .a(n_27805), .o(n_45132) );
na02f80 g740898 ( .a(n_44311), .b(n_39360), .o(n_39396) );
no02f80 g775681 ( .a(n_5306), .b(n_5256), .o(n_5458) );
na02f80 g752994 ( .a(n_27263), .b(n_27287), .o(n_27352) );
oa12f80 g756619 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_25_), .c(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23972) );
na02f80 FE_RC_4049_0 ( .a(FE_RN_1758_0), .b(FE_RN_1759_0), .o(FE_RN_1760_0) );
in01f80 g741244 ( .a(n_38984), .o(n_39030) );
ao12f80 g756222 ( .a(n_24741), .b(n_24740), .c(n_24739), .o(n_25138) );
in01f80 newInst_2450 ( .a(newNet_1013), .o(newNet_2450) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_15_ ( .ck(newNet_254), .d(n_46154), .o(delay_xor_ln22_unr6_stage3_stallmux_q_15_) );
ao22s80 g739548 ( .a(n_44028), .b(n_40629), .c(n_40639), .d(FE_OCP_RBN2132_n_40629), .o(n_40668) );
no02f80 g755305 ( .a(n_25470), .b(n_25110), .o(n_25528) );
na02f80 g770407 ( .a(n_10514), .b(n_44054), .o(n_10587) );
in01f80 newInst_3602 ( .a(newNet_50), .o(newNet_3602) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_22_ ( .ck(newNet_1845), .d(n_16927), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_) );
no02f80 g740168 ( .a(n_39816), .b(n_39978), .o(n_40001) );
no02f80 g738752 ( .a(FE_OCPN1013_n_41478), .b(n_41328), .o(n_41788) );
oa22f80 g751397 ( .a(n_28441), .b(n_28329), .c(n_28478), .d(n_28330), .o(n_29715) );
na02f80 g755882 ( .a(n_25089), .b(n_24299), .o(n_25005) );
in01f80 g767240 ( .a(n_13554), .o(n_13555) );
na02f80 g758184 ( .a(n_44277), .b(n_21076), .o(n_22231) );
in01f80 g779066 ( .a(n_2288), .o(n_2794) );
in01f80 newInst_2632 ( .a(newNet_2631), .o(newNet_2632) );
in01f80 g759476 ( .a(n_20735), .o(n_20736) );
in01f80 FE_OCP_RBC2911_n_30908 ( .a(n_30908), .o(FE_OCP_RBN2911_n_30908) );
in01f80 g757400 ( .a(n_22972), .o(n_23109) );
in01f80 g779042 ( .a(n_2074), .o(n_2075) );
no02f80 g761546 ( .a(n_18999), .b(n_18998), .o(n_19000) );
in01f80 g769826 ( .a(n_11235), .o(n_11284) );
in01f80 FE_OCP_RBC2350_n_38515 ( .a(n_38515), .o(FE_OCP_RBN2350_n_38515) );
in01f80 g755979 ( .a(FE_OFN788_n_25834), .o(n_29379) );
in01f80 g743479 ( .a(n_36567), .o(n_36551) );
in01f80 g762684 ( .a(n_17851), .o(n_17930) );
in01f80 g768092 ( .a(n_13210), .o(n_13161) );
no02f80 g776310 ( .a(n_4681), .b(n_4245), .o(n_4798) );
in01f80 g775151 ( .a(n_6034), .o(n_6035) );
na02f80 g750638 ( .a(n_29353), .b(n_28849), .o(n_29330) );
no02f80 g756540 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_27_), .o(n_23854) );
in01f80 FE_OCP_RBC2919_n_16084 ( .a(n_16084), .o(FE_OCP_RBN2919_n_16084) );
na02f80 g749449 ( .a(n_30464), .b(n_27014), .o(n_30515) );
na02f80 g751580 ( .a(n_28817), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n_28887) );
na02f80 g745020 ( .a(n_34947), .b(n_34894), .o(n_34948) );
in01f80 newInst_3225 ( .a(newNet_1072), .o(newNet_3225) );
in01f80 g777029 ( .a(n_4008), .o(n_4118) );
oa22f80 FE_RC_386_0 ( .a(n_1167), .b(FE_OCPN874_n_44672), .c(n_1154), .d(n_44637), .o(n_1314) );
no02f80 g751050 ( .a(n_30094), .b(n_30089), .o(n_30892) );
na02f80 g761651 ( .a(n_18682), .b(FE_OFN778_n_17093), .o(n_18721) );
na02f80 g761770 ( .a(n_18678), .b(n_18646), .o(n_18684) );
in01f80 g760553 ( .a(n_19942), .o(n_19943) );
in01f80 g738775 ( .a(n_41435), .o(n_41483) );
no02f80 g760880 ( .a(n_20017), .b(n_19732), .o(n_20056) );
na02f80 g776642 ( .a(n_4499), .b(n_4498), .o(n_4500) );
no02f80 g762965 ( .a(n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_9_), .o(n_17745) );
no02f80 g781112 ( .a(n_231), .b(n_99), .o(n_244) );
na02f80 g780215 ( .a(n_837), .b(n_812), .o(n_813) );
in01f80 g767517 ( .a(n_13225), .o(n_13226) );
na02f80 g743961 ( .a(n_35747), .b(n_35831), .o(n_35828) );
in01f80 g772336 ( .a(n_8688), .o(n_8689) );
oa22f80 FE_RC_1576_0 ( .a(n_13755), .b(n_13659), .c(n_13673), .d(n_13813), .o(n_13890) );
in01f80 g754388 ( .a(n_25783), .o(n_25813) );
in01f80 g760952 ( .a(n_19450), .o(n_19451) );
ao12f80 g762706 ( .a(n_17967), .b(FE_OCP_RBN2140_FE_OCPN861_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_13_), .o(n_17915) );
oa12f80 g739166 ( .a(n_40848), .b(n_40938), .c(n_40753), .o(n_40992) );
in01f80 newInst_1342 ( .a(newNet_1341), .o(newNet_1342) );
na02f80 g778225 ( .a(n_2619), .b(n_2326), .o(n_3208) );
no02f80 g749194 ( .a(n_30829), .b(FE_OCPN1486_n_27315), .o(n_30887) );
no02f80 FE_RC_3549_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .b(n_32525), .o(FE_RN_1539_0) );
na02f80 g743842 ( .a(n_35832), .b(n_35707), .o(n_35833) );
in01f80 g776525 ( .a(n_4177), .o(n_4178) );
na02f80 g743645 ( .a(n_44835), .b(n_36099), .o(n_36441) );
no02f80 g766368 ( .a(n_14099), .b(FE_OCP_RBN2249_n_13017), .o(n_14135) );
in01f80 FE_OCP_RBC2223_n_12902 ( .a(n_12902), .o(FE_OCP_RBN2223_n_12902) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_10_ ( .ck(newNet_2498), .d(n_31878), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_) );
in01f80 newInst_2316 ( .a(newNet_2210), .o(newNet_2316) );
in01f80 g748669 ( .a(n_31421), .o(n_31437) );
oa12f80 g779460 ( .a(n_2113), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_28_), .o(n_2683) );
no02f80 g775277 ( .a(n_5816), .b(n_5808), .o(n_5867) );
na02f80 g745774 ( .a(n_34242), .b(n_34258), .o(n_34304) );
ao12f80 g757942 ( .a(n_22027), .b(n_22085), .c(n_21970), .o(n_22172) );
in01f80 g769756 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_15_), .o(n_11298) );
in01f80 g758839 ( .a(n_21556), .o(n_21510) );
no02f80 g740626 ( .a(n_39628), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39638) );
in01f80 newInst_1176 ( .a(newNet_1175), .o(newNet_1176) );
ao22s80 FE_RC_807_0 ( .a(n_7661), .b(n_8704), .c(n_7660), .d(n_8703), .o(n_8842) );
na02f80 g758264 ( .a(FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .o(n_22645) );
na02f80 g756470 ( .a(n_23584), .b(n_23663), .o(n_23687) );
no02f80 g754972 ( .a(n_25152), .b(n_25151), .o(n_25153) );
in01f80 fopt783496 ( .a(n_45065), .o(n_45066) );
oa22f80 g773602 ( .a(n_7351), .b(n_6921), .c(n_7352), .d(n_6920), .o(n_7853) );
in01f80 g747647 ( .a(n_32384), .o(n_32358) );
in01f80 g769577 ( .a(n_11377), .o(n_11378) );
na02f80 g775722 ( .a(n_5335), .b(n_4009), .o(n_5357) );
in01f80 g742577 ( .a(n_37969), .o(n_38273) );
in01f80 g780602 ( .a(n_682), .o(n_690) );
ao12f80 g760169 ( .a(n_20900), .b(n_20899), .c(n_20898), .o(n_21562) );
na03f80 FE_RC_1127_0 ( .a(n_40915), .b(n_40732), .c(n_40743), .o(n_40946) );
no02f80 g755525 ( .a(n_24647), .b(n_23996), .o(n_24723) );
no02f80 g747622 ( .a(n_33394), .b(n_33393), .o(n_33395) );
oa12f80 g762425 ( .a(n_18352), .b(n_18351), .c(n_18350), .o(n_18660) );
in01f80 g741866 ( .a(n_38288), .o(n_38368) );
oa12f80 g754338 ( .a(n_26613), .b(FE_OCP_RBN3704_n_26231), .c(n_26855), .o(n_26944) );
oa12f80 g758668 ( .a(n_21782), .b(n_22363), .c(n_21779), .o(n_22431) );
in01f80 g780303 ( .a(n_1050), .o(n_1092) );
no02f80 g747374 ( .a(FE_OCP_RBN3333_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_4_), .o(n_32600) );
ao12f80 g743069 ( .a(n_37091), .b(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_13_), .o(n_37441) );
ao22s80 g775356 ( .a(FE_OCP_RBN2946_n_5428), .b(n_5093), .c(n_5428), .d(n_5094), .o(n_5555) );
no02f80 g764427 ( .a(n_16053), .b(n_14419), .o(n_16094) );
in01f80 newInst_389 ( .a(newNet_33), .o(newNet_389) );
na02f80 g738495 ( .a(n_41660), .b(n_41330), .o(n_41691) );
in01f80 newInst_3351 ( .a(newNet_2130), .o(newNet_3351) );
no02f80 g736803 ( .a(n_43391), .b(n_43390), .o(n_43425) );
in01f80 g770936 ( .a(n_10006), .o(n_10007) );
na02f80 g748809 ( .a(n_32454), .b(n_32487), .o(n_33084) );
oa22f80 g756951 ( .a(n_24059), .b(n_23897), .c(n_24188), .d(n_23341), .o(n_24300) );
no02f80 g771015 ( .a(n_9726), .b(n_9672), .o(n_9749) );
in01f80 newInst_2501 ( .a(newNet_2500), .o(newNet_2501) );
na02f80 g737681 ( .a(n_42392), .b(n_42483), .o(n_42485) );
in01f80 g749667 ( .a(n_30080), .o(n_30154) );
no02f80 g763905 ( .a(n_17256), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n_17363) );
in01f80 g774237 ( .a(n_6594), .o(n_6595) );
na02f80 FE_RC_2162_0 ( .a(FE_RN_765_0), .b(FE_RN_766_0), .o(n_15652) );
na02f80 g759408 ( .a(n_20823), .b(n_20732), .o(n_20854) );
oa22f80 g751527 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_17_), .c(n_28460), .d(n_27712), .o(n_29014) );
in01f80 g740250 ( .a(n_40365), .o(n_40366) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_28_ ( .ck(newNet_2456), .d(FE_OCP_RBN3142_n_32395), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_) );
in01f80 FE_OCP_RBC2388_n_13860 ( .a(n_13860), .o(FE_OCP_RBN2388_n_13860) );
no02f80 g774361 ( .a(n_6528), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n_6671) );
oa12f80 g766983 ( .a(n_13799), .b(n_13798), .c(n_13797), .o(n_14304) );
oa22f80 g737871 ( .a(n_42270), .b(n_41949), .c(n_42547), .d(n_41923), .o(n_42574) );
in01f80 g756757 ( .a(n_25092), .o(n_24236) );
na02f80 g764305 ( .a(n_16401), .b(n_16400), .o(n_16432) );
in01f80 newInst_1670 ( .a(newNet_1669), .o(newNet_1670) );
ao12f80 g747116 ( .a(FE_RN_193_0), .b(n_32721), .c(FE_OCPN1236_n_32791), .o(n_32761) );
in01f80 g765061 ( .a(FE_OCP_RBN3659_n_15314), .o(n_15351) );
na02f80 g740377 ( .a(n_39787), .b(n_39853), .o(n_39915) );
na02f80 g778412 ( .a(n_2470), .b(n_2444), .o(n_2607) );
na02f80 g759944 ( .a(FE_OCP_RBN3678_n_21051), .b(n_21625), .o(n_21825) );
no02f80 g766732 ( .a(n_13751), .b(FE_OCP_RBN2246_n_13017), .o(n_13775) );
na02f80 g737577 ( .a(n_42446), .b(n_42445), .o(n_42447) );
in01f80 newInst_2612 ( .a(newNet_2611), .o(newNet_2612) );
ao12f80 g742865 ( .a(n_36937), .b(n_37058), .c(n_36924), .o(n_37200) );
na02f80 g776111 ( .a(n_5048), .b(n_4467), .o(n_4940) );
na02f80 g777068 ( .a(n_3662), .b(n_3734), .o(n_3735) );
no02f80 FE_RC_2400_0 ( .a(FE_RN_945_0), .b(n_42843), .o(FE_RN_946_0) );
in01f80 g741081 ( .a(n_39187), .o(n_39188) );
no02f80 g748395 ( .a(FE_OCP_RBN3712_n_31466), .b(n_30492), .o(n_31554) );
oa12f80 g750489 ( .a(n_29560), .b(n_29559), .c(n_29558), .o(n_31012) );
na02f80 g738592 ( .a(n_41419), .b(n_41447), .o(n_41448) );
no02f80 g761699 ( .a(n_18715), .b(n_18600), .o(n_18794) );
in01f80 FE_RC_2190_0 ( .a(n_15009), .o(FE_RN_784_0) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_4_ ( .ck(newNet_909), .d(n_27749), .o(n_45202) );
na02f80 g752625 ( .a(n_27535), .b(n_27264), .o(n_27573) );
na02f80 g736659 ( .a(n_43405), .b(n_43393), .o(n_43564) );
ao12f80 g768135 ( .a(n_12386), .b(n_12591), .c(n_12424), .o(n_12629) );
na02f80 g768505 ( .a(n_12343), .b(n_10715), .o(n_12424) );
na02f80 FE_RC_191_0 ( .a(FE_OCP_RBN3483_n_13667), .b(FE_RN_64_0), .o(FE_RN_65_0) );
na02f80 g759493 ( .a(n_20851), .b(n_20822), .o(n_20935) );
oa12f80 g742887 ( .a(n_46254), .b(n_37073), .c(delay_add_ln22_unr23_stage9_stallmux_q_15_), .o(n_37129) );
no02f80 g750864 ( .a(n_30168), .b(n_30040), .o(n_30335) );
oa12f80 g753538 ( .a(n_26675), .b(n_26674), .c(n_26705), .o(n_26731) );
in01f80 g779780 ( .a(n_1415), .o(n_1480) );
in01f80 FE_OCPC1508_n_23414 ( .a(FE_OCPN1507_n_23414), .o(FE_OCPN1508_n_23414) );
ao12f80 g746718 ( .a(n_34232), .b(n_34231), .c(n_34230), .o(n_34735) );
na02f80 g771682 ( .a(n_9240), .b(n_44575), .o(n_9378) );
in01f80 newInst_1055 ( .a(newNet_1054), .o(newNet_1055) );
no03m80 g767911 ( .a(n_12992), .b(n_13080), .c(n_13079), .o(n_13252) );
in01f80 newInst_44 ( .a(newNet_43), .o(newNet_44) );
no02f80 g780411 ( .a(n_796), .b(n_788), .o(n_1180) );
in01f80 FE_OFC220_n_35655 ( .a(n_35655), .o(FE_OFN220_n_35655) );
oa22f80 FE_RC_186_0 ( .a(n_11734), .b(n_11788), .c(n_11735), .d(n_11789), .o(n_11941) );
no02f80 g741283 ( .a(n_44921), .b(n_38572), .o(n_38942) );
in01f80 g781265 ( .a(n_96), .o(n_97) );
na02f80 FE_RC_3171_0 ( .a(FE_RN_1403_0), .b(FE_RN_1404_0), .o(FE_RN_1405_0) );
in01f80 g742612 ( .a(n_46952), .o(n_37492) );
in01f80 g760997 ( .a(n_19445), .o(n_19446) );
in01f80 g758573 ( .a(n_21938), .o(n_21939) );
in01f80 g747852 ( .a(n_33762), .o(n_33239) );
in01f80 FE_RC_4008_0 ( .a(FE_OCPN1441_n_45060), .o(FE_RN_1740_0) );
na02f80 g754322 ( .a(n_45533), .b(n_25831), .o(n_25832) );
na02f80 g747334 ( .a(n_32810), .b(n_32684), .o(n_32686) );
na02f80 FE_RC_1897_0 ( .a(n_24262), .b(n_24222), .o(FE_RN_593_0) );
in01f80 g751762 ( .a(FE_OCPN989_n_28353), .o(n_28354) );
na02f80 g753290 ( .a(n_27287), .b(n_26048), .o(n_27463) );
oa12f80 g769013 ( .a(n_11538), .b(n_11473), .c(n_11477), .o(n_11603) );
in01f80 newInst_958 ( .a(newNet_957), .o(newNet_958) );
in01f80 g748510 ( .a(n_31447), .o(n_31471) );
oa22f80 g747357 ( .a(n_32525), .b(n_30905), .c(n_32432), .d(delay_sub_ln21_0_unr20_stage8_stallmux_q_0_), .o(n_33768) );
no02f80 g739976 ( .a(FE_OCP_RBN3717_n_39913), .b(n_40155), .o(n_40227) );
na02f80 g774971 ( .a(n_6163), .b(n_6127), .o(n_6237) );
na02f80 g754096 ( .a(n_26097), .b(n_23339), .o(n_26120) );
oa12f80 g751378 ( .a(n_29171), .b(n_29363), .c(n_29200), .o(n_29410) );
no02f80 g755471 ( .a(n_24579), .b(n_24626), .o(n_24656) );
in01f80 FE_OCP_RBC1094_n_45224 ( .a(n_45224), .o(FE_OCP_RBN1094_n_45224) );
in01f80 g772349 ( .a(n_8546), .o(n_8547) );
no02f80 g753105 ( .a(n_27295), .b(n_27601), .o(n_27396) );
in01f80 FE_OCP_RBC3483_n_13667 ( .a(FE_OCP_RBN3482_n_13667), .o(FE_OCP_RBN3483_n_13667) );
in01f80 g769604 ( .a(n_11415), .o(n_11416) );
no02f80 g770910 ( .a(n_10166), .b(n_10130), .o(n_10424) );
no02f80 g755074 ( .a(n_25554), .b(n_25532), .o(n_25615) );
in01f80 newInst_822 ( .a(newNet_716), .o(newNet_822) );
in01f80 FE_OCP_RBC2894_n_39575 ( .a(n_39575), .o(FE_OCP_RBN2894_n_39575) );
oa12f80 g753466 ( .a(n_26696), .b(n_26767), .c(n_26766), .o(n_26768) );
no02f80 g761513 ( .a(n_18921), .b(n_18942), .o(n_19054) );
no02f80 g769300 ( .a(n_11418), .b(n_11429), .o(n_11568) );
in01f80 newInst_3010 ( .a(newNet_3009), .o(newNet_3010) );
in01f80 newInst_211 ( .a(newNet_210), .o(newNet_211) );
in01f80 g760277 ( .a(n_20387), .o(n_20428) );
oa12f80 g768295 ( .a(n_12389), .b(n_44426), .c(n_12346), .o(n_12591) );
ao12f80 g778490 ( .a(n_3229), .b(n_2549), .c(FE_OCP_RBN2294_n_2438), .o(n_2735) );
in01f80 g775161 ( .a(n_6025), .o(n_6026) );
na02f80 g765192 ( .a(n_15881), .b(n_15749), .o(n_15882) );
na02f80 g780627 ( .a(n_890), .b(n_808), .o(n_1051) );
no02f80 g748918 ( .a(n_32375), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32390) );
oa12f80 g776527 ( .a(n_3873), .b(n_3992), .c(n_3983), .o(n_4154) );
na02f80 g768362 ( .a(n_12445), .b(n_12320), .o(n_12490) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_15_ ( .ck(newNet_1337), .d(n_1219), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_22_ ( .ck(newNet_1314), .d(n_1257), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_) );
na02f80 g751816 ( .a(n_28283), .b(n_28267), .o(n_28343) );
in01f80 newInst_217 ( .a(newNet_54), .o(newNet_217) );
oa22f80 g779073 ( .a(n_2076), .b(n_1830), .c(n_2065), .d(n_1829), .o(n_2127) );
ao12f80 g779470 ( .a(n_1770), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .o(n_1804) );
no02f80 g770835 ( .a(n_9978), .b(n_10008), .o(n_10089) );
no02f80 FE_RC_184_0 ( .a(FE_RN_60_0), .b(FE_RN_61_0), .o(FE_RN_62_0) );
no02f80 g766872 ( .a(n_14347), .b(n_14350), .o(n_14348) );
na02f80 g755361 ( .a(n_24912), .b(n_24959), .o(n_24960) );
no02f80 g779552 ( .a(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .o(n_1544) );
no02f80 g773436 ( .a(n_7551), .b(n_7550), .o(n_7552) );
in01f80 g771492 ( .a(n_9093), .o(n_9137) );
in01f80 g755787 ( .a(n_24346), .o(n_24402) );
in01f80 FE_OCPC3773_n_15371 ( .a(FE_OCPN3772_n_15371), .o(FE_OCPN3773_n_15371) );
oa12f80 g738603 ( .a(n_41686), .b(n_41713), .c(n_41326), .o(n_42061) );
na02f80 g771502 ( .a(n_9484), .b(n_9471), .o(n_9641) );
na02f80 g742637 ( .a(n_37522), .b(n_37521), .o(n_37523) );
na02f80 g765078 ( .a(n_15345), .b(n_15306), .o(n_15422) );
no02f80 g750055 ( .a(n_29896), .b(n_29081), .o(n_30018) );
no02f80 g742155 ( .a(n_38157), .b(n_38130), .o(n_38197) );
in01f80 g772393 ( .a(n_8491), .o(n_8492) );
na02f80 g770727 ( .a(n_10387), .b(n_10167), .o(n_10388) );
na02f80 g777279 ( .a(n_3912), .b(n_3911), .o(n_4090) );
in01f80 g760618 ( .a(n_19880), .o(n_19881) );
na02f80 g770174 ( .a(n_10759), .b(n_10735), .o(n_10809) );
no02f80 g755260 ( .a(n_25011), .b(n_24799), .o(n_25040) );
no02f80 g769595 ( .a(FE_OCP_RBN3063_n_11325), .b(n_11351), .o(n_11388) );
in01f80 newInst_1845 ( .a(newNet_1844), .o(newNet_1845) );
na02f80 g771213 ( .a(n_9881), .b(n_9880), .o(n_9882) );
no02f80 g737014 ( .a(n_43230), .b(n_43418), .o(n_43451) );
in01f80 g740903 ( .a(n_39288), .o(n_39289) );
in01f80 g779807 ( .a(n_1539), .o(n_1540) );
in01f80 g750502 ( .a(n_29585), .o(n_29586) );
na02f80 g781205 ( .a(n_95), .b(n_155), .o(n_156) );
no02f80 g755944 ( .a(n_24186), .b(n_23824), .o(n_24274) );
oa12f80 g740763 ( .a(n_39183), .b(n_39493), .c(n_39206), .o(n_39516) );
no02f80 g778204 ( .a(n_2795), .b(n_2794), .o(n_2830) );
no02f80 g744721 ( .a(n_35172), .b(n_35168), .o(n_35230) );
no02f80 g740151 ( .a(n_39781), .b(n_39841), .o(n_39982) );
no02f80 g780830 ( .a(n_478), .b(n_467), .o(n_484) );
na02f80 g770242 ( .a(n_10801), .b(FE_OCP_RBN3003_n_10805), .o(n_10925) );
no02f80 g743102 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_), .o(n_37109) );
no02f80 FE_RC_2812_0 ( .a(n_9726), .b(n_9723), .o(FE_RN_1204_0) );
no02f80 g752907 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n_27991) );
in01f80 newInst_3057 ( .a(newNet_877), .o(newNet_3057) );
na02f80 g780165 ( .a(n_1075), .b(n_882), .o(n_948) );
in01f80 FE_RC_376_0 ( .a(n_12457), .o(FE_RN_112_0) );
ao12f80 g737500 ( .a(n_42497), .b(n_42498), .c(n_42225), .o(n_42555) );
na02f80 g780878 ( .a(n_521), .b(n_424), .o(n_567) );
no02f80 g761356 ( .a(n_19054), .b(FE_OCP_DRV_N1550_n_19053), .o(n_19130) );
na02f80 g746726 ( .a(n_34212), .b(n_33740), .o(n_34233) );
in01f80 g757128 ( .a(n_24059), .o(n_27796) );
no02f80 g739620 ( .a(FE_OCP_RBN3339_n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n_40655) );
in01f80 g740058 ( .a(n_40145), .o(n_40146) );
na02f80 g755108 ( .a(n_24161), .b(n_25178), .o(n_25205) );
na02f80 g766208 ( .a(n_14472), .b(n_14473), .o(n_14505) );
na02f80 g780452 ( .a(n_855), .b(n_580), .o(n_881) );
in01f80 newInst_149 ( .a(newNet_148), .o(newNet_149) );
in01f80 FE_OCPC1527_n_26296 ( .a(n_26296), .o(FE_OCPN1527_n_26296) );
in01f80 FE_OCP_RBC2250_n_13017 ( .a(FE_OCP_RBN2248_n_13017), .o(FE_OCP_RBN2250_n_13017) );
in01f80 g765163 ( .a(n_15972), .o(n_15973) );
na02f80 g758225 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_), .o(n_22732) );
no02f80 FE_RC_2487_0 ( .a(FE_RN_1002_0), .b(FE_RN_1005_0), .o(n_10551) );
in01f80 g744511 ( .a(n_35444), .o(n_35425) );
no02f80 g754413 ( .a(n_25676), .b(n_25379), .o(n_25706) );
ao22s80 g751508 ( .a(FE_OCP_RBN3402_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_23_), .c(n_28597), .d(n_28606), .o(n_28699) );
no02f80 g778998 ( .a(n_2077), .b(n_1629), .o(n_2101) );
na02f80 g751466 ( .a(n_28547), .b(n_28466), .o(n_28496) );
in01f80 newInst_545 ( .a(newNet_194), .o(newNet_545) );
in01f80 g777160 ( .a(n_5328), .o(n_5260) );
na02f80 g774587 ( .a(n_6363), .b(n_5648), .o(n_6397) );
no02f80 FE_RC_2631_0 ( .a(n_12350), .b(delay_add_ln22_unr8_stage4_stallmux_q_10_), .o(FE_RN_1095_0) );
in01f80 newInst_225 ( .a(newNet_224), .o(newNet_225) );
no02f80 g753404 ( .a(n_27010), .b(n_27009), .o(n_27024) );
oa12f80 g737225 ( .a(n_42363), .b(n_42888), .c(n_42280), .o(n_42933) );
in01f80 newInst_1298 ( .a(newNet_1297), .o(newNet_1298) );
in01f80 g762949 ( .a(n_17725), .o(n_17674) );
in01f80 g770822 ( .a(n_10017), .o(n_10059) );
in01f80 newInst_3280 ( .a(newNet_828), .o(newNet_3280) );
no02f80 g772726 ( .a(n_8147), .b(n_7886), .o(n_8148) );
na02f80 g763687 ( .a(n_16750), .b(n_16734), .o(n_16827) );
in01f80 g756487 ( .a(n_23879), .o(n_23880) );
na02f80 g749648 ( .a(n_30283), .b(n_30265), .o(n_30266) );
no02f80 g750697 ( .a(n_29263), .b(n_28740), .o(n_29301) );
in01f80 g763235 ( .a(n_17279), .o(n_17280) );
in01f80 g757024 ( .a(n_23905), .o(n_23862) );
ao12f80 g774168 ( .a(n_7099), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .o(n_7245) );
ao12f80 g741216 ( .a(n_38925), .b(FE_OCP_RBN3581_n_44944), .c(n_38892), .o(n_39228) );
no02f80 g780632 ( .a(n_779), .b(n_828), .o(n_887) );
no02f80 g771120 ( .a(n_9553), .b(n_9552), .o(n_9554) );
in01f80 g738399 ( .a(n_41703), .o(n_41704) );
na02f80 g749320 ( .a(n_30611), .b(n_30585), .o(n_30652) );
no02f80 g758139 ( .a(n_22415), .b(n_22291), .o(n_22416) );
oa12f80 g736597 ( .a(n_306), .b(n_43191), .c(FE_OFN5_n_43918), .o(n_43337) );
in01f80 g780568 ( .a(n_742), .o(n_743) );
no02f80 g766606 ( .a(n_14435), .b(n_14007), .o(n_14457) );
na02f80 g755594 ( .a(n_45633), .b(n_24555), .o(n_24639) );
in01f80 g773126 ( .a(n_7741), .o(n_7782) );
na02f80 g742113 ( .a(n_37928), .b(n_37965), .o(n_38000) );
oa22f80 g784560 ( .a(FE_OFN800_n_46285), .b(n_10705), .c(FE_OCP_RBN3709_n_46337), .d(n_10636), .o(n_46381) );
no02f80 g739213 ( .a(n_40692), .b(n_40707), .o(n_40796) );
no02f80 g744651 ( .a(n_35267), .b(n_35252), .o(n_35349) );
in01f80 g752367 ( .a(n_27783), .o(n_27756) );
oa22f80 g739830 ( .a(n_40412), .b(n_40365), .c(n_40432), .d(n_40366), .o(n_40457) );
in01f80 g757465 ( .a(n_22835), .o(n_22804) );
in01f80 newInst_1616 ( .a(newNet_1615), .o(newNet_1616) );
oa22f80 g784372 ( .a(FE_OFN806_n_46196), .b(FE_OCP_RBN3115_n_6379), .c(FE_OFN84_n_46137), .d(n_6379), .o(n_46178) );
na02f80 g778378 ( .a(n_2453), .b(n_2206), .o(n_2469) );
in01f80 g761123 ( .a(n_19300), .o(n_19498) );
in01f80 FE_OCP_RBC3133_n_27736 ( .a(n_27736), .o(FE_OCP_RBN3133_n_27736) );
no02f80 g743116 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_), .o(n_37205) );
ao12f80 g740805 ( .a(n_39280), .b(n_39381), .c(n_39279), .o(n_39466) );
in01f80 g737601 ( .a(n_42489), .o(n_42490) );
na02f80 g756582 ( .a(n_23574), .b(n_22630), .o(n_23682) );
no02f80 g774330 ( .a(FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_5_), .o(n_6531) );
oa12f80 g766468 ( .a(n_14066), .b(n_14065), .c(n_14064), .o(n_15935) );
in01f80 newInst_1581 ( .a(newNet_1580), .o(newNet_1581) );
na02f80 g771459 ( .a(n_9305), .b(n_9304), .o(n_9486) );
no02f80 g746549 ( .a(n_34442), .b(n_34441), .o(n_34443) );
oa12f80 g777816 ( .a(n_2710), .b(n_3212), .c(n_2651), .o(n_3410) );
in01f80 g744694 ( .a(n_36575), .o(n_36576) );
in01f80 g753727 ( .a(n_26557), .o(n_26558) );
in01f80 newInst_2022 ( .a(newNet_1665), .o(newNet_2022) );
in01f80 newInst_3726 ( .a(newNet_3725), .o(newNet_3726) );
in01f80 g777821 ( .a(n_3299), .o(n_3300) );
oa12f80 g757457 ( .a(n_22959), .b(n_22935), .c(n_44083), .o(n_23172) );
no02f80 FE_RC_3017_0 ( .a(n_35122), .b(FE_RN_1323_0), .o(n_35178) );
in01f80 g736853 ( .a(n_43619), .o(n_43620) );
na02f80 g752829 ( .a(n_27469), .b(n_26464), .o(n_27510) );
no02f80 g743865 ( .a(n_35987), .b(n_35827), .o(n_35988) );
na02f80 FE_RC_3260_0 ( .a(FE_RN_1437_0), .b(FE_RN_1438_0), .o(FE_RN_1439_0) );
in01f80 g758422 ( .a(FE_OFN738_n_22641), .o(n_23354) );
in01f80 g769378 ( .a(n_11935), .o(n_11936) );
oa22f80 g784361 ( .a(FE_OFN774_n_46137), .b(n_6212), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_6233), .o(n_46167) );
in01f80 g746626 ( .a(n_34911), .o(n_34912) );
na02f80 g777781 ( .a(n_3379), .b(n_3378), .o(n_3457) );
no02f80 g751045 ( .a(n_30090), .b(n_29995), .o(n_30616) );
ao12f80 g741229 ( .a(n_39000), .b(FE_OCP_RBN3580_n_44944), .c(n_38912), .o(n_39453) );
oa12f80 g760486 ( .a(n_19930), .b(n_20423), .c(n_19911), .o(n_20624) );
ao12f80 g774212 ( .a(n_6658), .b(n_6591), .c(n_6630), .o(n_6753) );
no02f80 g766938 ( .a(n_14293), .b(n_14208), .o(n_15029) );
na02f80 g761015 ( .a(n_19285), .b(n_19218), .o(n_19322) );
in01f80 g740280 ( .a(n_40361), .o(n_40362) );
no02f80 g764685 ( .a(n_16030), .b(n_15938), .o(n_15945) );
na02f80 g757657 ( .a(n_22613), .b(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n_22994) );
in01f80 g776510 ( .a(n_4542), .o(n_4601) );
no02f80 FE_RC_1414_0 ( .a(FE_RN_411_0), .b(FE_RN_412_0), .o(FE_RN_413_0) );
no02f80 g781310 ( .a(n_7), .b(n_47), .o(n_48) );
ao22s80 g780229 ( .a(n_970), .b(FE_OFN761_n_45813), .c(n_904), .d(n_1203), .o(n_1028) );
no02f80 g738062 ( .a(n_42087), .b(n_41881), .o(n_42109) );
in01f80 g779690 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .o(n_1370) );
in01f80 g738870 ( .a(n_41347), .o(n_41637) );
in01f80 g747501 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_3_), .o(n_32351) );
in01f80 g766551 ( .a(n_13995), .o(n_13996) );
in01f80 newInst_2281 ( .a(newNet_479), .o(newNet_2281) );
in01f80 g739203 ( .a(n_40863), .o(n_40864) );
na02f80 g752151 ( .a(n_28667), .b(n_28666), .o(n_28668) );
in01f80 g777357 ( .a(n_4999), .o(n_5000) );
na02f80 g757320 ( .a(n_23002), .b(n_23020), .o(n_23137) );
na02f80 g780186 ( .a(n_1128), .b(n_45814), .o(n_1162) );
no02f80 g754739 ( .a(n_26160), .b(n_25684), .o(n_26381) );
in01f80 fopt783994 ( .a(n_45718), .o(n_45717) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_4_ ( .ck(newNet_554), .d(n_16863), .o(delay_xor_ln22_unr12_stage5_stallmux_q_4_) );
na02f80 g743392 ( .a(n_36657), .b(n_36589), .o(n_36658) );
no02f80 g745847 ( .a(n_34140), .b(n_34139), .o(n_34141) );
in01f80 newInst_1898 ( .a(newNet_1897), .o(newNet_1898) );
in01f80 newInst_1822 ( .a(newNet_1821), .o(newNet_1822) );
no02f80 g777167 ( .a(n_4901), .b(n_4818), .o(n_5873) );
no02f80 g776072 ( .a(n_5021), .b(n_5010), .o(n_5093) );
na03f80 FE_RC_3579_0 ( .a(n_14478), .b(FE_RN_1556_0), .c(FE_RN_1557_0), .o(FE_RN_1558_0) );
in01f80 g742294 ( .a(FE_OCP_RBN2257_n_37844), .o(n_37945) );
na02f80 g742750 ( .a(n_37393), .b(n_37392), .o(n_37394) );
in01f80 g749616 ( .a(n_30526), .o(n_30505) );
no02f80 g749712 ( .a(n_31290), .b(n_31342), .o(n_31348) );
na02f80 g760191 ( .a(n_20433), .b(n_20391), .o(n_20526) );
no02f80 g770416 ( .a(n_10586), .b(n_10508), .o(n_10609) );
in01f80 g744629 ( .a(n_35328), .o(n_35396) );
oa12f80 g746571 ( .a(n_34609), .b(n_34666), .c(n_34585), .o(n_35071) );
oa12f80 g762665 ( .a(n_17870), .b(n_17928), .c(n_17822), .o(n_18000) );
na02f80 g750015 ( .a(n_30924), .b(n_30267), .o(n_31044) );
in01f80 g745181 ( .a(n_34712), .o(n_34676) );
in01f80 g780360 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_), .o(n_944) );
in01f80 FE_RC_812_0 ( .a(n_29092), .o(FE_RN_244_0) );
in01f80 g740635 ( .a(n_39989), .o(n_39605) );
na02f80 g775536 ( .a(FE_OCP_RBN2942_n_5454), .b(FE_OCP_RBN2733_n_4219), .o(n_5522) );
in01f80 newInst_611 ( .a(newNet_610), .o(newNet_611) );
na02f80 g741642 ( .a(n_38541), .b(n_38555), .o(n_38912) );
in01f80 g749780 ( .a(n_31388), .o(n_31389) );
no02f80 g738246 ( .a(n_41896), .b(n_41675), .o(n_41897) );
in01f80 g773505 ( .a(n_7560), .o(n_7543) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_2_ ( .ck(newNet_3497), .d(n_21173), .o(delay_add_ln22_unr14_stage6_stallmux_q_2_) );
in01f80 g769235 ( .a(n_12493), .o(n_12494) );
no02f80 g781148 ( .a(n_209), .b(n_264), .o(n_213) );
in01f80 FE_OCP_RBC3005_n_11087 ( .a(n_11087), .o(FE_OCP_RBN3005_n_11087) );
in01f80 g739757 ( .a(n_40472), .o(n_40505) );
na02f80 g749108 ( .a(n_30879), .b(n_30912), .o(n_31026) );
na02f80 g762750 ( .a(n_18197), .b(n_17615), .o(n_18235) );
in01f80 g756497 ( .a(n_23943), .o(n_23944) );
no02f80 g737788 ( .a(n_42187), .b(n_42204), .o(n_42208) );
na02f80 g772356 ( .a(n_8477), .b(n_8413), .o(n_8478) );
na02f80 g747842 ( .a(n_33238), .b(n_33336), .o(n_33391) );
no02f80 g763289 ( .a(n_17045), .b(n_16952), .o(n_17043) );
in01f80 g766530 ( .a(n_14062), .o(n_14063) );
in01f80 newInst_1023 ( .a(newNet_1022), .o(newNet_1023) );
na02f80 g762198 ( .a(n_18190), .b(n_17922), .o(n_18192) );
no02f80 g748928 ( .a(n_30967), .b(n_30890), .o(n_31014) );
in01f80 g754630 ( .a(n_27246), .o(n_27518) );
in01f80 FE_OCP_RBC2872_n_39542 ( .a(n_39542), .o(FE_OCP_RBN2872_n_39542) );
na02f80 g769564 ( .a(n_11425), .b(n_11424), .o(n_11464) );
ao12f80 g749144 ( .a(n_31529), .b(n_32116), .c(n_31570), .o(n_32206) );
na02f80 g774287 ( .a(n_6830), .b(n_6703), .o(n_6704) );
in01f80 g780862 ( .a(FE_OFN50_n_1045), .o(n_563) );
na02f80 g767023 ( .a(FE_OCP_RBN3529_n_13765), .b(n_13961), .o(n_14108) );
in01f80 g772462 ( .a(n_8540), .o(n_8541) );
oa12f80 g770560 ( .a(n_10162), .b(n_10170), .c(n_10261), .o(n_10481) );
na02f80 g775391 ( .a(n_5436), .b(n_5057), .o(n_5480) );
na02f80 g778650 ( .a(n_2382), .b(n_2027), .o(n_2441) );
in01f80 g778078 ( .a(n_4642), .o(n_3025) );
in01f80 g741237 ( .a(n_38882), .o(n_38915) );
in01f80 g758809 ( .a(n_21807), .o(n_21808) );
no02f80 g740036 ( .a(n_39845), .b(n_39872), .o(n_39873) );
oa12f80 g772512 ( .a(n_8646), .b(n_8645), .c(n_8644), .o(n_9478) );
no02f80 g764631 ( .a(n_16071), .b(FE_OCP_RBN2483_n_14326), .o(n_16180) );
in01f80 FE_OCP_RBC2869_n_10480 ( .a(n_10480), .o(FE_OCP_RBN2869_n_10480) );
na02f80 g774147 ( .a(n_6654), .b(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n_6655) );
oa12f80 g770767 ( .a(n_9601), .b(n_10255), .c(n_9695), .o(n_10373) );
in01f80 FE_OCP_RBC1149_n_27962 ( .a(n_27962), .o(FE_OCP_RBN1149_n_27962) );
in01f80 g753949 ( .a(n_26219), .o(n_26258) );
in01f80 fopt782858 ( .a(n_22028), .o(n_44288) );
in01f80 g752149 ( .a(n_28090), .o(n_28091) );
na02f80 g778677 ( .a(n_2277), .b(n_2270), .o(n_2331) );
oa12f80 g768478 ( .a(n_12406), .b(n_45659), .c(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .o(n_12454) );
na02f80 g769390 ( .a(n_11377), .b(FE_OCP_RBN2861_n_10399), .o(n_11407) );
na02f80 g776436 ( .a(n_4378), .b(n_3951), .o(n_4625) );
no02f80 g767361 ( .a(n_13435), .b(FE_OCPN1472_n_13434), .o(n_13451) );
in01f80 FE_OCP_DRV_C3158_n_27062 ( .a(FE_OCP_DRV_N3157_n_27062), .o(FE_OCP_DRV_N3158_n_27062) );
in01f80 g742892 ( .a(n_37419), .o(n_37078) );
no02f80 g741941 ( .a(n_38185), .b(n_37654), .o(n_38203) );
in01f80 g757477 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_10_), .o(n_23033) );
in01f80 newInst_2122 ( .a(newNet_2121), .o(newNet_2122) );
in01f80 g756805 ( .a(n_23471), .o(n_23472) );
no02f80 g742257 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37901), .o(n_38266) );
in01f80 g744659 ( .a(n_36599), .o(n_36600) );
in01f80 g773876 ( .a(n_7028), .o(n_7015) );
in01f80 newInst_188 ( .a(newNet_76), .o(newNet_188) );
na02f80 g739568 ( .a(n_40608), .b(n_45513), .o(n_40629) );
no02f80 g748651 ( .a(n_31400), .b(n_31074), .o(n_31422) );
in01f80 newInst_1631 ( .a(newNet_1630), .o(newNet_1631) );
na02f80 g777177 ( .a(n_3940), .b(n_3816), .o(n_4084) );
no02f80 g769120 ( .a(n_11623), .b(n_11608), .o(n_11747) );
ms00f80 cos_out_reg_21_ ( .ck(newNet_3719), .d(n_43865), .o(cos_out_21) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_14_ ( .ck(newNet_2409), .d(n_36345), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_14_) );
in01f80 g743535 ( .a(n_36629), .o(n_36607) );
in01f80 g739279 ( .a(n_44026), .o(n_40780) );
in01f80 g768552 ( .a(n_12328), .o(n_12329) );
na02f80 g738513 ( .a(n_41582), .b(n_41291), .o(n_41694) );
oa22f80 FE_RC_1139_0 ( .a(n_36301), .b(n_36560), .c(n_36302), .d(n_36546), .o(n_36669) );
na02f80 g784078 ( .a(n_7598), .b(n_45824), .o(n_45825) );
in01f80 g748849 ( .a(n_31111), .o(n_31112) );
in01f80 g766246 ( .a(n_14547), .o(n_14498) );
in01f80 FE_OCP_RBC2994_n_35539 ( .a(FE_OCP_RBN2991_n_35539), .o(FE_OCP_RBN2994_n_35539) );
no02f80 g747324 ( .a(n_32440), .b(n_44962), .o(n_32527) );
oa12f80 g745860 ( .a(n_44112), .b(n_34004), .c(n_33942), .o(n_34429) );
oa12f80 g769102 ( .a(n_45685), .b(n_12014), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_24_), .o(n_12085) );
na02f80 g763306 ( .a(n_17040), .b(n_16915), .o(n_17085) );
in01f80 FE_RC_2505_0 ( .a(n_17765), .o(FE_RN_1017_0) );
oa12f80 g750350 ( .a(n_29727), .b(n_29739), .c(n_29737), .o(n_29789) );
na02f80 g778105 ( .a(n_2965), .b(n_2999), .o(n_3026) );
in01f80 newInst_2907 ( .a(newNet_2906), .o(newNet_2907) );
na02f80 g741190 ( .a(FE_OCP_RBN2636_n_38806), .b(n_38919), .o(n_39009) );
in01f80 newInst_812 ( .a(newNet_811), .o(newNet_812) );
na02f80 g778318 ( .a(n_2910), .b(delay_add_ln22_unr2_stage2_stallmux_q_30_), .o(n_2927) );
in01f80 g753269 ( .a(n_27462), .o(n_27415) );
na02f80 FE_RC_2551_0 ( .a(n_34078), .b(FE_RN_1044_0), .o(n_34124) );
no02f80 g768867 ( .a(n_11736), .b(n_11821), .o(n_11958) );
ao12f80 g775746 ( .a(n_5291), .b(n_5367), .c(n_5290), .o(n_5418) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_30_ ( .ck(newNet_1699), .d(n_22689), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_30_) );
no02f80 g757393 ( .a(n_44084), .b(delay_xor_ln21_unr15_stage6_stallmux_q_8_), .o(n_23229) );
no02f80 g764973 ( .a(n_15610), .b(n_15609), .o(n_15541) );
oa22f80 g748703 ( .a(n_32460), .b(n_32479), .c(n_32539), .d(n_32480), .o(n_33240) );
no02f80 g777623 ( .a(n_3481), .b(n_2759), .o(n_3559) );
ao12f80 g759796 ( .a(n_21446), .b(n_21714), .c(n_21481), .o(n_22176) );
oa12f80 g777014 ( .a(n_3668), .b(n_3689), .c(n_3029), .o(n_3764) );
oa12f80 g764666 ( .a(n_15373), .b(n_15808), .c(n_15806), .o(n_15820) );
no02f80 g762280 ( .a(n_18584), .b(n_18609), .o(n_19159) );
na02f80 g773473 ( .a(n_7491), .b(n_7278), .o(n_7558) );
no02f80 g741948 ( .a(n_38110), .b(n_38167), .o(n_38168) );
na02f80 g757427 ( .a(n_22964), .b(n_22988), .o(n_23100) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_1_ ( .ck(newNet_2564), .d(n_26365), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_1_) );
in01f80 newInst_1980 ( .a(newNet_820), .o(newNet_1980) );
in01f80 g739046 ( .a(n_41121), .o(n_41122) );
na02f80 g740539 ( .a(n_39714), .b(n_39715), .o(n_39746) );
na02f80 g775712 ( .a(n_5159), .b(n_5071), .o(n_5160) );
in01f80 newInst_1857 ( .a(newNet_1856), .o(newNet_1857) );
in01f80 g757890 ( .a(n_23026), .o(n_23008) );
no02f80 g749271 ( .a(n_30843), .b(n_30760), .o(n_30869) );
ms00f80 sin_out_reg_19_ ( .ck(newNet_64), .d(n_43896), .o(sin_out_19) );
no02f80 g778122 ( .a(n_2845), .b(n_2534), .o(n_2924) );
oa12f80 g770637 ( .a(n_10094), .b(n_10181), .c(n_10025), .o(n_10328) );
no02f80 g744121 ( .a(n_47265), .b(n_35900), .o(n_35901) );
na02f80 g761653 ( .a(n_19403), .b(n_18811), .o(n_19495) );
in01f80 g764237 ( .a(n_16516), .o(n_16580) );
ao12f80 g757627 ( .a(n_22078), .b(n_45721), .c(n_22079), .o(n_22619) );
na02f80 FE_RC_2399_0 ( .a(FE_RN_944_0), .b(n_42592), .o(FE_RN_945_0) );
no02f80 g779177 ( .a(n_1898), .b(delay_add_ln22_unr2_stage2_stallmux_q_10_), .o(n_1903) );
ao12f80 g751333 ( .a(n_29512), .b(n_29511), .c(n_29510), .o(n_29940) );
in01f80 FE_OCPC992_n_22249 ( .a(FE_OCPN990_n_22249), .o(FE_OCPN992_n_22249) );
no02f80 g778682 ( .a(n_45903), .b(n_2606), .o(n_2249) );
na02f80 g771256 ( .a(n_9350), .b(n_9288), .o(n_9457) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_1_ ( .ck(newNet_3056), .d(n_1122), .o(delay_add_ln22_unr2_stage2_stallmux_q_1_) );
in01f80 g753630 ( .a(n_26661), .o(n_26662) );
in01f80 newInst_1244 ( .a(newNet_561), .o(newNet_1244) );
in01f80 FE_OCP_RBC2728_n_4219 ( .a(FE_OCP_RBN2725_n_4219), .o(FE_OCP_RBN2728_n_4219) );
in01f80 g763217 ( .a(n_17009), .o(n_17048) );
in01f80 g778050 ( .a(n_3066), .o(n_3067) );
no03m80 g743347 ( .a(n_37726), .b(n_37789), .c(n_37731), .o(n_37790) );
in01f80 g754402 ( .a(n_45533), .o(n_25808) );
in01f80 FE_OCPC1489_n_30823 ( .a(n_30823), .o(FE_OCPN1489_n_30823) );
ao12f80 g760757 ( .a(n_20089), .b(n_20088), .c(n_20087), .o(n_20156) );
in01f80 g767386 ( .a(n_13446), .o(n_13447) );
no02f80 g769682 ( .a(n_11209), .b(n_46424), .o(n_11227) );
no02f80 g741267 ( .a(FE_OCP_RBN3582_n_44944), .b(n_38553), .o(n_39395) );
na02f80 g756435 ( .a(n_23855), .b(n_23816), .o(n_24040) );
ao12f80 g739384 ( .a(n_40904), .b(n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n_40969) );
no02f80 g761477 ( .a(n_19845), .b(n_19900), .o(n_19954) );
in01f80 g768673 ( .a(n_12240), .o(n_12189) );
na02f80 g773168 ( .a(n_7721), .b(n_7771), .o(n_7921) );
in01f80 g765697 ( .a(n_16338), .o(n_17584) );
in01f80 g738999 ( .a(n_41186), .o(n_41207) );
na02f80 g750820 ( .a(n_29188), .b(n_29187), .o(n_29189) );
na02f80 g753238 ( .a(n_27110), .b(n_45533), .o(n_27175) );
na02f80 g754872 ( .a(n_25564), .b(n_25543), .o(n_25622) );
in01f80 g769158 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_2_), .o(n_11594) );
no02f80 g769278 ( .a(n_11582), .b(n_11581), .o(n_11583) );
in01f80 g780542 ( .a(n_778), .o(n_724) );
in01f80 g746854 ( .a(n_33059), .o(n_33060) );
in01f80 g744821 ( .a(n_36476), .o(n_36494) );
in01f80 g775084 ( .a(n_6106), .o(n_6107) );
in01f80 FE_RC_3716_0 ( .a(n_5677), .o(FE_RN_1634_0) );
in01f80 newInst_3288 ( .a(newNet_3287), .o(newNet_3288) );
oa22f80 g747766 ( .a(n_33571), .b(n_33362), .c(n_33372), .d(n_33396), .o(n_33758) );
na02f80 g741757 ( .a(n_38369), .b(n_38168), .o(n_38506) );
no02f80 g778712 ( .a(n_2438), .b(n_2057), .o(n_3108) );
na02f80 g774460 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n_6864) );
oa12f80 g758912 ( .a(n_22059), .b(n_22058), .c(n_22057), .o(n_22116) );
ao12f80 g763776 ( .a(n_17093), .b(n_17261), .c(n_17057), .o(n_17262) );
na02f80 g737069 ( .a(n_43097), .b(n_43123), .o(n_43165) );
in01f80 FE_RC_2358_0 ( .a(n_18884), .o(FE_RN_910_0) );
na02f80 g780701 ( .a(n_638), .b(n_637), .o(n_639) );
in01f80 g748230 ( .a(n_32072), .o(n_32073) );
na02f80 g740086 ( .a(n_40003), .b(n_39941), .o(n_40004) );
in01f80 g753567 ( .a(n_26778), .o(n_26779) );
in01f80 g766185 ( .a(n_14572), .o(n_14593) );
in01f80 g772474 ( .a(n_8388), .o(n_8750) );
in01f80 newInst_3361 ( .a(newNet_3360), .o(newNet_3361) );
na02f80 g750042 ( .a(n_29846), .b(n_28831), .o(n_29968) );
na02f80 g762391 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18487), .o(n_18608) );
ao12f80 g764509 ( .a(n_46980), .b(n_16154), .c(n_16111), .o(n_16155) );
in01f80 g737925 ( .a(n_42514), .o(n_42515) );
oa12f80 g770843 ( .a(n_10133), .b(n_10132), .c(n_10171), .o(n_10213) );
na02f80 FE_RC_2351_0 ( .a(n_1682), .b(n_1681), .o(FE_RN_904_0) );
in01f80 g751986 ( .a(n_28905), .o(n_28878) );
na02f80 g756386 ( .a(n_23692), .b(n_23479), .o(n_23795) );
no03m80 g746101 ( .a(FE_OCP_RBN1355_n_44259), .b(n_33698), .c(n_33782), .o(n_33833) );
no02f80 g769296 ( .a(FE_OCP_RBN3093_n_11475), .b(n_10936), .o(n_11578) );
in01f80 g769635 ( .a(n_11279), .o(n_11280) );
no02f80 g736725 ( .a(n_43029), .b(n_43042), .o(n_43074) );
oa22f80 g780534 ( .a(n_890), .b(n_422), .c(n_923), .d(n_412), .o(n_1109) );
oa22f80 g750037 ( .a(FE_OCPN1786_n_30134), .b(FE_OCP_RBN2341_n_29470), .c(FE_OCP_RBN2571_n_29922), .d(n_45489), .o(n_30385) );
in01f80 g744223 ( .a(n_36287), .o(n_36288) );
oa12f80 g750658 ( .a(n_28798), .b(n_29279), .c(n_28804), .o(n_29329) );
in01f80 FE_RC_3070_0 ( .a(n_26176), .o(FE_RN_1350_0) );
ao12f80 g738457 ( .a(n_41509), .b(n_41508), .c(n_41507), .o(n_42211) );
in01f80 newInst_1912 ( .a(newNet_1911), .o(newNet_1912) );
in01f80 newInst_365 ( .a(newNet_364), .o(newNet_365) );
oa22f80 g741099 ( .a(FE_OCP_RBN3629_n_38870), .b(n_38493), .c(FE_OCPN957_n_39096), .d(n_38516), .o(n_39500) );
no02f80 g754698 ( .a(n_26231), .b(n_26348), .o(n_26716) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_27_ ( .ck(newNet_1493), .d(n_32342), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_) );
no02f80 g779766 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_5_), .o(n_1543) );
in01f80 g764034 ( .a(n_17900), .o(n_18032) );
ao22s80 FE_RC_1938_0 ( .a(FE_OFN788_n_25834), .b(FE_OCP_RBN2346_n_29448), .c(n_29561), .d(n_29448), .o(n_29545) );
no02f80 g760574 ( .a(n_19888), .b(n_19816), .o(n_19889) );
in01f80 g756503 ( .a(n_23786), .o(n_23787) );
in01f80 g739847 ( .a(n_40349), .o(n_40383) );
no02f80 g771228 ( .a(n_9791), .b(n_9790), .o(n_9918) );
in01f80 newInst_952 ( .a(newNet_226), .o(newNet_952) );
in01f80 g774930 ( .a(n_6268), .o(n_6269) );
in01f80 g759396 ( .a(n_21118), .o(n_22076) );
oa12f80 g749374 ( .a(n_31348), .b(n_31981), .c(n_31341), .o(n_32008) );
in01f80 newInst_3599 ( .a(newNet_3598), .o(newNet_3599) );
no02f80 g751037 ( .a(n_30094), .b(n_30059), .o(n_30159) );
in01f80 newInst_1832 ( .a(newNet_1831), .o(newNet_1832) );
in01f80 FE_OCP_RBC3242_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3242_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
in01f80 FE_OCP_RBC1729_n_20903 ( .a(n_20903), .o(FE_OCP_RBN1729_n_20903) );
in01f80 g773241 ( .a(n_7600), .o(n_7601) );
in01f80 g743386 ( .a(n_36718), .o(n_36719) );
no02f80 g774293 ( .a(n_6684), .b(n_6683), .o(n_7056) );
oa12f80 g738447 ( .a(n_41523), .b(FE_OCPN953_n_41540), .c(n_41433), .o(n_41841) );
ms00f80 delay_sub_ln23_0_unr17_stage7_stallmux_q_reg ( .ck(newNet_1671), .d(n_24188), .o(n_44722) );
in01f80 g778216 ( .a(n_2778), .o(n_2852) );
na02f80 g750172 ( .a(n_30923), .b(n_30900), .o(n_30901) );
na02f80 g769323 ( .a(FE_OCPN867_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_21_), .o(n_11894) );
na02f80 g779229 ( .a(n_1823), .b(delay_add_ln22_unr2_stage2_stallmux_q_8_), .o(n_1892) );
oa22f80 FE_RC_718_0 ( .a(FE_OCP_RBN2337_n_8269), .b(FE_OCP_RBN3453_FE_OCPN1240_n_7721), .c(n_8269), .d(FE_OCPN940_n_7712), .o(n_8107) );
na02f80 g781020 ( .a(cos_out_9), .b(FE_OFN2_n_43918), .o(n_314) );
oa12f80 g776266 ( .a(n_4365), .b(n_4323), .c(n_4248), .o(n_4454) );
no02f80 g753887 ( .a(n_26297), .b(FE_OCPN1528_n_26296), .o(n_26403) );
in01f80 g763397 ( .a(n_16996), .o(n_17035) );
no02f80 g757225 ( .a(n_23470), .b(n_22853), .o(n_23523) );
no02f80 g746801 ( .a(n_33102), .b(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n_33103) );
no02f80 g742411 ( .a(FE_OCP_RBN2212_n_37720), .b(n_38047), .o(n_37743) );
in01f80 newInst_1015 ( .a(newNet_1014), .o(newNet_1015) );
oa12f80 g780029 ( .a(n_866), .b(n_1250), .c(n_929), .o(n_1259) );
oa22f80 FE_RC_989_0 ( .a(n_24350), .b(n_27805), .c(n_27796), .d(n_45132), .o(n_27863) );
na02f80 g737418 ( .a(n_42736), .b(n_42428), .o(n_42796) );
in01f80 FE_OCP_RBC3067_n_43230 ( .a(n_43230), .o(FE_OCP_RBN3067_n_43230) );
in01f80 newInst_3485 ( .a(newNet_3484), .o(newNet_3485) );
in01f80 g751177 ( .a(n_30000), .o(n_29939) );
ao12f80 g772699 ( .a(n_8102), .b(n_8204), .c(n_8158), .o(n_8275) );
in01f80 FE_RC_3219_0 ( .a(FE_RN_1429_0), .o(FE_RN_1428_0) );
no02f80 g766008 ( .a(n_14668), .b(n_14649), .o(n_14774) );
in01f80 g742019 ( .a(n_38042), .o(n_38012) );
ao12f80 g760979 ( .a(n_19272), .b(n_19278), .c(n_19169), .o(n_19279) );
in01f80 g777830 ( .a(n_3255), .o(n_3293) );
na02f80 g759771 ( .a(n_20712), .b(n_20634), .o(n_20754) );
na02f80 g761161 ( .a(n_19104), .b(n_19057), .o(n_19168) );
no02f80 g776097 ( .a(n_5048), .b(FE_OCP_RBN2669_n_4158), .o(n_5021) );
in01f80 g753207 ( .a(n_27425), .o(n_27343) );
in01f80 g759568 ( .a(n_20878), .o(n_20904) );
in01f80 newInst_1234 ( .a(newNet_1233), .o(newNet_1234) );
no02f80 g746539 ( .a(n_34546), .b(n_34496), .o(n_34915) );
in01f80 g749460 ( .a(n_30514), .o(n_30535) );
in01f80 g756254 ( .a(n_24767), .o(n_24768) );
ao12f80 g748205 ( .a(n_32764), .b(n_32780), .c(n_32763), .o(n_33281) );
oa12f80 g755424 ( .a(n_25527), .b(n_25526), .c(n_25525), .o(n_26230) );
na02f80 g744604 ( .a(n_35293), .b(n_35292), .o(n_35317) );
na02f80 g755819 ( .a(n_24314), .b(n_24013), .o(n_24315) );
in01f80 FE_OCPC1761_n_37877 ( .a(n_37877), .o(FE_OCPN1761_n_37877) );
in01f80 g754813 ( .a(n_25363), .o(n_25364) );
oa22f80 FE_RC_2933_0 ( .a(n_44463), .b(FE_OCP_RBN2917_n_10644), .c(FE_OCP_RBN3646_n_44490), .d(n_10644), .o(FE_RN_1278_0) );
na02f80 g738979 ( .a(n_41155), .b(n_41208), .o(n_41209) );
in01f80 g760087 ( .a(n_20375), .o(n_20409) );
na02f80 g740193 ( .a(n_39796), .b(n_39795), .o(n_39814) );
in01f80 g741394 ( .a(FE_OCP_RBN2639_n_38806), .o(n_38847) );
oa22f80 g775571 ( .a(n_5236), .b(n_5169), .c(n_5206), .d(n_5170), .o(n_5397) );
oa12f80 g761901 ( .a(n_18467), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n_18637) );
no02f80 g765294 ( .a(n_15781), .b(n_15869), .o(n_15827) );
in01f80 g770272 ( .a(n_10736), .o(n_10737) );
no02f80 g745069 ( .a(n_36233), .b(n_35654), .o(n_36313) );
in01f80 newInst_1449 ( .a(newNet_1448), .o(newNet_1449) );
na02f80 g773164 ( .a(n_7802), .b(n_7794), .o(n_7889) );
in01f80 FE_RC_3615_0 ( .a(n_20422), .o(n_20445) );
na02f80 g765873 ( .a(n_14796), .b(n_14859), .o(n_14860) );
no02f80 g767861 ( .a(n_12922), .b(n_12435), .o(n_13084) );
no02f80 g773736 ( .a(n_7240), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_15_), .o(n_7262) );
in01f80 newInst_2678 ( .a(newNet_144), .o(newNet_2678) );
na02f80 g772495 ( .a(n_8590), .b(n_8591), .o(n_8685) );
oa12f80 g756391 ( .a(n_23834), .b(n_24259), .c(n_24169), .o(n_24301) );
in01f80 newInst_2550 ( .a(newNet_1938), .o(newNet_2550) );
no02f80 g776335 ( .a(n_4197), .b(n_4065), .o(n_4319) );
no02f80 g775620 ( .a(n_5458), .b(n_4606), .o(n_5512) );
in01f80 g777881 ( .a(n_3239), .o(n_3261) );
na02f80 g739132 ( .a(n_40991), .b(n_41006), .o(n_41055) );
in01f80 newInst_764 ( .a(newNet_763), .o(newNet_764) );
no02f80 g748711 ( .a(n_32539), .b(n_32508), .o(n_32509) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_23_ ( .ck(newNet_1508), .d(n_32274), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_) );
in01f80 g744620 ( .a(n_35329), .o(n_35346) );
no02f80 g742174 ( .a(n_44887), .b(n_38270), .o(n_38307) );
no02f80 g765881 ( .a(n_14800), .b(n_14856), .o(n_14857) );
oa12f80 g739696 ( .a(n_40211), .b(n_40543), .c(n_40251), .o(n_40565) );
in01f80 g753484 ( .a(n_26915), .o(n_26916) );
ao12f80 g738110 ( .a(n_42084), .b(n_42105), .c(n_42083), .o(n_42158) );
ao12f80 g756510 ( .a(n_23878), .b(n_23783), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_25_), .o(n_23917) );
no02f80 g776292 ( .a(n_4604), .b(n_4160), .o(n_4733) );
ao12f80 g778218 ( .a(n_2668), .b(n_2667), .c(n_2709), .o(n_4339) );
no02f80 g773005 ( .a(n_7775), .b(n_7807), .o(n_7831) );
no02f80 g773794 ( .a(n_7137), .b(n_7033), .o(n_7159) );
na02f80 g746023 ( .a(n_33719), .b(n_33646), .o(n_33787) );
in01f80 FE_OFC745_n_23604 ( .a(FE_OFN744_n_23604), .o(FE_OFN745_n_23604) );
in01f80 g769572 ( .a(n_11495), .o(n_11605) );
na02f80 FE_RC_3020_0 ( .a(n_47268), .b(FE_RN_1324_0), .o(n_16735) );
na02f80 g775263 ( .a(n_5834), .b(n_5866), .o(n_5972) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_6_ ( .ck(newNet_3102), .d(n_40427), .o(delay_add_ln22_unr27_stage10_stallmux_q_6_) );
na02f80 g739222 ( .a(n_40740), .b(n_40739), .o(n_40741) );
no02f80 g773833 ( .a(n_7103), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .o(n_7132) );
oa12f80 g770538 ( .a(n_46420), .b(n_10465), .c(FE_OCP_RBN3560_n_8809), .o(n_10554) );
in01f80 g741308 ( .a(n_38902), .o(n_38903) );
in01f80 g776024 ( .a(n_5140), .o(n_5141) );
na02f80 g775333 ( .a(n_5863), .b(n_5862), .o(n_5864) );
ao12f80 g752456 ( .a(n_27411), .b(n_27648), .c(n_27337), .o(n_27696) );
in01f80 g757672 ( .a(n_22640), .o(n_22617) );
no02f80 g753944 ( .a(n_26173), .b(FE_OCPN1508_n_23414), .o(n_26222) );
oa22f80 FE_RC_553_0 ( .a(FE_OCP_RBN2828_n_30731), .b(FE_OCP_DRV_N3158_n_27062), .c(FE_OCPN1410_n_27014), .d(n_30731), .o(n_30847) );
in01f80 newInst_1509 ( .a(newNet_137), .o(newNet_1509) );
in01f80 FE_OCP_RBC3058_n_36515 ( .a(n_36515), .o(FE_OCP_RBN3058_n_36515) );
na02f80 g753253 ( .a(n_27287), .b(n_25851), .o(n_27334) );
in01f80 newInst_915 ( .a(newNet_914), .o(newNet_915) );
in01f80 FE_RC_4184_0 ( .a(FE_RN_1829_0), .o(FE_RN_1821_0) );
na02f80 g766999 ( .a(n_13497), .b(FE_OCPN860_n_12880), .o(n_13567) );
in01f80 g771965 ( .a(n_9770), .o(n_9870) );
in01f80 g754655 ( .a(FE_OCPN1410_n_27014), .o(n_27131) );
no02f80 g778234 ( .a(n_2667), .b(n_2709), .o(n_2668) );
oa12f80 g752776 ( .a(n_26875), .b(n_27075), .c(n_26960), .o(n_27193) );
no02f80 g742180 ( .a(n_44867), .b(n_37935), .o(n_38003) );
oa22f80 g750992 ( .a(n_28890), .b(n_28914), .c(n_28933), .d(n_28915), .o(n_30399) );
in01f80 g742954 ( .a(n_37193), .o(n_37194) );
in01f80 newInst_1447 ( .a(newNet_1446), .o(newNet_1447) );
no02f80 g739283 ( .a(n_40773), .b(n_40813), .o(n_40856) );
na03f80 FE_RC_3442_0 ( .a(FE_OCP_RBN3857_FE_RN_779_0), .b(n_22185), .c(FE_RN_1286_0), .o(FE_RN_1287_0) );
oa22f80 g749111 ( .a(n_32201), .b(n_31617), .c(n_32202), .d(n_31618), .o(n_32257) );
na02f80 g767050 ( .a(FE_OCP_RBN3529_n_13765), .b(n_13502), .o(n_14006) );
in01f80 g743039 ( .a(n_37178), .o(n_37179) );
na02f80 g753896 ( .a(n_26294), .b(n_26293), .o(n_26295) );
in01f80 g780347 ( .a(n_990), .o(n_1014) );
in01f80 g740994 ( .a(n_39065), .o(n_38971) );
in01f80 g739361 ( .a(n_40785), .o(n_40758) );
no03m80 g742786 ( .a(n_37343), .b(n_37333), .c(n_37146), .o(n_37442) );
ao12f80 g773383 ( .a(n_7555), .b(n_7558), .c(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n_7574) );
in01f80 g758773 ( .a(n_21707), .o(n_21734) );
no02f80 g743931 ( .a(n_35951), .b(n_44223), .o(n_36039) );
no02f80 g767014 ( .a(FE_OCP_RBN2457_n_13765), .b(n_13325), .o(n_13904) );
no02f80 g756926 ( .a(n_24234), .b(n_24256), .o(n_24543) );
in01f80 g766657 ( .a(n_13931), .o(n_14051) );
no02f80 g739992 ( .a(n_40154), .b(FE_OCP_RBN2834_n_39586), .o(n_40155) );
na02f80 g746616 ( .a(n_34473), .b(n_34472), .o(n_34545) );
in01f80 g777949 ( .a(n_47020), .o(n_3231) );
in01f80 g781335 ( .a(n_70), .o(n_71) );
no02f80 g761324 ( .a(n_19714), .b(n_19713), .o(n_19767) );
in01f80 fopt783257 ( .a(n_44826), .o(n_44825) );
no02f80 g752342 ( .a(n_27823), .b(FE_OCP_RBN3306_n_44722), .o(n_27889) );
na02f80 g736916 ( .a(n_43038), .b(n_42803), .o(n_43183) );
na02f80 g778338 ( .a(n_2607), .b(n_2606), .o(n_2624) );
in01f80 g748155 ( .a(n_32101), .o(n_32102) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_10_ ( .ck(newNet_3658), .d(n_16183), .o(delay_add_ln22_unr11_stage5_stallmux_q_10_) );
ao22s80 g762598 ( .a(n_18000), .b(n_17925), .c(n_17949), .d(n_17924), .o(n_19590) );
in01f80 g764172 ( .a(n_16598), .o(n_16599) );
in01f80 g761966 ( .a(n_18316), .o(n_18317) );
oa22f80 g784370 ( .a(FE_OFN775_n_46137), .b(n_5613), .c(FE_OFN805_n_46196), .d(n_5645), .o(n_46176) );
na02f80 FE_RC_2496_0 ( .a(FE_OCP_RBN3306_n_44722), .b(FE_RN_1011_0), .o(n_27884) );
in01f80 g753911 ( .a(n_27067), .o(n_27063) );
na02f80 g773674 ( .a(n_7320), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_), .o(n_7371) );
in01f80 FE_RC_2841_0 ( .a(n_13618), .o(FE_RN_1222_0) );
na02f80 g775311 ( .a(n_5798), .b(n_5584), .o(n_5799) );
na02f80 g741340 ( .a(n_44944), .b(n_38496), .o(n_38900) );
no02f80 g753639 ( .a(n_26657), .b(n_26656), .o(n_26692) );
oa12f80 g739241 ( .a(n_40788), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_6_), .o(n_41001) );
ao12f80 g746255 ( .a(n_34610), .b(n_34944), .c(n_34616), .o(n_35087) );
in01f80 newInst_3302 ( .a(newNet_3301), .o(newNet_3302) );
no02f80 g779527 ( .a(n_1433), .b(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n_1515) );
in01f80 g773550 ( .a(n_7486), .o(n_7487) );
in01f80 FE_OCP_RBC2989_n_35539 ( .a(FE_OCP_RBN3698_n_35543), .o(FE_OCP_RBN2989_n_35539) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_12_ ( .ck(newNet_2023), .d(n_46988), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_12_) );
na02f80 g751957 ( .a(n_28919), .b(n_28669), .o(n_29242) );
na02f80 g766630 ( .a(n_13783), .b(n_13817), .o(n_13930) );
in01f80 g765489 ( .a(n_15920), .o(n_15921) );
in01f80 newInst_3511 ( .a(newNet_3510), .o(newNet_3511) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_31_ ( .ck(newNet_2914), .d(n_6720), .o(delay_add_ln22_unr5_stage3_stallmux_q_31_) );
in01f80 g749281 ( .a(FE_OCP_RBN3673_n_30820), .o(n_31655) );
in01f80 newInst_2345 ( .a(newNet_2344), .o(newNet_2345) );
in01f80 g773081 ( .a(n_8118), .o(n_8119) );
in01f80 newInst_3757 ( .a(newNet_3756), .o(newNet_3757) );
in01f80 g769162 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n_11593) );
in01f80 FE_OCP_RBC3032_n_43000 ( .a(n_43000), .o(FE_OCP_RBN3032_n_43000) );
oa12f80 g762897 ( .a(n_17069), .b(n_17599), .c(n_17042), .o(n_17600) );
in01f80 fopt783590 ( .a(n_35012), .o(n_45221) );
na02f80 g755723 ( .a(n_24402), .b(n_24052), .o(n_24407) );
in01f80 FE_RC_680_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_5_), .o(FE_RN_219_0) );
na02f80 g757964 ( .a(n_23116), .b(n_23054), .o(n_23532) );
oa22f80 FE_RC_3800_0 ( .a(FE_OCP_RBN2432_n_14018), .b(n_14367), .c(FE_OCP_RBN2431_n_14018), .d(n_14366), .o(n_14544) );
in01f80 g736586 ( .a(n_43682), .o(n_43678) );
na02f80 g747715 ( .a(n_32264), .b(n_32107), .o(n_32279) );
na02f80 FE_RC_2473_0 ( .a(FE_RN_993_0), .b(FE_RN_997_0), .o(n_14564) );
na02f80 FE_RC_677_0 ( .a(FE_RN_216_0), .b(FE_RN_217_0), .o(FE_RN_218_0) );
no02f80 g747049 ( .a(n_34043), .b(n_34042), .o(n_34044) );
ao12f80 g754590 ( .a(n_26609), .b(n_26856), .c(n_26546), .o(n_26890) );
ao12f80 g746045 ( .a(n_35161), .b(n_35190), .c(n_35160), .o(n_35259) );
no02f80 g736507 ( .a(n_43665), .b(n_43234), .o(n_43675) );
oa12f80 g762765 ( .a(n_18142), .b(n_18158), .c(n_18141), .o(n_18422) );
na02f80 g766179 ( .a(n_14511), .b(n_14510), .o(n_14545) );
in01f80 FE_RC_2726_0 ( .a(n_18356), .o(FE_RN_1153_0) );
oa22f80 FE_RC_788_0 ( .a(n_11802), .b(n_12023), .c(n_11801), .d(n_11988), .o(n_12211) );
na02f80 g745299 ( .a(n_36021), .b(n_35932), .o(n_36052) );
na02f80 g750062 ( .a(n_29869), .b(n_29111), .o(n_30053) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_27_ ( .ck(newNet_2169), .d(n_1009), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_27_) );
in01f80 g742724 ( .a(n_37849), .o(n_37352) );
no02f80 g754964 ( .a(n_25868), .b(n_25839), .o(n_25840) );
na02f80 g768742 ( .a(n_12128), .b(n_12127), .o(n_12273) );
no02f80 g764898 ( .a(n_15680), .b(n_15677), .o(n_15888) );
in01f80 fopt783144 ( .a(n_1282), .o(n_44650) );
na02f80 g739130 ( .a(n_40976), .b(n_40831), .o(n_40995) );
na02f80 g755844 ( .a(n_24314), .b(n_24015), .o(n_24313) );
no02f80 g770877 ( .a(n_10007), .b(n_9744), .o(n_10134) );
na02f80 g747379 ( .a(FE_OCP_RBN2102_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_10_), .o(n_32665) );
in01f80 g741138 ( .a(n_39151), .o(n_39152) );
in01f80 g749785 ( .a(n_31627), .o(n_31628) );
na02f80 g775714 ( .a(n_5409), .b(n_5344), .o(n_5459) );
no02f80 g772006 ( .a(n_44511), .b(n_8811), .o(n_11041) );
na02f80 g754234 ( .a(n_26744), .b(n_26743), .o(n_26745) );
in01f80 newInst_3570 ( .a(newNet_3569), .o(newNet_3570) );
na02f80 FE_RC_2845_0 ( .a(FE_RN_1224_0), .b(n_11240), .o(n_11313) );
no02f80 g744232 ( .a(n_36816), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n_36862) );
ao12f80 g752303 ( .a(n_28050), .b(n_28457), .c(n_27949), .o(n_28479) );
in01f80 FE_RC_4193_0 ( .a(FE_RN_1719_0), .o(FE_RN_1837_0) );
in01f80 FE_OCPC1231_n_42201 ( .a(FE_OCPN1230_n_42201), .o(FE_OCPN1231_n_42201) );
in01f80 g757381 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_12_), .o(n_23106) );
no02f80 g767694 ( .a(n_13256), .b(n_13255), .o(n_13346) );
no02f80 g758128 ( .a(n_22212), .b(n_22333), .o(n_22335) );
in01f80 newInst_470 ( .a(newNet_469), .o(newNet_470) );
na02f80 g770088 ( .a(n_10672), .b(n_10357), .o(n_10732) );
in01f80 g771366 ( .a(n_9261), .o(n_9194) );
in01f80 g739306 ( .a(n_41009), .o(n_41010) );
in01f80 g755704 ( .a(n_24547), .o(n_24548) );
in01f80 g755315 ( .a(n_25685), .o(n_25547) );
na02f80 g772020 ( .a(n_44463), .b(n_9681), .o(n_9733) );
na02f80 g757241 ( .a(n_23495), .b(n_22924), .o(n_23535) );
in01f80 g778456 ( .a(n_2511), .o(n_2512) );
no02f80 g763356 ( .a(FE_OCP_RBN3213_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .o(n_17133) );
na02f80 g754108 ( .a(n_25998), .b(FE_OCPN1440_n_23339), .o(n_26064) );
in01f80 newInst_2850 ( .a(newNet_2849), .o(newNet_2850) );
in01f80 newInst_2182 ( .a(newNet_2181), .o(newNet_2182) );
na02f80 g740864 ( .a(n_39217), .b(n_39332), .o(n_39398) );
in01f80 newInst_2445 ( .a(newNet_2444), .o(newNet_2445) );
in01f80 g781308 ( .a(n_57), .o(n_102) );
no02f80 g773405 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_26_), .o(n_8742) );
no02f80 g738767 ( .a(n_41357), .b(n_40863), .o(n_41370) );
in01f80 g761639 ( .a(n_18797), .o(n_18949) );
no02f80 g768973 ( .a(n_11596), .b(n_11608), .o(n_11609) );
in01f80 FE_OCPC1496_n_26528 ( .a(FE_OCPN1495_n_26528), .o(FE_OCPN1496_n_26528) );
in01f80 FE_OCP_RBC2982_n_26767 ( .a(n_26767), .o(FE_OCP_RBN2982_n_26767) );
oa22f80 g741515 ( .a(n_38673), .b(n_38624), .c(n_38674), .d(n_38637), .o(n_38747) );
ao12f80 g736297 ( .a(n_43357), .b(n_43859), .c(n_43645), .o(n_43882) );
oa22f80 g778514 ( .a(n_2608), .b(n_2090), .c(n_2530), .d(n_2091), .o(n_2672) );
in01f80 g773328 ( .a(n_8232), .o(n_8362) );
ao12f80 g751719 ( .a(n_28147), .b(n_28322), .c(n_28187), .o(n_28373) );
in01f80 g770283 ( .a(n_10517), .o(n_10518) );
na02f80 g773204 ( .a(n_7674), .b(n_7673), .o(n_7681) );
na02f80 g744305 ( .a(n_44174), .b(n_36062), .o(n_36089) );
na02f80 g781085 ( .a(n_282), .b(state_cordic_1_), .o(n_43918) );
oa12f80 g770921 ( .a(n_9838), .b(n_10049), .c(n_9918), .o(n_10182) );
na02f80 g775655 ( .a(n_5314), .b(n_5345), .o(n_5424) );
oa12f80 g749703 ( .a(n_31540), .b(n_31481), .c(FE_OCP_RBN3011_n_31117), .o(n_31635) );
na02f80 g770906 ( .a(n_10132), .b(n_10171), .o(n_10133) );
na02f80 g764448 ( .a(n_16220), .b(FE_OCPN3775_n_14730), .o(n_16219) );
no03m80 FE_RC_624_0 ( .a(n_40986), .b(n_41293), .c(n_41294), .o(n_41314) );
no02f80 g737694 ( .a(n_42216), .b(n_41797), .o(n_42288) );
no02f80 g767559 ( .a(n_13050), .b(n_12283), .o(n_13183) );
in01f80 g765497 ( .a(n_15867), .o(n_15868) );
na02f80 g739104 ( .a(n_41002), .b(n_41001), .o(n_41003) );
na02f80 g743929 ( .a(n_35825), .b(n_44222), .o(n_35913) );
ao12f80 g779488 ( .a(n_2083), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_26_), .o(n_2090) );
in01f80 g771986 ( .a(n_9601), .o(n_9602) );
no02f80 g763033 ( .a(n_17455), .b(n_17022), .o(n_17514) );
in01f80 FE_OCP_RBC2432_n_14018 ( .a(FE_OCP_RBN2431_n_14018), .o(FE_OCP_RBN2432_n_14018) );
no02f80 g766377 ( .a(n_14278), .b(FE_OCPN3765_FE_OCP_RBN2222_n_13010), .o(n_14318) );
oa22f80 g780030 ( .a(n_1251), .b(n_1070), .c(n_1250), .d(n_1071), .o(n_1260) );
in01f80 g745263 ( .a(n_35968), .o(n_35941) );
oa22f80 g745341 ( .a(n_36049), .b(n_35525), .c(FE_OCP_RBN2994_n_35539), .d(n_36022), .o(n_36211) );
in01f80 g747452 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_30_), .o(n_32354) );
oa12f80 g764811 ( .a(n_15723), .b(n_15888), .c(n_15790), .o(n_16029) );
na02f80 g771069 ( .a(n_9715), .b(FE_OCPN903_n_44581), .o(n_9716) );
in01f80 newInst_2942 ( .a(newNet_2333), .o(newNet_2942) );
in01f80 newInst_1485 ( .a(newNet_1344), .o(newNet_1485) );
in01f80 g772202 ( .a(n_8895), .o(n_8896) );
na02f80 g775872 ( .a(n_5475), .b(n_5374), .o(n_5697) );
no02f80 g742133 ( .a(n_38266), .b(n_38276), .o(n_38309) );
in01f80 g746865 ( .a(n_33447), .o(n_33448) );
no02f80 g757403 ( .a(n_22942), .b(n_22941), .o(n_22967) );
no02f80 g755751 ( .a(n_24402), .b(n_24039), .o(n_24403) );
in01f80 newInst_570 ( .a(newNet_569), .o(newNet_570) );
in01f80 FE_RC_4056_0 ( .a(n_26401), .o(FE_RN_1764_0) );
in01f80 g776752 ( .a(n_3981), .o(n_3982) );
no02f80 g741576 ( .a(n_38629), .b(n_38630), .o(n_38666) );
in01f80 g746584 ( .a(n_34885), .o(n_34886) );
in01f80 newInst_2727 ( .a(newNet_408), .o(newNet_2727) );
in01f80 g742834 ( .a(n_37240), .o(n_37241) );
no02f80 g762323 ( .a(n_18160), .b(n_18159), .o(n_18185) );
in01f80 g756141 ( .a(n_24906), .o(n_24902) );
ao22s80 g742036 ( .a(FE_OCP_RBN3445_n_37945), .b(n_37364), .c(FE_OCP_RBN3442_n_37945), .d(n_37393), .o(n_38359) );
in01f80 g751293 ( .a(FE_OCPN1478_n_28775), .o(n_28776) );
in01f80 g770103 ( .a(n_10889), .o(n_10890) );
no02f80 FE_RC_2071_0 ( .a(n_24923), .b(n_24924), .o(FE_RN_706_0) );
na02f80 g759786 ( .a(n_21773), .b(n_21825), .o(n_21861) );
in01f80 newInst_1896 ( .a(newNet_1895), .o(newNet_1896) );
in01f80 FE_RC_1965_0 ( .a(n_23914), .o(FE_RN_635_0) );
no02f80 g736728 ( .a(n_43200), .b(n_43136), .o(n_43227) );
in01f80 g741265 ( .a(n_39318), .o(n_39319) );
no02f80 FE_RC_2471_0 ( .a(FE_RN_994_0), .b(FE_RN_995_0), .o(FE_RN_996_0) );
na02f80 g737745 ( .a(FE_OCPN885_n_42216), .b(n_42064), .o(n_42449) );
no02f80 g784115 ( .a(n_47176), .b(n_45858), .o(n_45865) );
in01f80 newInst_1424 ( .a(newNet_1423), .o(newNet_1424) );
ao12f80 g780426 ( .a(n_878), .b(n_1099), .c(FE_OFN50_n_1045), .o(n_907) );
in01f80 g748736 ( .a(n_31399), .o(n_31357) );
no02f80 g758893 ( .a(n_21609), .b(n_21462), .o(n_21703) );
no02f80 g747820 ( .a(n_33238), .b(n_33294), .o(n_33311) );
na02f80 g749605 ( .a(n_31582), .b(n_31580), .o(n_31581) );
in01f80 g764938 ( .a(n_45502), .o(n_15656) );
na02f80 g780458 ( .a(n_1098), .b(FE_OFN50_n_1045), .o(n_834) );
na02f80 FE_RC_2022_0 ( .a(FE_RN_669_0), .b(FE_RN_670_0), .o(FE_RN_671_0) );
ao12f80 FE_RC_2502_0 ( .a(FE_RN_1014_0), .b(FE_RN_1015_0), .c(n_42038), .o(n_42100) );
no02f80 g772781 ( .a(n_8097), .b(n_8096), .o(n_8098) );
no02f80 g752963 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_), .o(n_28106) );
in01f80 newInst_486 ( .a(newNet_485), .o(newNet_486) );
na02f80 g767477 ( .a(n_13225), .b(n_12321), .o(n_13338) );
na02f80 g769263 ( .a(n_11556), .b(n_10910), .o(n_11671) );
in01f80 g780760 ( .a(n_695), .o(n_550) );
no02f80 g751060 ( .a(n_30381), .b(n_29939), .o(n_30520) );
oa12f80 g772907 ( .a(n_7935), .b(n_7934), .c(n_7933), .o(n_9605) );
na02f80 g771837 ( .a(n_9650), .b(n_9735), .o(n_10351) );
in01f80 g737457 ( .a(n_42792), .o(n_42771) );
in01f80 g761349 ( .a(n_18982), .o(n_19034) );
no02f80 g744514 ( .a(n_35413), .b(n_35283), .o(n_35423) );
in01f80 g777018 ( .a(n_3875), .o(n_3876) );
in01f80 g771931 ( .a(n_9001), .o(n_9002) );
no02f80 g773190 ( .a(n_7612), .b(n_8174), .o(n_7627) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_29_ ( .ck(newNet_3123), .d(n_40593), .o(delay_add_ln22_unr27_stage10_stallmux_q_29_) );
ao12f80 g784435 ( .a(n_46226), .b(n_46197), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n_46247) );
in01f80 FE_RC_3227_0 ( .a(n_8709), .o(FE_RN_1430_0) );
na02f80 g743546 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n_36475) );
in01f80 g769701 ( .a(n_11331), .o(n_11332) );
no02f80 g738702 ( .a(n_41483), .b(n_41492), .o(n_41571) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_25_ ( .ck(newNet_2842), .d(n_12068), .o(delay_add_ln22_unr8_stage4_stallmux_q_25_) );
na02f80 g759354 ( .a(n_21006), .b(n_45091), .o(n_21077) );
in01f80 g736314 ( .a(n_43876), .o(n_43877) );
oa12f80 g758780 ( .a(n_22180), .b(n_22209), .c(n_22179), .o(n_22244) );
in01f80 FE_OCP_RBC2260_n_18899 ( .a(n_18899), .o(FE_OCP_RBN2260_n_18899) );
in01f80 FE_OCPC1408_n_672 ( .a(FE_OCPN1407_n_672), .o(FE_OCPN1408_n_672) );
na02f80 g771356 ( .a(FE_OCP_RBN3569_n_9188), .b(n_8309), .o(n_9295) );
in01f80 newInst_1068 ( .a(newNet_1067), .o(newNet_1068) );
no02f80 g764274 ( .a(n_16297), .b(n_16337), .o(n_16471) );
no02f80 g743915 ( .a(n_36100), .b(n_36141), .o(n_36246) );
in01f80 g746542 ( .a(n_34525), .o(n_34526) );
no02f80 g743133 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .o(n_37036) );
na02f80 g773860 ( .a(n_7127), .b(n_7010), .o(n_7125) );
no02f80 g740680 ( .a(n_39552), .b(n_45841), .o(n_39589) );
no02f80 g742674 ( .a(n_37457), .b(n_37456), .o(n_37458) );
in01f80 newInst_3586 ( .a(newNet_3585), .o(newNet_3586) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_12_ ( .ck(newNet_267), .d(n_46161), .o(delay_xor_ln22_unr6_stage3_stallmux_q_12_) );
na02f80 g769785 ( .a(n_11208), .b(n_10982), .o(n_11238) );
no02f80 g742242 ( .a(FE_OCP_RBN2240_n_44881), .b(n_37719), .o(n_38213) );
no02f80 g765005 ( .a(n_15644), .b(n_15643), .o(n_15581) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_10_ ( .ck(newNet_1042), .d(n_17654), .o(delay_xor_ln21_unr12_stage5_stallmux_q_10_) );
in01f80 g746675 ( .a(n_34612), .o(n_34666) );
in01f80 g756196 ( .a(n_24791), .o(n_24792) );
no02f80 g743009 ( .a(n_37147), .b(n_37091), .o(n_37157) );
in01f80 g775867 ( .a(n_5249), .o(n_5250) );
in01f80 g749738 ( .a(n_31292), .o(n_31349) );
in01f80 newInst_2414 ( .a(newNet_2404), .o(newNet_2414) );
oa22f80 FE_RC_4125_0 ( .a(n_20226), .b(n_20210), .c(n_20209), .d(n_20241), .o(n_20336) );
na02f80 g755899 ( .a(n_24229), .b(n_24228), .o(n_24322) );
in01f80 g758315 ( .a(n_22149), .o(n_22333) );
in01f80 g779149 ( .a(n_2025), .o(n_2003) );
no02f80 g766991 ( .a(n_13770), .b(n_13769), .o(n_13771) );
no02f80 g753936 ( .a(n_26158), .b(n_26206), .o(n_26262) );
na02f80 g746006 ( .a(n_34010), .b(n_34009), .o(n_34063) );
oa22f80 FE_RC_3438_0 ( .a(n_22961), .b(n_22902), .c(n_20252), .d(n_22862), .o(n_22962) );
in01f80 newInst_839 ( .a(newNet_183), .o(newNet_839) );
oa12f80 g752599 ( .a(n_27436), .b(n_27568), .c(n_27277), .o(n_27628) );
na02f80 g758056 ( .a(n_23052), .b(n_23051), .o(n_23642) );
no02f80 g762313 ( .a(n_18056), .b(n_18055), .o(n_18078) );
in01f80 FE_OCP_RBC2509_n_13896 ( .a(FE_OCP_RBN2508_n_13896), .o(FE_OCP_RBN2509_n_13896) );
no02f80 g754955 ( .a(n_25481), .b(n_24635), .o(n_25588) );
no02f80 g761970 ( .a(n_18963), .b(n_18931), .o(n_18992) );
ao12f80 g745092 ( .a(n_34489), .b(n_34661), .c(n_34368), .o(n_34768) );
na02f80 g764104 ( .a(n_16517), .b(n_16369), .o(n_16569) );
no02f80 g755555 ( .a(n_24617), .b(n_24600), .o(n_24718) );
in01f80 g771074 ( .a(n_9928), .o(n_9888) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_16_ ( .ck(newNet_3158), .d(n_40457), .o(delay_add_ln22_unr27_stage10_stallmux_q_16_) );
na02f80 g737438 ( .a(n_42716), .b(n_42425), .o(n_42733) );
na02f80 g741543 ( .a(n_38655), .b(n_38652), .o(n_38656) );
in01f80 FE_RC_2696_0 ( .a(n_8710), .o(FE_RN_1130_0) );
no02f80 g768586 ( .a(n_12233), .b(n_11860), .o(n_12267) );
in01f80 g757731 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n_22562) );
no02f80 FE_RC_3526_0 ( .a(FE_RN_1524_0), .b(n_27476), .o(n_27535) );
no02f80 g740751 ( .a(n_39356), .b(n_39258), .o(n_39416) );
na02f80 g784138 ( .a(n_45879), .b(n_45884), .o(n_45889) );
na02f80 g743468 ( .a(n_36520), .b(n_36750), .o(n_36521) );
ao12f80 g778293 ( .a(n_2525), .b(n_2524), .c(n_2523), .o(n_2674) );
na02f80 g771620 ( .a(n_9201), .b(n_9071), .o(n_9242) );
no02f80 g740063 ( .a(n_40117), .b(n_40116), .o(n_40143) );
no02f80 g768109 ( .a(n_12698), .b(n_12415), .o(n_12761) );
in01f80 FE_RC_125_0 ( .a(n_11769), .o(FE_RN_30_0) );
na02f80 g759495 ( .a(n_20959), .b(n_20957), .o(n_21054) );
no02f80 g765526 ( .a(n_15599), .b(n_15086), .o(n_15834) );
ao12f80 g768702 ( .a(n_12148), .b(n_45659), .c(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .o(n_12238) );
no02f80 g748410 ( .a(FE_OCPN1052_n_31674), .b(n_30643), .o(n_31787) );
in01f80 FE_OCPC1743_n_24962 ( .a(n_24962), .o(FE_OCPN1743_n_24962) );
no02f80 g737523 ( .a(n_42532), .b(n_42531), .o(n_42533) );
no02f80 g754074 ( .a(n_26067), .b(n_26093), .o(n_26167) );
in01f80 g758793 ( .a(n_21617), .o(n_21654) );
oa22f80 FE_RC_1707_0 ( .a(n_22961), .b(n_46965), .c(n_22580), .d(n_22594), .o(n_22671) );
in01f80 g779516 ( .a(n_1567), .o(n_1568) );
in01f80 g769292 ( .a(n_11560), .o(n_11684) );
in01f80 g772944 ( .a(n_7894), .o(n_7895) );
oa12f80 g749671 ( .a(n_30026), .b(n_30057), .c(n_30025), .o(n_31719) );
in01f80 FE_RC_3746_0 ( .a(FE_RN_1643_0), .o(FE_RN_1644_0) );
oa12f80 g752250 ( .a(n_28212), .b(FE_OCP_RBN2179_FE_RN_526_0), .c(n_28259), .o(n_28559) );
na02f80 g763693 ( .a(n_16749), .b(n_16726), .o(n_16784) );
no02f80 g743437 ( .a(n_36551), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36586) );
in01f80 newInst_3591 ( .a(newNet_1098), .o(newNet_3591) );
in01f80 g756536 ( .a(n_23586), .o(n_23639) );
ao12f80 g762842 ( .a(n_17740), .b(n_17839), .c(n_17791), .o(n_17843) );
no02f80 g753679 ( .a(n_26586), .b(n_26533), .o(n_26674) );
na02f80 g736736 ( .a(n_43306), .b(n_43324), .o(n_43360) );
oa12f80 g768100 ( .a(n_12598), .b(n_12597), .c(n_12596), .o(n_13800) );
no02f80 g769837 ( .a(n_46987), .b(n_9682), .o(n_11283) );
in01f80 newInst_2874 ( .a(newNet_71), .o(newNet_2874) );
na02f80 g764679 ( .a(n_15706), .b(n_14524), .o(n_15743) );
na02f80 g764361 ( .a(n_16288), .b(n_16157), .o(n_16289) );
na02f80 g772016 ( .a(FE_OCP_RBN3644_n_44490), .b(n_9768), .o(n_9874) );
ao12f80 g767546 ( .a(n_13217), .b(n_13216), .c(n_13215), .o(n_13324) );
no02f80 g757006 ( .a(n_23305), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .o(n_23371) );
in01f80 g751016 ( .a(n_30067), .o(n_30127) );
in01f80 newInst_3685 ( .a(newNet_3576), .o(newNet_3685) );
in01f80 fopt783526 ( .a(n_45139), .o(n_45137) );
oa22f80 g780010 ( .a(n_1270), .b(n_1044), .c(n_1271), .d(n_1043), .o(n_1275) );
in01f80 g738840 ( .a(n_41313), .o(n_41325) );
na02f80 g763163 ( .a(n_17281), .b(n_17274), .o(n_17405) );
na02f80 g760354 ( .a(n_20782), .b(n_20781), .o(n_20783) );
na02f80 g773148 ( .a(n_7674), .b(n_7163), .o(n_7716) );
oa12f80 g736477 ( .a(n_323), .b(n_43672), .c(FE_OFN3_n_43918), .o(n_43707) );
no02f80 g771148 ( .a(n_9839), .b(n_9918), .o(n_10004) );
no02f80 g745311 ( .a(n_34386), .b(n_34385), .o(n_34387) );
no03m80 g766843 ( .a(n_13939), .b(n_13943), .c(n_13821), .o(n_13940) );
in01f80 g779465 ( .a(n_1854), .o(n_1855) );
no02f80 g771411 ( .a(n_9562), .b(n_9608), .o(n_9785) );
in01f80 g776601 ( .a(n_4233), .o(n_4234) );
na02f80 g750077 ( .a(n_29869), .b(n_30214), .o(n_30215) );
no02f80 g760300 ( .a(n_20834), .b(n_19933), .o(n_20953) );
in01f80 newInst_1459 ( .a(newNet_379), .o(newNet_1459) );
in01f80 newInst_2760 ( .a(newNet_1419), .o(newNet_2760) );
ao12f80 g741803 ( .a(n_38307), .b(n_38388), .c(n_38347), .o(n_38491) );
in01f80 newInst_3290 ( .a(newNet_3289), .o(newNet_3290) );
in01f80 newInst_1019 ( .a(newNet_1018), .o(newNet_1019) );
in01f80 g773842 ( .a(n_7163), .o(n_7164) );
na02f80 g759180 ( .a(n_21157), .b(n_45023), .o(n_21317) );
in01f80 g756129 ( .a(n_25188), .o(n_25160) );
no02f80 g773099 ( .a(n_7996), .b(n_7995), .o(n_8588) );
in01f80 g753457 ( .a(n_26980), .o(n_26981) );
na02f80 g743267 ( .a(n_36761), .b(n_36692), .o(n_36783) );
no02f80 g754726 ( .a(FE_OCP_RBN2966_n_26231), .b(n_26542), .o(n_26636) );
na02f80 g751595 ( .a(n_28597), .b(n_28606), .o(n_28598) );
in01f80 g738534 ( .a(n_41408), .o(n_41409) );
na02f80 g751961 ( .a(n_28919), .b(n_29067), .o(n_29305) );
in01f80 newInst_3474 ( .a(newNet_3473), .o(newNet_3474) );
no02f80 g746739 ( .a(n_33037), .b(n_33023), .o(n_33067) );
ao12f80 g771097 ( .a(n_9721), .b(n_9921), .c(n_9786), .o(n_10045) );
no02f80 g771937 ( .a(n_8700), .b(n_8699), .o(n_8701) );
no02f80 g749880 ( .a(n_29900), .b(n_29896), .o(n_29967) );
no02f80 g746003 ( .a(n_33979), .b(n_34032), .o(n_34061) );
no02f80 g749039 ( .a(n_31094), .b(n_31093), .o(n_31149) );
na02f80 g750429 ( .a(n_29553), .b(n_25859), .o(n_29554) );
na02f80 FE_RC_915_0 ( .a(n_31029), .b(n_30939), .o(FE_RN_271_0) );
ao12f80 g779219 ( .a(n_1819), .b(n_1818), .c(n_1817), .o(n_2255) );
na02f80 g740197 ( .a(FE_OCP_RBN3722_n_39913), .b(n_40177), .o(n_40291) );
no02f80 g778142 ( .a(n_2930), .b(n_2929), .o(n_2964) );
oa12f80 g751409 ( .a(n_28455), .b(n_28477), .c(n_28454), .o(n_29765) );
in01f80 g775678 ( .a(n_5611), .o(n_5612) );
na02f80 g746083 ( .a(n_33937), .b(n_33448), .o(n_33955) );
no02f80 g738598 ( .a(n_41365), .b(n_40930), .o(n_41388) );
na02f80 g743750 ( .a(n_37305), .b(n_37304), .o(n_37307) );
ao12f80 g742616 ( .a(n_37425), .b(n_37424), .c(n_37423), .o(n_38298) );
in01f80 FE_OCP_RBC2210_n_37694 ( .a(n_37694), .o(FE_OCP_RBN2210_n_37694) );
oa22f80 FE_RC_3648_0 ( .a(n_17321), .b(n_17514), .c(n_17322), .d(n_17493), .o(n_17686) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_2_ ( .ck(newNet_1010), .d(n_16730), .o(delay_xor_ln21_unr12_stage5_stallmux_q_2_) );
na02f80 g740365 ( .a(n_39787), .b(n_39810), .o(n_39811) );
oa22f80 FE_RC_3802_0 ( .a(FE_OCP_RBN1176_n_18981), .b(n_19249), .c(FE_OCP_RBN1177_n_18981), .d(n_19271), .o(n_19437) );
in01f80 FE_OCP_RBC2144_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2142_FE_OCPN861_n_45450), .o(FE_OCP_RBN2144_FE_OCPN861_n_45450) );
na02f80 g748794 ( .a(n_32455), .b(n_32454), .o(n_32456) );
no02f80 g753892 ( .a(n_26279), .b(n_26362), .o(n_26426) );
in01f80 g757935 ( .a(n_22926), .o(n_22884) );
in01f80 newInst_2105 ( .a(newNet_2104), .o(newNet_2105) );
in01f80 newInst_4 ( .a(newNet_3), .o(newNet_4) );
oa12f80 g738302 ( .a(n_41485), .b(n_41757), .c(n_41593), .o(n_41865) );
no02f80 g752931 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_), .o(n_28108) );
no02f80 g761814 ( .a(n_18379), .b(n_18377), .o(n_18378) );
in01f80 g768082 ( .a(n_13103), .o(n_13104) );
in01f80 g752856 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_), .o(n_28342) );
no02f80 g767550 ( .a(n_12875), .b(n_12947), .o(n_12948) );
na02f80 g742995 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_7_), .b(delay_add_ln22_unr23_stage9_stallmux_q_7_), .o(n_36964) );
in01f80 newInst_1536 ( .a(newNet_1535), .o(newNet_1536) );
no02f80 g744329 ( .a(n_44180), .b(n_35195), .o(n_36063) );
in01f80 g778578 ( .a(n_2485), .o(n_2486) );
no02f80 g756753 ( .a(n_23870), .b(n_23671), .o(n_23939) );
in01f80 g779436 ( .a(n_1829), .o(n_1830) );
in01f80 FE_OCPC1777_n_37744 ( .a(n_37744), .o(FE_OCPN1777_n_37744) );
in01f80 FE_OCPC1502_n_20723 ( .a(FE_OCPN1501_n_20723), .o(FE_OCPN1502_n_20723) );
no02f80 g762038 ( .a(n_18780), .b(n_18779), .o(n_18781) );
na02f80 g777001 ( .a(n_3960), .b(n_4098), .o(n_4143) );
in01f80 g746262 ( .a(n_33687), .o(n_33688) );
na02f80 g750549 ( .a(n_29422), .b(n_30111), .o(n_29454) );
in01f80 g775675 ( .a(n_5620), .o(n_5621) );
in01f80 FE_RC_2016_0 ( .a(n_13419), .o(FE_RN_667_0) );
ao12f80 g753789 ( .a(n_26861), .b(n_27067), .c(n_26547), .o(n_27095) );
no02f80 g750782 ( .a(n_29145), .b(n_28679), .o(n_29195) );
in01f80 g765813 ( .a(n_15091), .o(n_15331) );
ao12f80 g767083 ( .a(n_13719), .b(n_13718), .c(n_13717), .o(n_14257) );
oa22f80 g784146 ( .a(n_36898), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .c(n_45890), .d(n_37023), .o(n_45896) );
in01f80 newInst_1305 ( .a(newNet_676), .o(newNet_1305) );
na02f80 g768756 ( .a(n_12174), .b(n_12173), .o(n_12175) );
ao12f80 g751363 ( .a(n_28908), .b(n_29361), .c(n_28991), .o(n_29463) );
in01f80 newInst_1915 ( .a(newNet_1914), .o(newNet_1915) );
oa12f80 g741874 ( .a(n_38348), .b(n_38244), .c(n_38301), .o(n_38416) );
oa12f80 g744504 ( .a(n_36685), .b(n_36682), .c(n_36049), .o(n_36728) );
in01f80 g763341 ( .a(n_17376), .o(n_17377) );
ao12f80 g745060 ( .a(n_35718), .b(n_36232), .c(n_35769), .o(n_36315) );
in01f80 FE_OCP_RBC2307_n_24288 ( .a(n_24288), .o(FE_OCP_RBN2307_n_24288) );
no02f80 g743749 ( .a(n_37292), .b(n_37246), .o(n_37308) );
no02f80 g766882 ( .a(n_14389), .b(n_14350), .o(n_15244) );
na02f80 g749945 ( .a(n_30349), .b(n_30371), .o(n_30369) );
no02f80 g770038 ( .a(n_10922), .b(FE_OCP_RBN3643_n_44490), .o(n_10955) );
in01f80 g754010 ( .a(n_26158), .o(n_26182) );
na02f80 g765316 ( .a(FE_OCP_RBN3507_n_13860), .b(FE_OCP_RBN2681_n_15048), .o(n_15273) );
no02f80 g774339 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_18_), .o(n_7121) );
na02f80 g750727 ( .a(n_29196), .b(n_28769), .o(n_29198) );
in01f80 g780907 ( .a(n_478), .o(n_472) );
na02f80 g743815 ( .a(n_46251), .b(n_46202), .o(n_37202) );
in01f80 g765630 ( .a(n_15047), .o(n_15116) );
in01f80 g759618 ( .a(n_20872), .o(n_20873) );
no02f80 g780564 ( .a(n_890), .b(n_661), .o(n_1027) );
oa22f80 g746226 ( .a(n_33844), .b(n_33768), .c(n_33706), .d(n_32574), .o(n_35106) );
in01f80 g752923 ( .a(n_27813), .o(n_27789) );
no02f80 g771828 ( .a(n_10037), .b(n_10081), .o(n_10082) );
na02f80 g751343 ( .a(n_29489), .b(n_29048), .o(n_29601) );
no02f80 g741564 ( .a(n_38646), .b(n_38632), .o(n_38676) );
no02f80 g775816 ( .a(n_5233), .b(n_5200), .o(n_5304) );
in01f80 g737425 ( .a(n_42782), .o(n_42751) );
na02f80 g745322 ( .a(n_35679), .b(n_35678), .o(n_35680) );
in01f80 g740924 ( .a(n_39368), .o(n_39369) );
in01f80 g771980 ( .a(n_9516), .o(n_9517) );
na02f80 g762020 ( .a(n_18390), .b(n_18460), .o(n_18506) );
in01f80 newInst_1043 ( .a(newNet_36), .o(newNet_1043) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_13_ ( .ck(newNet_1425), .d(n_36528), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_) );
in01f80 g759312 ( .a(n_21259), .o(n_21260) );
na02f80 g743515 ( .a(n_36534), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36562) );
na02f80 g760774 ( .a(n_19558), .b(n_19528), .o(n_19597) );
oa22f80 FE_RC_779_0 ( .a(n_8366), .b(FE_OCP_RBN2513_n_8533), .c(n_8348), .d(n_8533), .o(n_8677) );
in01f80 g761958 ( .a(n_18397), .o(n_18553) );
no02f80 g739217 ( .a(n_40786), .b(n_40785), .o(n_40827) );
in01f80 g767967 ( .a(n_13274), .o(n_13275) );
no02f80 g742738 ( .a(n_37442), .b(n_37441), .o(n_37443) );
in01f80 g753074 ( .a(n_27923), .o(n_27733) );
no02f80 g778341 ( .a(n_2495), .b(n_2494), .o(n_2526) );
in01f80 g740774 ( .a(n_46950), .o(n_39548) );
in01f80 FE_OCP_RBC2206_n_12907 ( .a(n_12907), .o(FE_OCP_RBN2206_n_12907) );
na02f80 g739334 ( .a(n_45180), .b(n_40695), .o(n_40732) );
no02f80 g767809 ( .a(n_12873), .b(n_12918), .o(n_12951) );
na02f80 g742440 ( .a(n_37657), .b(n_36947), .o(n_37737) );
no02f80 g762788 ( .a(n_17887), .b(n_17886), .o(n_17912) );
in01f80 g745365 ( .a(n_35849), .o(n_35938) );
in01f80 newInst_2639 ( .a(newNet_2638), .o(newNet_2639) );
oa22f80 g752448 ( .a(n_27610), .b(n_27487), .c(n_27624), .d(n_27486), .o(n_27720) );
ao12f80 g751366 ( .a(n_28515), .b(n_28536), .c(n_28514), .o(n_28582) );
in01f80 g781302 ( .a(n_44), .o(n_45) );
in01f80 newInst_395 ( .a(newNet_394), .o(newNet_395) );
in01f80 g774359 ( .a(n_6985), .o(n_6986) );
no02f80 g761134 ( .a(n_19088), .b(n_18358), .o(n_19116) );
in01f80 g752138 ( .a(n_28139), .o(n_28140) );
no02f80 g767954 ( .a(n_12749), .b(n_12748), .o(n_12750) );
na02f80 g779318 ( .a(n_1675), .b(n_1402), .o(n_1712) );
na02f80 g751326 ( .a(n_29537), .b(n_29536), .o(n_29538) );
no02f80 g751913 ( .a(n_28902), .b(n_28923), .o(n_28903) );
in01f80 newInst_596 ( .a(newNet_595), .o(newNet_596) );
in01f80 g754759 ( .a(n_26132), .o(n_26133) );
na02f80 FE_RC_3713_0 ( .a(FE_RN_636_0), .b(FE_RN_1633_0), .o(n_24436) );
na02f80 g770802 ( .a(n_10218), .b(n_10217), .o(n_10219) );
ms00f80 cos_out_reg_13_ ( .ck(newNet_3746), .d(n_43796), .o(cos_out_13) );
na02f80 g738510 ( .a(FE_OCPN952_n_41540), .b(n_41576), .o(n_41814) );
no02f80 g770137 ( .a(n_10730), .b(n_44490), .o(n_10762) );
in01f80 g737131 ( .a(n_43030), .o(n_43171) );
in01f80 g771555 ( .a(n_9506), .o(n_9606) );
na03f80 FE_RC_1701_0 ( .a(n_24422), .b(n_24574), .c(FE_OCP_RBN1162_n_24701), .o(n_46963) );
na02f80 g751440 ( .a(n_28528), .b(n_28493), .o(n_28529) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_28_ ( .ck(newNet_2164), .d(n_902), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_28_) );
in01f80 g739313 ( .a(n_40887), .o(n_40763) );
in01f80 g760070 ( .a(n_20273), .o(n_20295) );
na02f80 g746346 ( .a(n_33610), .b(n_33609), .o(n_33611) );
in01f80 g766645 ( .a(n_13981), .o(n_13982) );
ao12f80 g750287 ( .a(n_29734), .b(n_29733), .c(n_29735), .o(n_31206) );
na02f80 g770587 ( .a(FE_OCP_RBN2794_n_10106), .b(FE_OCP_RBN3570_n_9188), .o(n_10359) );
no02f80 g738332 ( .a(n_41647), .b(n_41624), .o(n_41712) );
na02f80 g764266 ( .a(n_16432), .b(n_16393), .o(n_16460) );
ao12f80 g751307 ( .a(n_29333), .b(n_29599), .c(n_29043), .o(n_29693) );
ao22s80 g773807 ( .a(n_7153), .b(n_7025), .c(n_7131), .d(n_7024), .o(n_7201) );
no02f80 g738760 ( .a(n_41382), .b(n_41063), .o(n_41683) );
na02f80 g761156 ( .a(FE_OCP_RBN1352_n_19148), .b(FE_OCP_RBN1176_n_18981), .o(n_19236) );
ao12f80 g779474 ( .a(n_2073), .b(n_1800), .c(delay_xor_ln22_unr3_stage2_stallmux_q_25_), .o(n_2496) );
no02f80 g770452 ( .a(n_10401), .b(n_44464), .o(n_10442) );
ao12f80 g749581 ( .a(n_30449), .b(n_30448), .c(n_30447), .o(n_30527) );
in01f80 FE_RC_3545_0 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_), .o(FE_RN_1536_0) );
in01f80 g752635 ( .a(n_27565), .o(n_27566) );
in01f80 g738820 ( .a(n_41353), .o(n_41344) );
in01f80 g745054 ( .a(n_34828), .o(n_35861) );
na02f80 g767027 ( .a(n_14758), .b(n_14168), .o(n_14427) );
in01f80 newInst_464 ( .a(newNet_195), .o(newNet_464) );
in01f80 g764556 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_9_), .o(n_17886) );
na02f80 g766053 ( .a(n_14582), .b(n_14473), .o(n_14615) );
na02f80 g775565 ( .a(n_5515), .b(n_5513), .o(n_5608) );
in01f80 FE_OCPC1438_FE_OCP_RBN1330_n_18866 ( .a(FE_OCPN1437_FE_OCP_RBN1330_n_18866), .o(FE_OCPN1438_FE_OCP_RBN1330_n_18866) );
no02f80 g758845 ( .a(n_21508), .b(n_21507), .o(n_21552) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_17_ ( .ck(newNet_650), .d(n_46348), .o(delay_xor_ln21_unr9_stage4_stallmux_q_17_) );
no02f80 g756240 ( .a(n_24070), .b(n_22089), .o(n_24099) );
no02f80 g776574 ( .a(n_4389), .b(n_3959), .o(n_4449) );
in01f80 FE_OCP_RBC3022_n_39942 ( .a(n_39942), .o(FE_OCP_RBN3022_n_39942) );
in01f80 FE_OCP_RBC1203_n_26121 ( .a(n_26121), .o(FE_OCP_RBN1203_n_26121) );
in01f80 FE_OCP_RBC3371_n_27970 ( .a(n_27970), .o(FE_OCP_RBN3371_n_27970) );
na02f80 g756716 ( .a(n_23480), .b(n_23503), .o(n_23794) );
in01f80 g760467 ( .a(n_20046), .o(n_20047) );
in01f80 newInst_1481 ( .a(newNet_1480), .o(newNet_1481) );
na02f80 FE_RC_3478_0 ( .a(n_39980), .b(n_40013), .o(FE_RN_1495_0) );
in01f80 g773785 ( .a(n_7157), .o(n_7158) );
in01f80 g741967 ( .a(n_38116), .o(n_38117) );
na02f80 g772934 ( .a(n_7934), .b(n_7933), .o(n_7935) );
no02f80 g759461 ( .a(n_20879), .b(n_20966), .o(n_21036) );
in01f80 g780461 ( .a(n_815), .o(n_847) );
no02f80 g757608 ( .a(n_22601), .b(n_22473), .o(n_22686) );
ao12f80 g784609 ( .a(n_42930), .b(n_42914), .c(n_42610), .o(n_46937) );
oa12f80 g742452 ( .a(n_37715), .b(n_37687), .c(n_37716), .o(n_37764) );
in01f80 g776233 ( .a(n_4602), .o(n_4603) );
in01f80 newInst_862 ( .a(newNet_861), .o(newNet_862) );
oa22f80 FE_RC_2681_0 ( .a(n_2998), .b(n_4057), .c(n_2997), .d(n_4131), .o(n_4238) );
na02f80 g737881 ( .a(n_42201), .b(n_42104), .o(n_42363) );
in01f80 g755041 ( .a(n_25355), .o(n_25356) );
na02f80 g774491 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_), .o(n_6737) );
na02f80 FE_RC_627_0 ( .a(FE_RN_192_0), .b(FE_RN_193_0), .o(FE_RN_194_0) );
oa12f80 g739739 ( .a(n_40399), .b(n_40513), .c(n_40130), .o(n_40540) );
na02f80 g754686 ( .a(FE_OCP_RBN2959_n_26231), .b(n_26544), .o(n_26606) );
na02f80 g767987 ( .a(n_13077), .b(n_13031), .o(n_13651) );
in01f80 newInst_1403 ( .a(newNet_982), .o(newNet_1403) );
na02f80 g746136 ( .a(n_35111), .b(n_35110), .o(n_35112) );
ao22s80 g742961 ( .a(n_37082), .b(n_36994), .c(n_46256), .d(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n_37056) );
in01f80 newInst_1428 ( .a(newNet_833), .o(newNet_1428) );
no02f80 g736755 ( .a(n_43205), .b(n_43223), .o(n_43274) );
in01f80 g741261 ( .a(n_39199), .o(n_39200) );
no02f80 g764264 ( .a(n_16438), .b(n_16272), .o(n_16439) );
na02f80 g774718 ( .a(n_6298), .b(n_6288), .o(n_6331) );
ao12f80 g741218 ( .a(n_38927), .b(FE_OCP_RBN2550_n_44944), .c(n_38890), .o(n_39269) );
oa22f80 g741820 ( .a(n_38368), .b(n_38376), .c(n_38285), .d(n_38377), .o(n_38908) );
na02f80 g772649 ( .a(n_8368), .b(n_8364), .o(n_8393) );
ao12f80 g760895 ( .a(n_19458), .b(n_19457), .c(n_19456), .o(n_21212) );
in01f80 g753168 ( .a(n_27521), .o(n_27522) );
na02f80 g763676 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_), .o(n_17610) );
na02f80 g773065 ( .a(n_8059), .b(n_8018), .o(n_8060) );
na02f80 g756031 ( .a(n_24998), .b(n_25090), .o(n_25030) );
na02f80 FE_RC_2357_0 ( .a(n_18722), .b(n_18810), .o(FE_RN_909_0) );
in01f80 g739711 ( .a(n_40515), .o(n_40516) );
no02f80 g779795 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_13_), .o(n_1484) );
in01f80 FE_OCP_RBC3066_n_36547 ( .a(n_36547), .o(FE_OCP_RBN3066_n_36547) );
no02f80 g748818 ( .a(n_32483), .b(n_32404), .o(n_32763) );
in01f80 g777102 ( .a(n_3760), .o(n_3778) );
no02f80 g755344 ( .a(n_25410), .b(n_25142), .o(n_25472) );
in01f80 FE_OCP_RBC2613_n_9075 ( .a(n_9075), .o(FE_OCP_RBN2613_n_9075) );
no02f80 g780996 ( .a(n_283), .b(n_129), .o(n_354) );
na02f80 g751606 ( .a(FE_OCPN1032_n_28448), .b(n_28424), .o(n_28463) );
ao12f80 g779454 ( .a(n_1797), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .o(n_2050) );
in01f80 newInst_2462 ( .a(newNet_2461), .o(newNet_2462) );
no02f80 g741299 ( .a(n_44955), .b(n_38892), .o(n_38925) );
in01f80 newInst_2572 ( .a(newNet_2571), .o(newNet_2572) );
na02f80 g737902 ( .a(n_42201), .b(n_41868), .o(n_42225) );
na02f80 g762792 ( .a(n_18156), .b(n_17614), .o(n_18197) );
ao12f80 g776867 ( .a(n_3918), .b(n_3955), .c(n_3753), .o(n_4026) );
na02f80 g750365 ( .a(n_29628), .b(FE_OCPN1406_n_25859), .o(n_29671) );
no02f80 FE_RC_1219_0 ( .a(FE_RN_366_0), .b(FE_RN_367_0), .o(FE_RN_368_0) );
no02f80 g744893 ( .a(n_35046), .b(n_30588), .o(n_35133) );
in01f80 newInst_3495 ( .a(newNet_898), .o(newNet_3495) );
oa12f80 g767319 ( .a(n_13347), .b(n_13636), .c(n_13316), .o(n_13697) );
oa12f80 g753610 ( .a(n_26595), .b(n_26594), .c(n_26599), .o(n_26668) );
in01f80 g764519 ( .a(n_16053), .o(n_16052) );
no02f80 g763381 ( .a(FE_OCP_RBN3724_n_16975), .b(FE_OCPN3789_n_15708), .o(n_17325) );
na02f80 g744798 ( .a(n_35097), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35200) );
no02f80 FE_RC_2724_0 ( .a(n_8332), .b(FE_RN_1151_0), .o(FE_RN_1152_0) );
na02f80 g760135 ( .a(n_20456), .b(FE_OCP_RBN1703_n_19560), .o(n_20750) );
na02f80 g760198 ( .a(FE_OCPN1261_n_20242), .b(n_20265), .o(n_20626) );
no02f80 g770326 ( .a(n_10537), .b(n_44463), .o(n_10696) );
in01f80 g759385 ( .a(n_20804), .o(n_20805) );
in01f80 newInst_3096 ( .a(newNet_3095), .o(newNet_3096) );
na02f80 g751832 ( .a(n_28207), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_7_), .o(n_28285) );
oa22f80 g773886 ( .a(n_7008), .b(n_7004), .c(n_7009), .d(n_7055), .o(n_7973) );
in01f80 FE_OCP_RBC3700_n_43015 ( .a(FE_OCP_RBN3699_n_43015), .o(FE_OCP_RBN3700_n_43015) );
na02f80 g738407 ( .a(n_41787), .b(n_41825), .o(n_41887) );
no02f80 g767414 ( .a(n_13401), .b(n_13400), .o(n_13402) );
na03f80 g746472 ( .a(n_33274), .b(n_33273), .c(n_32944), .o(n_33275) );
oa22f80 FE_RC_3233_0 ( .a(n_19419), .b(FE_RN_652_0), .c(FE_OCP_DRV_N1556_n_19384), .d(FE_RN_653_0), .o(n_19555) );
no02f80 g745217 ( .a(n_36226), .b(n_35809), .o(n_35810) );
ao22s80 g779355 ( .a(n_1604), .b(n_1633), .c(n_1662), .d(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n_1708) );
in01f80 newInst_1102 ( .a(newNet_1101), .o(newNet_1102) );
in01f80 g774367 ( .a(n_7097), .o(n_7098) );
na02f80 g751470 ( .a(n_28426), .b(n_28425), .o(n_28427) );
in01f80 g736794 ( .a(n_43554), .o(n_43555) );
na02f80 g780520 ( .a(n_794), .b(n_841), .o(n_1212) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_3_ ( .ck(newNet_3595), .d(n_15303), .o(delay_add_ln22_unr11_stage5_stallmux_q_3_) );
in01f80 FE_RC_3856_0 ( .a(n_45024), .o(FE_RN_1683_0) );
in01f80 newInst_2368 ( .a(newNet_2367), .o(newNet_2368) );
in01f80 g741736 ( .a(n_38531), .o(n_38532) );
ao12f80 g764121 ( .a(n_16134), .b(n_16930), .c(n_16261), .o(n_16960) );
in01f80 newInst_3046 ( .a(newNet_3045), .o(newNet_3046) );
no02f80 FE_RC_1050_0 ( .a(n_14563), .b(n_15287), .o(FE_RN_307_0) );
in01f80 g740204 ( .a(n_40016), .o(n_39976) );
in01f80 FE_RC_2299_0 ( .a(n_25160), .o(FE_RN_867_0) );
in01f80 g744808 ( .a(n_36479), .o(n_36480) );
no02f80 g750589 ( .a(n_29405), .b(n_29387), .o(n_29470) );
no03m80 FE_RC_28_0 ( .a(n_6244), .b(n_6321), .c(n_6231), .o(n_6358) );
in01f80 g761213 ( .a(n_19104), .o(n_19135) );
no02f80 g759227 ( .a(n_21220), .b(n_21219), .o(n_21269) );
na02f80 g742435 ( .a(n_37702), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37756) );
na02f80 g764570 ( .a(n_15911), .b(n_14419), .o(n_15953) );
in01f80 g754602 ( .a(n_26886), .o(n_26887) );
in01f80 g771675 ( .a(n_9269), .o(n_9379) );
no02f80 g743419 ( .a(n_36627), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36672) );
no02f80 g778039 ( .a(n_2991), .b(n_2990), .o(n_2992) );
no02f80 g767977 ( .a(n_13034), .b(n_12782), .o(n_13443) );
no02f80 g763913 ( .a(n_17255), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_10_), .o(n_17354) );
in01f80 newInst_2391 ( .a(newNet_2390), .o(newNet_2391) );
no02f80 g779760 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(n_1569) );
in01f80 newInst_1849 ( .a(newNet_1848), .o(newNet_1849) );
in01f80 FE_OCPC993_n_15552 ( .a(n_15552), .o(FE_OCPN993_n_15552) );
no02f80 g737276 ( .a(n_42869), .b(n_42616), .o(n_42890) );
in01f80 g777248 ( .a(n_3616), .o(n_3625) );
na02f80 g745761 ( .a(n_34197), .b(n_34158), .o(n_34248) );
in01f80 g775618 ( .a(n_5472), .o(n_5473) );
in01f80 FE_OCP_RBC3509_n_13860 ( .a(FE_OCP_RBN3508_n_13860), .o(FE_OCP_RBN3509_n_13860) );
na02f80 g768804 ( .a(n_11853), .b(n_11776), .o(n_11989) );
no02f80 g762017 ( .a(n_18590), .b(n_18541), .o(n_18633) );
no02f80 g752235 ( .a(FE_OCPN877_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .o(n_27916) );
na02f80 g761453 ( .a(n_20086), .b(n_19825), .o(n_20133) );
in01f80 g747391 ( .a(n_32678), .o(n_32679) );
no02f80 g761557 ( .a(n_18858), .b(n_18866), .o(n_18942) );
in01f80 g740744 ( .a(n_39969), .o(n_39519) );
no03m80 g768826 ( .a(n_11927), .b(n_11918), .c(n_11919), .o(n_12026) );
in01f80 g775467 ( .a(n_5820), .o(n_5821) );
ao12f80 g748720 ( .a(n_32507), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n_33127) );
ao12f80 g768324 ( .a(n_12489), .b(n_12490), .c(n_12488), .o(n_12538) );
ao12f80 g768895 ( .a(n_11846), .b(n_11845), .c(delay_add_ln22_unr8_stage4_stallmux_q_0_), .o(n_11944) );
ao22s80 FE_RC_3363_0 ( .a(n_31800), .b(n_45518), .c(n_31801), .d(n_45516), .o(n_32266) );
in01f80 g769768 ( .a(n_11263), .o(n_11264) );
in01f80 g749149 ( .a(n_30890), .o(n_30857) );
in01f80 newInst_2166 ( .a(newNet_2165), .o(newNet_2166) );
in01f80 FE_OCP_RBC2695_n_14814 ( .a(n_14814), .o(FE_OCP_RBN2695_n_14814) );
no02f80 g739032 ( .a(n_41135), .b(n_41134), .o(n_41136) );
in01f80 g777751 ( .a(n_4228), .o(n_3385) );
na02f80 g781066 ( .a(sin_out_7), .b(FE_OFN3_n_43918), .o(n_323) );
na02f80 g773110 ( .a(n_7741), .b(n_7710), .o(n_7757) );
na02f80 g760392 ( .a(n_20739), .b(n_20041), .o(n_20835) );
in01f80 g780552 ( .a(n_754), .o(n_749) );
na02f80 g780049 ( .a(n_1239), .b(n_888), .o(n_1245) );
no02f80 g773827 ( .a(n_7065), .b(n_7064), .o(n_7066) );
na02f80 g763112 ( .a(n_17505), .b(n_17580), .o(n_17634) );
no02f80 g756302 ( .a(n_24542), .b(n_24036), .o(n_24665) );
ao22s80 FE_RC_1593_0 ( .a(n_29732), .b(n_45489), .c(FE_OCP_RBN2341_n_29470), .d(n_29719), .o(n_29813) );
na02f80 g773634 ( .a(n_7354), .b(n_7353), .o(n_7403) );
no02f80 g777654 ( .a(n_3428), .b(n_2913), .o(n_3429) );
in01f80 g739112 ( .a(n_41083), .o(n_41072) );
na02f80 FE_RC_2482_0 ( .a(FE_RN_1001_0), .b(n_40495), .o(n_40511) );
in01f80 g760526 ( .a(n_21244), .o(n_20485) );
no02f80 g743111 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n_37088) );
in01f80 FE_OCP_RBC3801_delay_xor_ln22_unr12_stage5_stallmux_q_1_ ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_1_), .o(FE_OCP_RBN3801_delay_xor_ln22_unr12_stage5_stallmux_q_1_) );
no02f80 g746901 ( .a(FE_OCP_RBN3384_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_23_), .o(n_33233) );
na02f80 g773700 ( .a(n_7284), .b(n_7283), .o(n_7285) );
in01f80 g758249 ( .a(n_22918), .o(n_22876) );
na02f80 g778553 ( .a(n_2299), .b(n_2233), .o(n_2340) );
na02f80 g760184 ( .a(n_20657), .b(n_20604), .o(n_20703) );
na02f80 g771743 ( .a(n_8787), .b(FE_OCP_RBN3540_n_8784), .o(n_8850) );
in01f80 newInst_899 ( .a(newNet_271), .o(newNet_899) );
in01f80 g774842 ( .a(n_6435), .o(n_6407) );
na02f80 g760612 ( .a(n_19783), .b(FE_OCPN1790_n_18119), .o(n_19862) );
na02f80 g766336 ( .a(n_14184), .b(n_14185), .o(n_14329) );
in01f80 newInst_3109 ( .a(newNet_3108), .o(newNet_3109) );
no02f80 g759150 ( .a(n_21082), .b(n_21049), .o(n_21230) );
in01f80 g764741 ( .a(n_16415), .o(n_16480) );
na02f80 g778533 ( .a(n_2618), .b(n_2701), .o(n_2729) );
no03m80 FE_RC_2237_0 ( .a(FE_RN_816_0), .b(n_23006), .c(n_23181), .o(FE_RN_817_0) );
in01f80 FE_OCPC1511_n_22280 ( .a(n_22280), .o(FE_OCPN1511_n_22280) );
na02f80 g765955 ( .a(n_14752), .b(n_14751), .o(n_14829) );
na02f80 g736834 ( .a(n_43034), .b(n_43051), .o(n_43064) );
oa12f80 g773395 ( .a(n_7535), .b(n_7558), .c(delay_add_ln22_unr5_stage3_stallmux_q_31_), .o(n_7588) );
no02f80 FE_RC_4173_0 ( .a(FE_RN_1819_0), .b(n_33407), .o(FE_RN_1820_0) );
no02f80 g762142 ( .a(n_18882), .b(n_18812), .o(n_19577) );
in01f80 newInst_2487 ( .a(newNet_2486), .o(newNet_2487) );
no02f80 g754928 ( .a(n_25481), .b(n_24774), .o(n_25648) );
in01f80 g770126 ( .a(n_10850), .o(n_10851) );
no02f80 g761499 ( .a(n_18971), .b(n_18996), .o(n_19024) );
na02f80 g739415 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_7_), .o(n_40726) );
no02f80 g760368 ( .a(n_20104), .b(n_20103), .o(n_20105) );
no02f80 g768382 ( .a(n_12504), .b(n_12239), .o(n_12505) );
na02f80 g766092 ( .a(n_14609), .b(n_14583), .o(n_14716) );
ao12f80 g754529 ( .a(n_25465), .b(n_25464), .c(n_25463), .o(n_27099) );
in01f80 g780290 ( .a(n_970), .o(n_904) );
in01f80 g740330 ( .a(n_40394), .o(n_40395) );
no02f80 g753682 ( .a(n_26537), .b(n_26318), .o(n_26538) );
ao12f80 g751269 ( .a(n_29725), .b(n_29724), .c(n_29723), .o(n_29767) );
na02f80 g737198 ( .a(n_42948), .b(n_42815), .o(n_42964) );
in01f80 newInst_414 ( .a(newNet_413), .o(newNet_414) );
no02f80 g749076 ( .a(n_30957), .b(n_30926), .o(n_31019) );
in01f80 newInst_2311 ( .a(newNet_2310), .o(newNet_2311) );
na02f80 g752551 ( .a(n_27595), .b(n_27396), .o(n_27609) );
in01f80 newInst_2563 ( .a(newNet_2562), .o(newNet_2563) );
na02f80 g764799 ( .a(n_15730), .b(n_15621), .o(n_15731) );
in01f80 g771341 ( .a(n_9057), .o(n_9058) );
no02f80 g745151 ( .a(n_34784), .b(n_34783), .o(n_34785) );
in01f80 g759762 ( .a(n_21564), .o(n_21565) );
na02f80 g773431 ( .a(n_46992), .b(n_6509), .o(n_7581) );
no02f80 g751172 ( .a(n_29909), .b(n_30086), .o(n_30157) );
ao12f80 g777200 ( .a(n_2734), .b(n_3492), .c(n_2656), .o(n_3593) );
in01f80 g774486 ( .a(n_6878), .o(n_6879) );
ao12f80 g737632 ( .a(n_42333), .b(n_42392), .c(n_42374), .o(n_42698) );
in01f80 newInst_905 ( .a(newNet_904), .o(newNet_905) );
in01f80 FE_RC_1107_0 ( .a(FE_RN_332_0), .o(n_2823) );
in01f80 FE_OCP_RBC3376_n_6822 ( .a(n_6822), .o(FE_OCP_RBN3376_n_6822) );
no02f80 g775138 ( .a(n_5989), .b(n_5988), .o(n_6080) );
oa12f80 g759969 ( .a(n_21103), .b(n_21102), .c(n_21101), .o(n_21694) );
in01f80 g765207 ( .a(n_15378), .o(n_15379) );
na02f80 g749767 ( .a(n_31287), .b(n_31187), .o(n_31319) );
na02f80 g784407 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n_46219) );
na02f80 FE_RC_641_0 ( .a(FE_RN_201_0), .b(FE_RN_202_0), .o(FE_RN_203_0) );
no03m80 g739069 ( .a(n_41120), .b(n_41109), .c(n_40816), .o(n_41178) );
no02f80 g737626 ( .a(n_42440), .b(n_42385), .o(n_42461) );
in01f80 g749464 ( .a(n_30599), .o(n_30600) );
in01f80 g759935 ( .a(n_21446), .o(n_21447) );
in01f80 newInst_2698 ( .a(newNet_2697), .o(newNet_2698) );
na02f80 g772520 ( .a(n_8395), .b(n_8399), .o(n_8457) );
in01f80 g764423 ( .a(n_16168), .o(n_16226) );
ao12f80 g781223 ( .a(n_11), .b(n_62), .c(beta_31), .o(n_99) );
oa22f80 FE_RC_771_0 ( .a(n_10032), .b(n_10203), .c(n_10033), .d(n_10200), .o(n_10399) );
in01f80 g739868 ( .a(n_40347), .o(n_40348) );
in01f80 FE_OCPC1249_n_44267 ( .a(FE_OCPN1248_n_44267), .o(FE_OCPN1249_n_44267) );
in01f80 g739937 ( .a(FE_OCP_RBN3046_n_40231), .o(n_40258) );
na02f80 g746382 ( .a(n_33489), .b(n_33488), .o(n_33490) );
in01f80 FE_RC_3074_0 ( .a(n_27126), .o(FE_RN_1353_0) );
no02f80 g754170 ( .a(n_25922), .b(n_25945), .o(n_26021) );
no02f80 g761300 ( .a(n_18925), .b(n_18901), .o(n_19008) );
in01f80 g771888 ( .a(n_8703), .o(n_8704) );
ao22s80 FE_RC_3708_0 ( .a(n_43534), .b(n_43881), .c(n_43533), .d(n_43880), .o(n_43907) );
no02f80 g757555 ( .a(n_22797), .b(n_44061), .o(n_22864) );
na02f80 g744052 ( .a(FE_OCPN3751_n_44222), .b(n_35665), .o(n_36264) );
in01f80 FE_OCP_RBC3705_n_11146 ( .a(n_11146), .o(FE_OCP_RBN3705_n_11146) );
oa22f80 g784544 ( .a(n_11605), .b(FE_OFN801_n_46285), .c(n_11495), .d(FE_OCP_RBN3044_n_46337), .o(n_46365) );
in01f80 g774963 ( .a(n_6198), .o(n_6218) );
in01f80 g742854 ( .a(n_37274), .o(n_37275) );
no02f80 g777385 ( .a(n_3477), .b(n_3364), .o(n_3514) );
oa12f80 g746231 ( .a(n_35073), .b(n_35072), .c(n_35071), .o(n_35629) );
in01f80 FE_RC_79_0 ( .a(n_17742), .o(FE_RN_22_0) );
na02f80 g746526 ( .a(n_34551), .b(FE_OCP_RBN2600_n_34388), .o(n_34616) );
in01f80 g759928 ( .a(n_21448), .o(n_21517) );
in01f80 fopt783094 ( .a(n_8875), .o(n_44570) );
in01f80 g779112 ( .a(n_2237), .o(n_2717) );
no02f80 g739431 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_20_), .o(n_40813) );
na02f80 g744546 ( .a(n_36662), .b(n_36681), .o(n_36685) );
no02f80 g744686 ( .a(n_35184), .b(n_35146), .o(n_35185) );
in01f80 FE_OCP_RBC3069_n_43230 ( .a(FE_OCP_RBN3067_n_43230), .o(FE_OCP_RBN3069_n_43230) );
oa22f80 g747137 ( .a(n_32755), .b(n_32734), .c(n_32756), .d(n_32774), .o(n_34009) );
in01f80 newInst_1005 ( .a(newNet_1004), .o(newNet_1005) );
in01f80 FE_RC_3568_0 ( .a(n_24305), .o(FE_RN_1550_0) );
oa22f80 FE_RC_3823_0 ( .a(n_23414), .b(n_26171), .c(n_23467), .d(FE_OCP_RBN3681_n_26171), .o(n_26320) );
ao12f80 g773386 ( .a(n_7566), .b(n_7565), .c(n_7564), .o(n_8030) );
in01f80 g781394 ( .a(rst), .o(n_264) );
in01f80 g745561 ( .a(n_34622), .o(n_34623) );
in01f80 g745777 ( .a(n_34447), .o(n_34448) );
na02f80 g742388 ( .a(n_37771), .b(n_37770), .o(n_37778) );
no02f80 g758714 ( .a(n_21658), .b(n_21507), .o(n_21688) );
na02f80 FE_RC_668_0 ( .a(FE_RN_210_0), .b(FE_RN_211_0), .o(FE_RN_212_0) );
na02f80 g780042 ( .a(n_1240), .b(n_963), .o(n_1248) );
in01f80 newInst_113 ( .a(newNet_65), .o(newNet_113) );
no02f80 g783786 ( .a(n_47008), .b(n_4182), .o(n_45462) );
na04m80 g747294 ( .a(n_32433), .b(n_32577), .c(n_32582), .d(n_32578), .o(n_32583) );
na02f80 g759897 ( .a(n_21374), .b(n_21514), .o(n_21670) );
na02f80 g752803 ( .a(n_28053), .b(n_28075), .o(n_28637) );
no02f80 FE_RC_3477_0 ( .a(FE_RN_1494_0), .b(n_36352), .o(n_36381) );
na02f80 g766130 ( .a(n_14450), .b(n_14476), .o(n_14557) );
no02f80 g767070 ( .a(n_13613), .b(n_13612), .o(n_13614) );
no02f80 g743246 ( .a(n_36783), .b(n_36742), .o(n_36801) );
na02f80 g737689 ( .a(n_42367), .b(n_41991), .o(n_42395) );
na02f80 g762739 ( .a(FE_OCPN854_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_19_), .o(n_17922) );
no02f80 FE_RC_1926_0 ( .a(n_35290), .b(FE_RN_608_0), .o(FE_RN_609_0) );
na02f80 g749123 ( .a(n_30914), .b(n_27518), .o(n_30915) );
no02f80 g739062 ( .a(n_41128), .b(n_41127), .o(n_41129) );
in01f80 g748034 ( .a(n_33000), .o(n_33001) );
in01f80 newInst_772 ( .a(newNet_771), .o(newNet_772) );
in01f80 g754143 ( .a(n_26027), .o(n_26059) );
na02f80 g755124 ( .a(n_25201), .b(n_24422), .o(n_25413) );
in01f80 g736815 ( .a(n_43621), .o(n_43622) );
no02f80 g768033 ( .a(n_12790), .b(n_12838), .o(n_12911) );
na02f80 g736386 ( .a(n_43759), .b(n_43433), .o(n_43789) );
in01f80 FE_OCPC1738_n_19052 ( .a(FE_OCPN1737_n_19052), .o(FE_OCPN1738_n_19052) );
in01f80 newInst_151 ( .a(newNet_150), .o(newNet_151) );
no02f80 g764184 ( .a(n_16497), .b(n_16496), .o(n_16588) );
in01f80 g770891 ( .a(n_9965), .o(n_9966) );
no02f80 g761762 ( .a(n_18564), .b(n_17661), .o(n_18566) );
in01f80 newInst_163 ( .a(newNet_162), .o(newNet_163) );
in01f80 newInst_3114 ( .a(newNet_3113), .o(newNet_3114) );
in01f80 newInst_2383 ( .a(newNet_2382), .o(newNet_2383) );
ao12f80 g746997 ( .a(n_34044), .b(n_34043), .c(n_34042), .o(n_34733) );
na02f80 g764788 ( .a(n_16359), .b(n_16358), .o(n_16360) );
oa12f80 g765255 ( .a(n_15574), .b(n_15573), .c(n_15572), .o(n_16100) );
in01f80 g753132 ( .a(n_27498), .o(n_27499) );
na02f80 g744666 ( .a(n_35215), .b(n_35239), .o(n_35316) );
no02f80 g775730 ( .a(n_5877), .b(n_5626), .o(n_5659) );
no02f80 g736732 ( .a(n_43325), .b(n_43270), .o(n_43326) );
na02f80 g761869 ( .a(n_18742), .b(n_18741), .o(n_18784) );
no02f80 g740004 ( .a(n_40038), .b(n_40152), .o(n_40153) );
na02f80 g770314 ( .a(n_10612), .b(FE_OCP_RBN3637_n_44490), .o(n_10724) );
in01f80 newInst_1510 ( .a(newNet_1283), .o(newNet_1510) );
oa22f80 g738157 ( .a(n_41981), .b(n_41851), .c(n_41980), .d(n_41852), .o(n_42046) );
na02f80 g768581 ( .a(n_12191), .b(n_12270), .o(n_12440) );
no02f80 g778092 ( .a(n_2942), .b(n_2217), .o(n_2943) );
na02f80 g774722 ( .a(n_6375), .b(n_6417), .o(n_6500) );
no02f80 g775646 ( .a(n_5173), .b(n_5190), .o(n_5308) );
na02f80 g758087 ( .a(n_44275), .b(FE_OCP_RBN1370_n_20763), .o(n_22311) );
in01f80 g757862 ( .a(n_22318), .o(n_22319) );
in01f80 newInst_350 ( .a(newNet_349), .o(newNet_350) );
in01f80 FE_OFC817_n_2285 ( .a(FE_OFN834_n_2285), .o(FE_OFN817_n_2285) );
no02f80 g747128 ( .a(n_32953), .b(n_32952), .o(n_32968) );
oa22f80 g749343 ( .a(n_31977), .b(n_31568), .c(n_31978), .d(n_31567), .o(n_32065) );
na02f80 g761913 ( .a(n_18302), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_), .o(n_18372) );
in01f80 g744477 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_), .o(n_36773) );
in01f80 g756548 ( .a(n_23993), .o(n_23994) );
no02f80 g737531 ( .a(n_42337), .b(n_42335), .o(n_42336) );
no02f80 g748373 ( .a(FE_OCPN1052_n_31674), .b(n_31795), .o(n_31823) );
na02f80 g780932 ( .a(n_457), .b(n_485), .o(n_489) );
no02f80 g751160 ( .a(n_30303), .b(n_30082), .o(n_30380) );
na02f80 g751530 ( .a(n_28453), .b(n_28452), .o(n_28506) );
in01f80 FE_OCP_RBC3444_n_37945 ( .a(n_37945), .o(FE_OCP_RBN3444_n_37945) );
oa12f80 g750166 ( .a(n_29764), .b(n_29755), .c(n_29728), .o(n_29795) );
no02f80 g763171 ( .a(n_16975), .b(n_17248), .o(n_17343) );
no02f80 g779775 ( .a(n_1780), .b(n_1381), .o(n_1444) );
in01f80 newInst_3153 ( .a(newNet_3152), .o(newNet_3153) );
no02f80 g740820 ( .a(n_39351), .b(n_39383), .o(n_39853) );
in01f80 newInst_244 ( .a(newNet_243), .o(newNet_244) );
no02f80 g775544 ( .a(n_5891), .b(n_5765), .o(n_5889) );
ao12f80 g756831 ( .a(n_24106), .b(n_24075), .c(n_24105), .o(n_24153) );
oa12f80 g771026 ( .a(n_9962), .b(n_10001), .c(n_9961), .o(n_10044) );
ao22s80 FE_RC_1542_0 ( .a(n_15450), .b(n_15989), .c(n_15449), .d(n_15990), .o(n_16146) );
no02f80 g753873 ( .a(n_26283), .b(n_26254), .o(n_26364) );
no02f80 FE_RC_4070_0 ( .a(n_35911), .b(n_35910), .o(FE_RN_1772_0) );
na02f80 g764824 ( .a(n_15652), .b(n_14618), .o(n_15730) );
no02f80 FE_RC_3405_0 ( .a(FE_RN_616_0), .b(FE_RN_1474_0), .o(n_19414) );
na02f80 g740812 ( .a(n_39438), .b(n_39405), .o(n_39535) );
na02f80 g768906 ( .a(n_44356), .b(n_11662), .o(n_11883) );
no02f80 g750557 ( .a(n_29354), .b(n_29326), .o(n_29425) );
in01f80 g757481 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .o(n_22803) );
no02f80 FE_RC_2838_0 ( .a(n_17881), .b(n_19148), .o(FE_RN_1220_0) );
no02f80 g761437 ( .a(n_18893), .b(n_17783), .o(n_18922) );
no02f80 g761751 ( .a(n_18565), .b(n_18599), .o(n_18795) );
in01f80 FE_RC_2930_0 ( .a(n_39371), .o(FE_RN_1277_0) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_17_ ( .ck(newNet_3327), .d(n_32085), .o(delay_add_ln22_unr20_stage8_stallmux_q_17_) );
na02f80 g776302 ( .a(n_4396), .b(n_4093), .o(n_4439) );
no02f80 g750621 ( .a(n_29339), .b(n_29304), .o(n_29401) );
no02f80 g738085 ( .a(n_42107), .b(n_42542), .o(n_42108) );
in01f80 g756800 ( .a(n_23473), .o(n_23474) );
ao12f80 g750220 ( .a(FE_OCP_RBN2446_n_29684), .b(n_29788), .c(n_29671), .o(n_29809) );
in01f80 newInst_2400 ( .a(newNet_1602), .o(newNet_2400) );
ao12f80 g756358 ( .a(n_23637), .b(n_23859), .c(n_23626), .o(n_23929) );
in01f80 g768003 ( .a(n_12819), .o(n_12820) );
in01f80 g767005 ( .a(n_14213), .o(n_14075) );
no02f80 g740417 ( .a(FE_OCP_RBN3022_n_39942), .b(n_39555), .o(n_40240) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_16_ ( .ck(newNet_183), .d(n_46351), .o(delay_xor_ln22_unr9_stage4_stallmux_q_16_) );
in01f80 g745571 ( .a(n_34351), .o(n_34322) );
no02f80 g760566 ( .a(n_19857), .b(n_19695), .o(n_19890) );
in01f80 g763436 ( .a(n_17069), .o(n_17070) );
in01f80 FE_OCP_RBC3673_n_30820 ( .a(n_30820), .o(FE_OCP_RBN3673_n_30820) );
na02f80 g779173 ( .a(n_1969), .b(n_1968), .o(n_2156) );
na02f80 g775545 ( .a(n_5553), .b(n_4862), .o(n_5716) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_14_ ( .ck(newNet_1761), .d(n_22144), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_) );
oa12f80 g745893 ( .a(n_35322), .b(n_35321), .c(n_35320), .o(n_35391) );
in01f80 g764064 ( .a(n_17093), .o(n_17498) );
in01f80 g738067 ( .a(n_42137), .o(n_42113) );
oa12f80 g774900 ( .a(n_6197), .b(n_6149), .c(n_6153), .o(n_6230) );
in01f80 g776845 ( .a(n_4126), .o(n_4127) );
in01f80 g766821 ( .a(n_14429), .o(n_14528) );
in01f80 g766857 ( .a(n_14044), .o(n_14081) );
na02f80 g772229 ( .a(n_8621), .b(n_7609), .o(n_8622) );
in01f80 FE_OCP_RBC2341_n_29470 ( .a(n_29470), .o(FE_OCP_RBN2341_n_29470) );
in01f80 FE_RC_819_0 ( .a(n_8986), .o(FE_RN_247_0) );
ao12f80 g767237 ( .a(n_13210), .b(n_13697), .c(n_13248), .o(n_13737) );
no02f80 g777728 ( .a(n_3326), .b(n_3314), .o(n_3315) );
no02f80 g775439 ( .a(n_5770), .b(n_47197), .o(n_5796) );
no02f80 g768660 ( .a(n_12154), .b(n_12153), .o(n_12155) );
in01f80 newInst_3300 ( .a(newNet_1600), .o(newNet_3300) );
no02f80 g765556 ( .a(FE_OCP_RBN2716_n_14982), .b(n_14514), .o(n_15180) );
na02f80 g765087 ( .a(n_16024), .b(n_15837), .o(n_16025) );
in01f80 FE_RC_3491_0 ( .a(n_37070), .o(FE_RN_1505_0) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_9_ ( .ck(newNet_3356), .d(n_27046), .o(delay_add_ln22_unr17_stage7_stallmux_q_9_) );
in01f80 newInst_1392 ( .a(newNet_1391), .o(newNet_1392) );
in01f80 FE_OCP_RBC3706_n_11146 ( .a(n_11146), .o(FE_OCP_RBN3706_n_11146) );
na02f80 g758048 ( .a(n_22732), .b(n_22456), .o(n_22733) );
no02f80 g778487 ( .a(n_2361), .b(n_2794), .o(n_2415) );
in01f80 g762329 ( .a(n_18096), .o(n_18115) );
na02f80 g757262 ( .a(n_23070), .b(n_21457), .o(n_23196) );
oa22f80 g739402 ( .a(FE_OCPN897_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_), .c(n_44775), .d(n_40480), .o(n_41043) );
in01f80 FE_OCPC990_n_22249 ( .a(n_22249), .o(FE_OCPN990_n_22249) );
in01f80 FE_OCP_DRV_C1541_n_26125 ( .a(n_26125), .o(FE_OCP_DRV_N1541_n_26125) );
no02f80 FE_RC_2542_0 ( .a(FE_RN_1038_0), .b(n_39143), .o(FE_RN_1039_0) );
no02f80 g762025 ( .a(n_18356), .b(n_18337), .o(n_18391) );
in01f80 g765405 ( .a(n_15151), .o(n_15189) );
in01f80 FE_OCP_RBC1375_n_20889 ( .a(n_20889), .o(FE_OCP_RBN1375_n_20889) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_13_ ( .ck(newNet_3254), .d(n_36422), .o(delay_add_ln22_unr23_stage9_stallmux_q_13_) );
na02f80 g748080 ( .a(n_31745), .b(n_31776), .o(n_31854) );
na02f80 FE_RC_3411_0 ( .a(FE_RN_1477_0), .b(FE_RN_739_0), .o(n_21236) );
na02f80 g759097 ( .a(n_21093), .b(FE_OCP_RBN3663_n_20750), .o(n_21130) );
no02f80 g760113 ( .a(FE_OCP_RBN2662_n_20333), .b(n_20332), .o(n_20463) );
ao22s80 FE_RC_1367_0 ( .a(n_39202), .b(n_39517), .c(n_39201), .d(n_39516), .o(n_39586) );
na02f80 g737890 ( .a(n_42270), .b(n_42569), .o(n_42656) );
in01f80 newInst_1111 ( .a(newNet_1110), .o(newNet_1111) );
in01f80 newInst_945 ( .a(newNet_867), .o(newNet_945) );
ao12f80 g750292 ( .a(n_30722), .b(n_30721), .c(n_30720), .o(n_31216) );
in01f80 FE_OCP_RBC3307_n_44722 ( .a(n_44722), .o(FE_OCP_RBN3307_n_44722) );
in01f80 FE_OCPC1509_n_44174 ( .a(n_44174), .o(FE_OCPN1509_n_44174) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_21_ ( .ck(newNet_2945), .d(n_6313), .o(delay_add_ln22_unr5_stage3_stallmux_q_21_) );
na02f80 g771381 ( .a(n_9401), .b(FE_OCP_RBN2605_FE_OCPN899_n_44593), .o(n_9586) );
na02f80 g759363 ( .a(n_21069), .b(n_20675), .o(n_21070) );
no02f80 g763847 ( .a(n_16682), .b(FE_OCP_RBN3062_FE_RN_640_0), .o(n_16728) );
na02f80 g777766 ( .a(n_3370), .b(n_4211), .o(n_3392) );
na03f80 FE_RC_2318_0 ( .a(FE_RN_881_0), .b(n_35959), .c(n_35927), .o(FE_RN_882_0) );
no02f80 g740752 ( .a(n_39311), .b(n_39366), .o(n_39413) );
ao12f80 g760840 ( .a(n_19565), .b(n_19287), .c(n_18032), .o(n_19441) );
in01f80 g769963 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_13_), .o(n_11101) );
in01f80 newInst_1413 ( .a(newNet_108), .o(newNet_1413) );
in01f80 g780623 ( .a(n_684), .o(n_685) );
in01f80 FE_OCP_RBC3464_n_7886 ( .a(n_7886), .o(FE_OCP_RBN3464_n_7886) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_6_ ( .ck(newNet_3368), .d(n_26810), .o(delay_add_ln22_unr17_stage7_stallmux_q_6_) );
na02f80 g766884 ( .a(n_14304), .b(n_14210), .o(n_14341) );
no02f80 g743906 ( .a(n_36942), .b(n_46237), .o(n_36927) );
na02f80 g773400 ( .a(n_7584), .b(n_7595), .o(n_7633) );
in01f80 g751995 ( .a(n_29004), .o(n_29488) );
in01f80 newInst_3501 ( .a(newNet_3500), .o(newNet_3501) );
in01f80 g780443 ( .a(n_796), .o(n_787) );
no02f80 g750668 ( .a(n_29325), .b(n_29302), .o(n_29421) );
in01f80 g768458 ( .a(n_12361), .o(n_12401) );
oa12f80 g757303 ( .a(n_23129), .b(n_23106), .c(n_44071), .o(n_23335) );
oa12f80 g761754 ( .a(n_19230), .b(n_19229), .c(n_19228), .o(n_19337) );
in01f80 g764397 ( .a(n_16330), .o(n_16278) );
in01f80 FE_RC_142_0 ( .a(FE_RN_41_0), .o(n_18268) );
no02f80 g736938 ( .a(n_43038), .b(n_46941), .o(n_43271) );
no02f80 g760640 ( .a(FE_OCP_RBN1182_n_19726), .b(FE_OCP_RBN3829_n_19204), .o(n_19780) );
no02f80 FE_RC_2491_0 ( .a(FE_RN_1008_0), .b(n_24068), .o(n_24081) );
na02f80 g757632 ( .a(n_22601), .b(n_22230), .o(n_22602) );
in01f80 FE_OCP_RBC2501_n_13896 ( .a(FE_OCP_RBN3528_n_13765), .o(FE_OCP_RBN2501_n_13896) );
in01f80 g738094 ( .a(n_42087), .o(n_42088) );
in01f80 newInst_844 ( .a(newNet_843), .o(newNet_844) );
no02f80 g744493 ( .a(n_35441), .b(n_35465), .o(n_35493) );
no02f80 FE_RC_91_0 ( .a(FE_RN_27_0), .b(FE_OCP_RBN3208_n_44365), .o(FE_RN_29_0) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_1_ ( .ck(newNet_919), .d(n_27725), .o(n_44422) );
in01f80 g748062 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_10_), .o(n_32861) );
no02f80 g760626 ( .a(n_19808), .b(FE_OFN815_n_19807), .o(n_19887) );
na02f80 g738582 ( .a(n_41536), .b(n_41663), .o(n_41925) );
oa22f80 FE_RC_4136_0 ( .a(n_22801), .b(n_22857), .c(n_22793), .d(n_22790), .o(n_22892) );
na02f80 g738369 ( .a(n_41702), .b(FE_OCP_RBN2316_n_41420), .o(n_41771) );
no02f80 g747869 ( .a(n_33131), .b(n_33130), .o(n_33132) );
in01f80 g751956 ( .a(n_29242), .o(n_29243) );
in01f80 g754694 ( .a(n_26812), .o(n_26813) );
no02f80 g770682 ( .a(n_10188), .b(n_10116), .o(n_10262) );
in01f80 newInst_345 ( .a(newNet_344), .o(newNet_345) );
na02f80 g750143 ( .a(n_29955), .b(n_29889), .o(n_30025) );
ao12f80 g769669 ( .a(n_11104), .b(n_11316), .c(n_47199), .o(n_11362) );
na02f80 g776490 ( .a(n_4425), .b(n_4393), .o(n_4490) );
na02f80 g739668 ( .a(n_44692), .b(n_40222), .o(n_40555) );
in01f80 g765806 ( .a(n_14889), .o(n_14890) );
in01f80 g778322 ( .a(n_3857), .o(n_2962) );
in01f80 FE_RC_908_0 ( .a(n_11478), .o(FE_RN_267_0) );
in01f80 g737268 ( .a(n_42906), .o(n_43170) );
no02f80 g760776 ( .a(n_19535), .b(n_19512), .o(n_19564) );
no02f80 g770142 ( .a(FE_OCP_RBN2899_n_44853), .b(n_10412), .o(n_10702) );
ao12f80 g740882 ( .a(n_38967), .b(n_39167), .c(n_38924), .o(n_39218) );
oa22f80 g748208 ( .a(FE_OCPN981_n_31961), .b(n_32076), .c(FE_OCPN880_n_31944), .d(n_30326), .o(n_32178) );
no02f80 g741508 ( .a(n_38723), .b(n_38719), .o(n_38743) );
in01f80 g743266 ( .a(n_36783), .o(n_36790) );
in01f80 g758154 ( .a(n_23148), .o(n_23149) );
na02f80 g767032 ( .a(FE_OCP_RBN3533_n_13765), .b(n_13975), .o(n_14041) );
na02f80 g740828 ( .a(n_39375), .b(n_39320), .o(n_39438) );
no02f80 g743972 ( .a(n_47264), .b(n_35905), .o(n_35951) );
in01f80 g761119 ( .a(n_19264), .o(n_19301) );
na02f80 g765099 ( .a(n_16347), .b(n_16346), .o(n_16348) );
in01f80 g743489 ( .a(n_36646), .o(n_36647) );
in01f80 g752026 ( .a(n_28102), .o(n_28149) );
na02f80 g767989 ( .a(n_13112), .b(n_13103), .o(n_13584) );
in01f80 newInst_913 ( .a(newNet_912), .o(newNet_913) );
ao12f80 g784390 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46200) );
na02f80 g763375 ( .a(FE_OCP_RBN3725_n_16975), .b(FE_OCP_RBN2812_n_15433), .o(n_17332) );
no02f80 g769358 ( .a(n_11784), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11838) );
na02f80 FE_RC_3923_0 ( .a(n_44061), .b(FE_RN_1696_0), .o(n_22820) );
in01f80 FE_OCP_RBC3674_FE_RN_1581_0 ( .a(FE_RN_1581_0), .o(FE_OCP_RBN3674_FE_RN_1581_0) );
in01f80 g744128 ( .a(n_36260), .o(n_36261) );
in01f80 g777550 ( .a(n_4182), .o(n_4556) );
na02f80 g741480 ( .a(n_38753), .b(n_38752), .o(n_38783) );
in01f80 g778737 ( .a(n_2609), .o(n_2643) );
in01f80 newInst_3717 ( .a(newNet_591), .o(newNet_3717) );
oa22f80 g779881 ( .a(FE_OCPN875_n_44672), .b(n_1040), .c(n_44637), .d(n_984), .o(n_1348) );
in01f80 g749538 ( .a(n_31782), .o(n_31815) );
in01f80 newInst_2627 ( .a(newNet_2626), .o(newNet_2627) );
oa12f80 g756417 ( .a(n_23856), .b(n_23766), .c(n_23821), .o(n_23857) );
oa12f80 g773115 ( .a(n_7960), .b(n_8232), .c(n_7982), .o(n_8820) );
ao12f80 g736535 ( .a(n_43489), .b(n_43659), .c(n_43553), .o(n_43696) );
no02f80 g752915 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_26_), .o(n_28128) );
in01f80 g770455 ( .a(n_10562), .o(n_10563) );
in01f80 g780401 ( .a(n_876), .o(n_858) );
no02f80 g761136 ( .a(n_19105), .b(n_18708), .o(n_19151) );
in01f80 newInst_1324 ( .a(newNet_1323), .o(newNet_1324) );
in01f80 g778395 ( .a(n_2505), .o(n_2506) );
na02f80 g774714 ( .a(n_6332), .b(n_6215), .o(n_6349) );
na02f80 g774895 ( .a(n_6303), .b(n_6276), .o(n_6419) );
na02f80 g778162 ( .a(n_2747), .b(n_2192), .o(n_2793) );
no02f80 g771433 ( .a(n_8975), .b(n_8189), .o(n_9089) );
no02f80 g747223 ( .a(n_33801), .b(n_33800), .o(n_33802) );
oa22f80 g752360 ( .a(n_27720), .b(n_24059), .c(n_27698), .d(n_27796), .o(n_27741) );
ao12f80 g757412 ( .a(n_22987), .b(n_22933), .c(n_22674), .o(n_23014) );
in01f80 newInst_1260 ( .a(newNet_1259), .o(newNet_1260) );
na02f80 g765663 ( .a(n_14962), .b(FE_OCP_RBN3485_n_13667), .o(n_14986) );
ao12f80 g772833 ( .a(n_7987), .b(n_7966), .c(n_7931), .o(n_8140) );
ao12f80 g741881 ( .a(n_38238), .b(n_38338), .c(n_38283), .o(n_38360) );
na02f80 g767637 ( .a(n_12804), .b(n_12772), .o(n_12907) );
in01f80 FE_RC_1882_0 ( .a(FE_RN_585_0), .o(n_28182) );
oa12f80 g777686 ( .a(n_3102), .b(n_3303), .c(n_3140), .o(n_3334) );
na02f80 g776277 ( .a(n_4521), .b(n_4439), .o(n_4652) );
no02f80 g748897 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .o(n_32603) );
in01f80 g768433 ( .a(n_12495), .o(n_12496) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_17_ ( .ck(newNet_3541), .d(n_22596), .o(delay_add_ln22_unr14_stage6_stallmux_q_17_) );
in01f80 g771844 ( .a(n_10123), .o(n_10208) );
ao22s80 g751332 ( .a(n_28612), .b(n_28416), .c(n_28552), .d(n_28415), .o(n_28656) );
no02f80 g742056 ( .a(FE_OCP_RBN2257_n_37844), .b(FE_OCPN1736_n_37877), .o(n_37979) );
na03f80 FE_RC_4156_0 ( .a(FE_RN_1808_0), .b(n_32919), .c(FE_RN_1708_0), .o(n_33207) );
in01f80 FE_OCP_RBC3040_n_46337 ( .a(n_46337), .o(FE_OCP_RBN3040_n_46337) );
na02f80 g749139 ( .a(n_30860), .b(n_30859), .o(n_30877) );
na02f80 g773772 ( .a(n_7222), .b(n_7221), .o(n_7223) );
in01f80 g754248 ( .a(n_25938), .o(n_25937) );
na02f80 g773002 ( .a(n_7713), .b(n_7683), .o(n_7777) );
in01f80 newInst_2909 ( .a(newNet_1547), .o(newNet_2909) );
na02f80 g767644 ( .a(n_13284), .b(n_13243), .o(n_13285) );
na02f80 g738115 ( .a(n_42046), .b(n_42500), .o(n_42047) );
no02f80 g777286 ( .a(n_4556), .b(n_4760), .o(n_5091) );
na02f80 g775199 ( .a(n_6008), .b(n_5961), .o(n_6032) );
na02f80 g763220 ( .a(n_17141), .b(FE_OCPN1756_n_16923), .o(n_17282) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_8_ ( .ck(newNet_2232), .d(n_40411), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_) );
no02f80 g777779 ( .a(n_3379), .b(n_3378), .o(n_3396) );
na02f80 g744023 ( .a(n_36065), .b(n_36096), .o(n_36097) );
in01f80 FE_OCP_RBC2708_n_15135 ( .a(FE_OCP_RBN3621_n_15135), .o(FE_OCP_RBN2708_n_15135) );
in01f80 g760434 ( .a(n_20030), .o(n_20031) );
no02f80 g762386 ( .a(n_45002), .b(n_18688), .o(n_18724) );
oa12f80 g784392 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_46202) );
no02f80 g763302 ( .a(n_17488), .b(n_16118), .o(n_17087) );
na02f80 g768963 ( .a(n_11779), .b(n_11762), .o(n_11881) );
no02f80 g741476 ( .a(n_38758), .b(n_38716), .o(n_38788) );
in01f80 newInst_3546 ( .a(newNet_3545), .o(newNet_3546) );
na02f80 g751556 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_22_), .o(n_28522) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_2_ ( .ck(newNet_380), .d(n_40588), .o(delay_xor_ln22_unr28_stage10_stallmux_q_2_) );
na02f80 g769721 ( .a(n_11173), .b(n_11106), .o(n_11242) );
no02f80 g771406 ( .a(n_9561), .b(n_9656), .o(n_9737) );
no02f80 g746270 ( .a(FE_OCP_RBN3411_n_33547), .b(FE_OCP_RBN1680_n_33491), .o(n_33592) );
no02f80 g771542 ( .a(n_8817), .b(n_7658), .o(n_8843) );
ao12f80 g746043 ( .a(n_35164), .b(n_35163), .c(n_35162), .o(n_35258) );
no02f80 g765778 ( .a(n_15362), .b(n_15361), .o(n_15363) );
no02f80 g741538 ( .a(n_38671), .b(n_38649), .o(n_38703) );
na02f80 g753391 ( .a(n_26988), .b(n_26963), .o(n_27027) );
no02f80 g763312 ( .a(n_17578), .b(n_17432), .o(n_17736) );
na02f80 g750784 ( .a(n_29121), .b(n_28724), .o(n_29165) );
in01f80 g769389 ( .a(n_11407), .o(n_11420) );
na02f80 g771833 ( .a(n_9323), .b(n_9226), .o(n_9558) );
no02f80 g776636 ( .a(n_4285), .b(n_4121), .o(n_4352) );
na02f80 g781057 ( .a(sin_out_17), .b(FE_OFN3_n_43918), .o(n_324) );
oa22f80 FE_RC_2402_0 ( .a(n_42585), .b(FE_OCP_RBN2970_n_42896), .c(n_42586), .d(n_42896), .o(n_42959) );
no02f80 g759903 ( .a(n_21406), .b(n_21246), .o(n_21774) );
in01f80 g755828 ( .a(n_25142), .o(n_25169) );
in01f80 g777664 ( .a(n_3386), .o(n_3401) );
na02f80 g736740 ( .a(n_43389), .b(n_43400), .o(n_43471) );
na02f80 g778615 ( .a(n_2741), .b(n_2752), .o(n_2814) );
no02f80 g757295 ( .a(n_23044), .b(FE_OCPN1020_n_23078), .o(n_23110) );
in01f80 g754847 ( .a(n_25593), .o(n_25594) );
in01f80 g763944 ( .a(n_16661), .o(n_16662) );
in01f80 g780307 ( .a(n_969), .o(n_1003) );
in01f80 g755502 ( .a(n_24652), .o(n_24687) );
in01f80 g763658 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .o(n_16830) );
na02f80 g779612 ( .a(n_1559), .b(n_1558), .o(n_1735) );
na02f80 g777730 ( .a(FE_OCP_RBN3539_n_3335), .b(n_2759), .o(n_3384) );
no02f80 g737709 ( .a(FE_OCPN885_n_42216), .b(n_42077), .o(n_42419) );
no02f80 g753085 ( .a(n_27146), .b(n_27121), .o(n_27305) );
in01f80 g763280 ( .a(n_17401), .o(n_17442) );
in01f80 newInst_2051 ( .a(newNet_1028), .o(newNet_2051) );
in01f80 g749339 ( .a(n_46958), .o(n_30814) );
in01f80 FE_OCPC947_n_41382 ( .a(n_41382), .o(FE_OCPN947_n_41382) );
no02f80 g763678 ( .a(n_17605), .b(n_17604), .o(n_18293) );
no02f80 g780480 ( .a(n_831), .b(n_795), .o(n_759) );
ao12f80 g751614 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .c(delay_add_ln22_unr17_stage7_stallmux_q_29_), .o(n_28761) );
in01f80 g768501 ( .a(n_12385), .o(n_12386) );
ao12f80 g753606 ( .a(n_26742), .b(n_27284), .c(n_26709), .o(n_27367) );
in01f80 g756320 ( .a(n_24585), .o(n_24586) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_4_ ( .ck(newNet_884), .d(n_32337), .o(delay_xor_ln21_unr21_stage8_stallmux_q_4_) );
no02f80 g746392 ( .a(n_33409), .b(n_32973), .o(n_33433) );
in01f80 g765586 ( .a(n_16136), .o(n_15744) );
no02f80 g769761 ( .a(n_11053), .b(n_11056), .o(n_11125) );
ao12f80 g768697 ( .a(n_11728), .b(n_44450), .c(n_11632), .o(n_12140) );
in01f80 g782661 ( .a(n_44055), .o(n_44056) );
oa12f80 g775105 ( .a(n_5788), .b(n_5996), .c(n_5769), .o(n_6067) );
in01f80 FE_OFC786_n_25834 ( .a(n_25834), .o(FE_OFN786_n_25834) );
oa22f80 FE_RC_3330_0 ( .a(n_29501), .b(n_29730), .c(n_29530), .d(n_29749), .o(n_29773) );
na02f80 FE_RC_4011_0 ( .a(FE_RN_1741_0), .b(n_30467), .o(n_30514) );
no02f80 g743286 ( .a(n_36743), .b(n_36711), .o(n_36759) );
ao12f80 g742527 ( .a(FE_OCP_RBN3393_n_37557), .b(FE_OCP_RBN2174_n_37559), .c(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37644) );
na03f80 g756289 ( .a(n_23838), .b(n_24610), .c(n_23722), .o(n_24770) );
in01f80 g778328 ( .a(n_2920), .o(n_2921) );
in01f80 FE_OCP_RBC2240_n_44881 ( .a(FE_OCP_RBN3427_n_44881), .o(FE_OCP_RBN2240_n_44881) );
in01f80 FE_OCP_DRV_C1599_n_21493 ( .a(n_21493), .o(FE_OCP_DRV_N1599_n_21493) );
no02f80 g736798 ( .a(n_43215), .b(n_43179), .o(n_43180) );
no02f80 g746374 ( .a(n_33411), .b(n_33163), .o(n_33473) );
no02f80 g747722 ( .a(n_33741), .b(n_33792), .o(n_34251) );
in01f80 FE_OCP_RBC3610_FE_OCPN1797_n_20333 ( .a(FE_OCPN1797_n_20333), .o(FE_OCP_RBN3610_FE_OCPN1797_n_20333) );
in01f80 g759370 ( .a(n_20802), .o(n_20803) );
na02f80 g742714 ( .a(n_37480), .b(n_37479), .o(n_37481) );
in01f80 g743925 ( .a(n_35868), .o(n_35914) );
in01f80 g771296 ( .a(n_9413), .o(n_9414) );
no02f80 g770941 ( .a(n_9747), .b(FE_OFN755_n_44461), .o(n_9868) );
no02f80 g757781 ( .a(n_22482), .b(n_22481), .o(n_22483) );
in01f80 g741799 ( .a(n_38493), .o(n_38516) );
ao22s80 g738771 ( .a(n_41339), .b(n_41343), .c(n_41324), .d(n_40658), .o(n_41369) );
no02f80 g746836 ( .a(n_33151), .b(n_33180), .o(n_33606) );
ao12f80 g748589 ( .a(n_31462), .b(n_31442), .c(n_31440), .o(n_31546) );
na02f80 g743984 ( .a(n_36034), .b(n_35976), .o(n_36100) );
in01f80 g736769 ( .a(n_43560), .o(n_43561) );
no02f80 g766683 ( .a(n_13729), .b(n_12869), .o(n_13757) );
no02f80 g767583 ( .a(n_13262), .b(n_13087), .o(n_13322) );
in01f80 g736465 ( .a(n_43742), .o(n_43768) );
in01f80 g763023 ( .a(n_17557), .o(n_17558) );
in01f80 g754486 ( .a(n_25568), .o(n_25597) );
in01f80 newInst_2421 ( .a(newNet_1227), .o(newNet_2421) );
in01f80 newInst_3341 ( .a(newNet_163), .o(newNet_3341) );
in01f80 newInst_1559 ( .a(newNet_1558), .o(newNet_1559) );
oa12f80 g779199 ( .a(n_1860), .b(n_1859), .c(n_1858), .o(n_2292) );
in01f80 newInst_2918 ( .a(newNet_2917), .o(newNet_2918) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_28_ ( .ck(newNet_3607), .d(n_44447), .o(delay_add_ln22_unr11_stage5_stallmux_q_28_) );
in01f80 FE_OFC802_n_46285 ( .a(FE_OFN798_n_46285), .o(FE_OFN802_n_46285) );
in01f80 FE_OCPC1756_n_16923 ( .a(FE_OCPN1755_n_16923), .o(FE_OCPN1756_n_16923) );
no02f80 g756456 ( .a(n_23851), .b(n_23850), .o(n_23852) );
in01f80 newInst_1990 ( .a(newNet_1989), .o(newNet_1990) );
na02f80 g754361 ( .a(n_25758), .b(n_25447), .o(n_25788) );
in01f80 newInst_2649 ( .a(newNet_2648), .o(newNet_2649) );
na02f80 g773610 ( .a(n_7360), .b(n_7308), .o(n_7361) );
no02f80 g780242 ( .a(n_1080), .b(n_1079), .o(n_1081) );
na02f80 g755268 ( .a(n_24944), .b(n_24943), .o(n_25018) );
in01f80 g755653 ( .a(FE_OCP_RBN2421_n_24505), .o(n_25104) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_1_ ( .ck(newNet_2857), .d(n_9760), .o(delay_add_ln22_unr8_stage4_stallmux_q_1_) );
in01f80 FE_RC_3754_0 ( .a(n_40711), .o(FE_RN_1649_0) );
na02f80 g750474 ( .a(n_29574), .b(n_29573), .o(n_29589) );
no02f80 g774303 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_10_), .o(n_6770) );
no02f80 g772499 ( .a(n_8487), .b(n_8488), .o(n_8570) );
na02f80 g765282 ( .a(n_15921), .b(n_15924), .o(n_16019) );
in01f80 FE_OCP_RBC3516_n_8498 ( .a(n_8498), .o(FE_OCP_RBN3516_n_8498) );
in01f80 g767430 ( .a(n_13397), .o(n_13491) );
in01f80 newInst_1862 ( .a(newNet_1861), .o(newNet_1862) );
in01f80 g749969 ( .a(n_30141), .o(n_30142) );
oa12f80 g770973 ( .a(n_9836), .b(n_10045), .c(n_9905), .o(n_10171) );
in01f80 g754104 ( .a(n_26204), .o(n_26144) );
no02f80 g761504 ( .a(n_18871), .b(n_18870), .o(n_18872) );
in01f80 FE_RC_820_0 ( .a(FE_RN_248_0), .o(n_9087) );
ao12f80 g751497 ( .a(n_28566), .b(n_28467), .c(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n_28701) );
in01f80 g757071 ( .a(n_23282), .o(n_23283) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_6_ ( .ck(newNet_1171), .d(n_4631), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_6_) );
no02f80 g771209 ( .a(n_9262), .b(FE_OCP_RBN2523_n_8951), .o(n_9358) );
ao12f80 g737618 ( .a(n_42294), .b(n_42308), .c(n_42270), .o(n_42400) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_1_ ( .ck(newNet_2759), .d(n_15065), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_) );
in01f80 g738798 ( .a(n_41537), .o(n_41564) );
in01f80 g779817 ( .a(n_1780), .o(n_1452) );
in01f80 newInst_3262 ( .a(newNet_2924), .o(newNet_3262) );
na02f80 g764883 ( .a(n_15543), .b(n_15586), .o(n_15619) );
na02f80 g739375 ( .a(n_40841), .b(n_40882), .o(n_41276) );
oa12f80 g749816 ( .a(n_31344), .b(FE_OCP_RBN3011_n_31117), .c(n_31277), .o(n_31617) );
no02f80 g776095 ( .a(n_4843), .b(n_4842), .o(n_4867) );
in01f80 FE_OCP_RBC3445_n_37945 ( .a(FE_OCP_RBN3442_n_37945), .o(FE_OCP_RBN3445_n_37945) );
no02f80 g748172 ( .a(n_32098), .b(n_32118), .o(n_32208) );
na02f80 g758863 ( .a(n_21437), .b(n_21398), .o(n_21587) );
na02f80 g744245 ( .a(n_46214), .b(n_36852), .o(n_37672) );
na02f80 g737963 ( .a(n_42170), .b(delay_sub_ln23_0_unr29_stage10_stallmux_q), .o(n_42177) );
na02f80 g774875 ( .a(n_6196), .b(FE_OCP_RBN2943_n_5454), .o(n_6205) );
in01f80 g746948 ( .a(n_32941), .o(n_32973) );
na02f80 g776941 ( .a(n_3973), .b(n_47022), .o(n_4149) );
no02f80 g747249 ( .a(FE_OCP_RBN2154_n_32772), .b(FE_OCPN1015_n_32820), .o(n_32815) );
in01f80 g763771 ( .a(n_17367), .o(n_17305) );
ms00f80 cos_out_reg_5_ ( .ck(newNet_3682), .d(n_43695), .o(cos_out_5) );
in01f80 g763216 ( .a(n_17048), .o(n_17049) );
no03m80 FE_RC_1379_0 ( .a(n_26306), .b(n_26217), .c(n_26225), .o(n_26378) );
in01f80 FE_OCPC852_n_694 ( .a(FE_OCPN851_n_694), .o(FE_OCPN852_n_694) );
no02f80 g771619 ( .a(n_9130), .b(n_9070), .o(n_9170) );
na02f80 g778692 ( .a(FE_OCP_RBN2290_n_2438), .b(n_2577), .o(n_2590) );
ao12f80 g768723 ( .a(n_11578), .b(n_11989), .c(n_11716), .o(n_11988) );
na02f80 g757488 ( .a(n_22935), .b(FE_OCP_RBN3819_n_44061), .o(n_22959) );
na02f80 g776991 ( .a(n_5384), .b(n_5355), .o(n_5403) );
in01f80 FE_OCP_RBC3715_n_39913 ( .a(FE_OCP_RBN3053_n_39913), .o(FE_OCP_RBN3715_n_39913) );
ao22s80 g776398 ( .a(FE_OCP_RBN2745_n_47011), .b(FE_OCPN960_n_3951), .c(n_47011), .d(n_4182), .o(n_4429) );
no02f80 g746090 ( .a(n_33831), .b(n_33830), .o(n_33832) );
in01f80 g740219 ( .a(n_40107), .o(n_40064) );
in01f80 newInst_3100 ( .a(newNet_2804), .o(newNet_3100) );
no02f80 g767088 ( .a(n_13606), .b(n_13608), .o(n_13617) );
no02f80 g762204 ( .a(n_18698), .b(n_18443), .o(n_18700) );
no02f80 g781105 ( .a(n_241), .b(n_549), .o(n_240) );
in01f80 FE_OCP_RBC2596_n_25181 ( .a(FE_OCP_RBN2593_n_25181), .o(FE_OCP_RBN2596_n_25181) );
na02f80 g777375 ( .a(n_4675), .b(FE_OFN825_n_5067), .o(n_5247) );
na02f80 g779098 ( .a(n_2005), .b(n_1977), .o(n_2317) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_8_ ( .ck(newNet_994), .d(n_17418), .o(delay_xor_ln21_unr12_stage5_stallmux_q_8_) );
na02f80 g766419 ( .a(n_14102), .b(n_14240), .o(n_14129) );
na02f80 g779246 ( .a(n_1828), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .o(n_1899) );
in01f80 newInst_15 ( .a(newNet_14), .o(newNet_15) );
in01f80 g760043 ( .a(n_21053), .o(n_21051) );
in01f80 g767704 ( .a(n_12898), .o(n_12899) );
no02f80 g766364 ( .a(n_14123), .b(n_13131), .o(n_14162) );
na02f80 g772045 ( .a(n_8710), .b(n_8652), .o(n_8793) );
in01f80 g743589 ( .a(n_37611), .o(n_37612) );
na02f80 g764567 ( .a(n_16007), .b(n_14452), .o(n_16008) );
in01f80 g749915 ( .a(n_30147), .o(n_30148) );
na02f80 g763476 ( .a(n_16880), .b(n_16879), .o(n_16908) );
no02f80 g770186 ( .a(n_10779), .b(n_10584), .o(n_10862) );
na02f80 g747813 ( .a(n_33392), .b(n_33441), .o(n_33413) );
in01f80 newInst_3348 ( .a(newNet_3347), .o(newNet_3348) );
na02f80 g746163 ( .a(n_33623), .b(n_33136), .o(n_33677) );
in01f80 g750761 ( .a(n_29262), .o(n_29296) );
na02f80 g776129 ( .a(n_4660), .b(FE_OCP_RBN2854_n_45462), .o(n_4915) );
na02f80 g760616 ( .a(n_20301), .b(n_19876), .o(n_20356) );
in01f80 g741848 ( .a(n_38495), .o(n_38436) );
no02f80 g771274 ( .a(n_9150), .b(n_9050), .o(n_9298) );
na02f80 g769229 ( .a(FE_OCP_RBN3093_n_11475), .b(n_10935), .o(n_11626) );
in01f80 FE_OCPC3173_n_38799 ( .a(n_38799), .o(FE_OCPN3173_n_38799) );
in01f80 FE_OCP_RBC2338_n_24325 ( .a(n_24325), .o(FE_OCP_RBN2338_n_24325) );
oa22f80 g784338 ( .a(FE_OCP_RBN3075_FE_OFN807_n_46195), .b(n_5913), .c(FE_OFN86_n_46137), .d(n_5906), .o(n_46143) );
in01f80 g749165 ( .a(n_30991), .o(n_31021) );
in01f80 FE_OCPC1384_n_18345 ( .a(FE_OCPN1383_n_18345), .o(FE_OCPN1384_n_18345) );
oa12f80 g739832 ( .a(n_40313), .b(n_40432), .c(n_40242), .o(n_40450) );
in01f80 FE_OCPC1390_n_9220 ( .a(FE_OCPN1389_n_9220), .o(FE_OCPN1390_n_9220) );
na02f80 g736929 ( .a(n_43038), .b(n_42792), .o(n_43087) );
no02f80 g751866 ( .a(n_28217), .b(n_28219), .o(n_28249) );
ao22s80 FE_RC_831_0 ( .a(n_23967), .b(n_24375), .c(n_23968), .d(n_24407), .o(n_24506) );
oa12f80 g764339 ( .a(n_16367), .b(n_16366), .c(n_16365), .o(n_16425) );
in01f80 g759816 ( .a(n_21855), .o(n_21856) );
no02f80 g737911 ( .a(n_42201), .b(n_41921), .o(n_42283) );
no02f80 g752183 ( .a(n_27940), .b(n_26566), .o(n_28068) );
na02f80 g748042 ( .a(n_32966), .b(n_32607), .o(n_33004) );
in01f80 g743724 ( .a(n_37362), .o(n_37363) );
in01f80 fopt782796 ( .a(n_44219), .o(n_44218) );
na02f80 g769366 ( .a(FE_OCPN867_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .o(n_11968) );
ao22s80 g756295 ( .a(n_23949), .b(n_23688), .c(n_24005), .d(n_23687), .o(n_24070) );
no02f80 g777843 ( .a(n_3204), .b(n_2425), .o(n_3205) );
in01f80 g747655 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(n_32171) );
no02f80 g740093 ( .a(n_39801), .b(n_39773), .o(n_39927) );
ao12f80 g746699 ( .a(n_32800), .b(n_33039), .c(n_32833), .o(n_33113) );
na02f80 g753622 ( .a(n_26597), .b(n_26591), .o(n_26669) );
na02f80 g781013 ( .a(sin_out_19), .b(FE_OFN3_n_43918), .o(n_328) );
in01f80 g778426 ( .a(n_2663), .o(n_3532) );
in01f80 g750137 ( .a(n_29832), .o(n_29833) );
in01f80 newInst_1636 ( .a(newNet_1635), .o(newNet_1636) );
na02f80 g769692 ( .a(n_11313), .b(n_11312), .o(n_11317) );
no02f80 FE_RC_3353_0 ( .a(FE_RN_1461_0), .b(FE_RN_1462_0), .o(FE_RN_1463_0) );
in01f80 g748767 ( .a(n_31375), .o(n_31376) );
no02f80 g750331 ( .a(n_30690), .b(n_30689), .o(n_30691) );
no02f80 g776725 ( .a(n_4330), .b(n_4276), .o(n_4499) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_1_ ( .ck(newNet_1936), .d(n_36766), .o(delay_sub_ln21_unr24_stage9_stallmux_q_1_) );
oa22f80 g750997 ( .a(FE_OCP_DRV_N1574_n_28869), .b(n_28913), .c(n_28870), .d(n_28912), .o(n_29892) );
in01f80 g779602 ( .a(n_1703), .o(n_1704) );
in01f80 g771862 ( .a(n_10246), .o(n_10247) );
in01f80 g757398 ( .a(FE_OCPN1020_n_23078), .o(n_22910) );
no02f80 g762069 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n_18505) );
oa22f80 g752477 ( .a(n_27714), .b(n_24059), .c(n_27683), .d(n_27845), .o(n_27737) );
na02f80 g753593 ( .a(n_26753), .b(FE_OCPN1518_n_26752), .o(n_26819) );
na02f80 g756809 ( .a(n_47245), .b(n_23032), .o(n_23439) );
no02f80 g776919 ( .a(n_3849), .b(n_3852), .o(n_3987) );
no02f80 g746577 ( .a(n_34810), .b(n_34547), .o(n_35069) );
na02f80 g754571 ( .a(n_26770), .b(n_26677), .o(n_26790) );
na02f80 g744288 ( .a(n_44180), .b(n_35774), .o(n_35899) );
no02f80 g779445 ( .a(n_1434), .b(n_1400), .o(n_1474) );
na02f80 g753270 ( .a(n_27377), .b(n_26110), .o(n_27462) );
in01f80 FE_OCP_RBC2891_n_10568 ( .a(n_10568), .o(FE_OCP_RBN2891_n_10568) );
oa12f80 g771304 ( .a(n_9310), .b(n_9654), .c(n_9311), .o(n_9884) );
in01f80 g779647 ( .a(n_1482), .o(n_1483) );
in01f80 g770554 ( .a(n_10433), .o(n_10434) );
no02f80 g750439 ( .a(n_29641), .b(n_29590), .o(n_29706) );
oa12f80 g736516 ( .a(n_311), .b(n_43663), .c(FE_OFN3_n_43918), .o(n_43703) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_5_ ( .ck(newNet_552), .d(n_17029), .o(delay_xor_ln22_unr12_stage5_stallmux_q_5_) );
no02f80 g747102 ( .a(n_32927), .b(delay_add_ln22_unr20_stage8_stallmux_q_8_), .o(n_32954) );
na02f80 g748852 ( .a(n_31199), .b(n_31180), .o(n_31328) );
no02f80 g753549 ( .a(n_26694), .b(n_26615), .o(n_26730) );
no02f80 g761929 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .o(n_18549) );
na02f80 g748597 ( .a(n_32723), .b(n_32538), .o(n_33146) );
in01f80 FE_RC_1810_0 ( .a(n_11770), .o(FE_RN_537_0) );
in01f80 FE_OCP_DRV_C3148_n_33225 ( .a(FE_OCP_DRV_N3147_n_33225), .o(FE_OCP_DRV_N3148_n_33225) );
na02f80 g751896 ( .a(n_29040), .b(n_29049), .o(n_29723) );
no02f80 FE_RC_2664_0 ( .a(n_2332), .b(FE_RN_1112_0), .o(FE_RN_1113_0) );
no02f80 FE_RC_1506_0 ( .a(FE_RN_421_0), .b(FE_RN_420_0), .o(FE_RN_422_0) );
no02f80 g754578 ( .a(n_25405), .b(n_25213), .o(n_25466) );
in01f80 g753028 ( .a(n_28336), .o(n_32287) );
in01f80 g754476 ( .a(n_26935), .o(n_26936) );
na02f80 g756747 ( .a(n_23513), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_), .o(n_23571) );
no02f80 g746912 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n_33186) );
no02f80 g742922 ( .a(n_37067), .b(n_37019), .o(n_37506) );
in01f80 FE_RC_1008_0 ( .a(n_17713), .o(FE_RN_292_0) );
na02f80 g752909 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n_27986) );
no02f80 g764694 ( .a(n_15812), .b(n_15810), .o(n_15811) );
in01f80 newInst_3205 ( .a(newNet_2418), .o(newNet_3205) );
no02f80 g778584 ( .a(n_2514), .b(n_2073), .o(n_2530) );
ao22s80 g736637 ( .a(n_43096), .b(n_43069), .c(n_43095), .d(n_43068), .o(n_43191) );
no02f80 g750097 ( .a(n_29857), .b(n_29892), .o(n_29918) );
oa12f80 g752673 ( .a(n_28261), .b(n_28178), .c(n_27923), .o(n_28260) );
na02f80 g763132 ( .a(n_17145), .b(n_17092), .o(n_17294) );
na02f80 g743173 ( .a(n_36930), .b(n_36943), .o(n_37227) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_22_ ( .ck(newNet_3221), .d(n_36468), .o(delay_add_ln22_unr23_stage9_stallmux_q_22_) );
no02f80 g754882 ( .a(n_25453), .b(n_25382), .o(n_25511) );
in01f80 g741257 ( .a(n_39451), .o(n_39452) );
in01f80 newInst_2882 ( .a(newNet_2881), .o(newNet_2882) );
oa12f80 g748192 ( .a(n_31467), .b(n_31424), .c(n_31447), .o(n_31506) );
in01f80 g761171 ( .a(n_19110), .o(n_19111) );
no02f80 g755285 ( .a(n_24900), .b(n_24808), .o(n_24975) );
in01f80 g741558 ( .a(n_38696), .o(n_38697) );
na02f80 g749790 ( .a(n_31282), .b(n_31570), .o(n_31313) );
no02f80 g755029 ( .a(n_25773), .b(n_25772), .o(n_25774) );
in01f80 g780887 ( .a(n_391), .o(n_392) );
na02f80 g777181 ( .a(n_4833), .b(n_4722), .o(n_5859) );
in01f80 g766558 ( .a(n_14023), .o(n_14024) );
in01f80 newInst_752 ( .a(newNet_751), .o(newNet_752) );
na02f80 g774467 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_6854) );
na02f80 g748221 ( .a(FE_OCP_RBN3732_n_31819), .b(n_32076), .o(n_32075) );
na02f80 g753397 ( .a(n_27041), .b(n_27040), .o(n_27125) );
oa12f80 g754136 ( .a(n_26948), .b(n_26947), .c(n_26946), .o(n_27001) );
no02f80 g760533 ( .a(n_20385), .b(n_20384), .o(n_20386) );
no02f80 g751630 ( .a(n_28391), .b(n_28371), .o(n_28372) );
no02f80 g743450 ( .a(n_36630), .b(n_36649), .o(n_36751) );
ao12f80 g748072 ( .a(n_32842), .b(n_32841), .c(n_32840), .o(n_33314) );
in01f80 FE_OCP_RBC2660_n_9292 ( .a(n_9292), .o(FE_OCP_RBN2660_n_9292) );
in01f80 newInst_2044 ( .a(newNet_2043), .o(newNet_2044) );
na02f80 g748637 ( .a(n_31301), .b(n_31308), .o(n_31302) );
na02f80 g753126 ( .a(n_27395), .b(n_27211), .o(n_27423) );
in01f80 FE_OCP_RBC2309_n_29298 ( .a(FE_OCP_RBN2308_n_29298), .o(FE_OCP_RBN2309_n_29298) );
ao12f80 g736680 ( .a(n_43023), .b(n_43028), .c(n_43043), .o(n_43075) );
no02f80 g770702 ( .a(n_9860), .b(n_9173), .o(n_9936) );
oa22f80 g736906 ( .a(n_43242), .b(n_43158), .c(FE_OCPN1247_n_43120), .d(n_46943), .o(n_43577) );
no02f80 g768805 ( .a(n_44859), .b(n_11847), .o(n_12024) );
na02f80 g773972 ( .a(n_6969), .b(n_6968), .o(n_7058) );
in01f80 FE_OCP_RBC3432_n_33664 ( .a(FE_OCP_RBN3431_n_33664), .o(FE_OCP_RBN3432_n_33664) );
na02f80 g772866 ( .a(n_8007), .b(n_8054), .o(n_8125) );
in01f80 g751216 ( .a(n_29818), .o(n_29837) );
na02f80 g780834 ( .a(n_499), .b(n_515), .o(n_649) );
in01f80 g747872 ( .a(n_32216), .o(n_32217) );
in01f80 g775183 ( .a(n_5787), .o(n_5788) );
in01f80 g745417 ( .a(n_35718), .o(n_35719) );
no02f80 g769689 ( .a(n_11268), .b(n_10246), .o(n_11333) );
ao12f80 g778925 ( .a(n_1749), .b(n_2144), .c(n_1743), .o(n_2166) );
no02f80 g738749 ( .a(n_41370), .b(n_41322), .o(n_41376) );
na02f80 g747952 ( .a(n_33125), .b(n_33124), .o(n_33126) );
in01f80 g776320 ( .a(n_4846), .o(n_4847) );
no02f80 g765891 ( .a(n_13659), .b(n_14829), .o(n_14877) );
in01f80 g781350 ( .a(beta_3), .o(n_12) );
no02f80 g770149 ( .a(n_10862), .b(n_10864), .o(n_10865) );
ao12f80 g764636 ( .a(n_15932), .b(n_16450), .c(n_15881), .o(n_16506) );
na02f80 FE_RC_2376_0 ( .a(FE_RN_923_0), .b(n_12119), .o(FE_RN_924_0) );
in01f80 g742210 ( .a(n_38249), .o(n_38250) );
in01f80 g768148 ( .a(FE_OCP_RBN2249_n_13017), .o(n_13916) );
oa12f80 g747755 ( .a(n_31810), .b(n_32000), .c(n_31686), .o(n_32169) );
na02f80 g768365 ( .a(n_12464), .b(delay_add_ln22_unr8_stage4_stallmux_q_13_), .o(n_12512) );
ao12f80 g756332 ( .a(n_23895), .b(n_23930), .c(n_23894), .o(n_25179) );
no02f80 g768534 ( .a(n_12310), .b(n_12227), .o(n_12317) );
in01f80 g780114 ( .a(n_1206), .o(n_1201) );
in01f80 g746688 ( .a(n_34390), .o(n_34388) );
in01f80 g779412 ( .a(n_1565), .o(n_1566) );
in01f80 g743739 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n_36465) );
in01f80 g772231 ( .a(n_8852), .o(n_8900) );
in01f80 g744824 ( .a(n_35102), .o(n_35155) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_26_ ( .ck(newNet_2928), .d(FE_OCP_RBN3140_n_6477), .o(delay_add_ln22_unr5_stage3_stallmux_q_26_) );
na02f80 g756376 ( .a(n_23973), .b(n_23856), .o(n_23999) );
in01f80 newInst_332 ( .a(newNet_331), .o(newNet_332) );
ao12f80 g760315 ( .a(n_20176), .b(n_20835), .c(n_20220), .o(n_20899) );
no02f80 g780012 ( .a(n_1266), .b(n_1027), .o(n_1269) );
ao12f80 g777954 ( .a(n_3091), .b(n_3090), .c(n_3089), .o(n_3717) );
no03m80 FE_RC_1046_0 ( .a(n_32643), .b(FE_RN_305_0), .c(n_32704), .o(n_32721) );
no02f80 g741047 ( .a(n_39081), .b(n_39056), .o(n_39077) );
no02f80 g744266 ( .a(n_44174), .b(n_35569), .o(n_35619) );
in01f80 g746879 ( .a(n_33855), .o(n_33870) );
na02f80 g766312 ( .a(n_14160), .b(n_14201), .o(n_14202) );
in01f80 g753037 ( .a(n_27948), .o(n_28336) );
in01f80 g778153 ( .a(n_2891), .o(n_2875) );
in01f80 g752998 ( .a(n_27427), .o(n_27428) );
na02f80 g779131 ( .a(n_2025), .b(n_1704), .o(n_2051) );
na02f80 g778610 ( .a(n_2388), .b(n_2452), .o(n_2456) );
in01f80 g738177 ( .a(n_42013), .o(n_42710) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_17_ ( .ck(newNet_3431), .d(n_27617), .o(delay_add_ln22_unr17_stage7_stallmux_q_17_) );
na02f80 g742372 ( .a(n_37801), .b(n_37800), .o(n_37810) );
in01f80 newInst_2702 ( .a(newNet_2701), .o(newNet_2702) );
na02f80 g742213 ( .a(n_44877), .b(n_37969), .o(n_37970) );
in01f80 FE_OCP_RBC2477_n_8599 ( .a(n_8599), .o(FE_OCP_RBN2477_n_8599) );
na02f80 g764497 ( .a(n_16573), .b(n_16572), .o(n_16574) );
oa12f80 g738237 ( .a(n_41932), .b(n_41931), .c(n_41930), .o(n_41955) );
no02f80 g742534 ( .a(n_37494), .b(n_37512), .o(n_37578) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_17_ ( .ck(newNet_1331), .d(n_1237), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_17_) );
in01f80 g776401 ( .a(n_4396), .o(n_4388) );
no02f80 g768493 ( .a(n_12336), .b(delay_add_ln22_unr8_stage4_stallmux_q_9_), .o(n_12353) );
in01f80 fopt783918 ( .a(n_27715), .o(n_45619) );
in01f80 g765100 ( .a(n_15420), .o(n_15421) );
na02f80 g755063 ( .a(n_25125), .b(n_25209), .o(n_25333) );
ao12f80 g743708 ( .a(n_35987), .b(n_36372), .c(n_35870), .o(n_36392) );
oa12f80 g747236 ( .a(n_33395), .b(n_33723), .c(n_33421), .o(n_33893) );
na02f80 g763059 ( .a(n_17579), .b(FE_OCP_RBN2139_n_17547), .o(n_17742) );
no02f80 g753923 ( .a(n_26187), .b(n_26212), .o(n_26425) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_22_ ( .ck(newNet_3313), .d(FE_OCP_RBN3113_n_32254), .o(delay_add_ln22_unr20_stage8_stallmux_q_22_) );
no02f80 g759642 ( .a(FE_OCP_RBN1706_n_20616), .b(FE_OCPN1504_n_47257), .o(n_20646) );
no02f80 g762013 ( .a(n_19014), .b(n_47248), .o(n_18338) );
in01f80 g770819 ( .a(n_10251), .o(n_10252) );
no02f80 g737003 ( .a(n_43097), .b(n_42992), .o(n_43464) );
na02f80 FE_RC_3990_0 ( .a(n_29872), .b(FE_RN_1730_0), .o(n_30079) );
na02f80 g741930 ( .a(n_38219), .b(n_38186), .o(n_38220) );
in01f80 g760827 ( .a(n_19685), .o(n_19616) );
ms00f80 cos_out_reg_0_ ( .ck(newNet_3757), .d(n_43154), .o(cos_out_0) );
no02f80 g739474 ( .a(n_40715), .b(n_40714), .o(n_40753) );
na02f80 g757507 ( .a(n_23343), .b(n_23342), .o(n_23344) );
na02f80 g745431 ( .a(FE_OCP_RBN2987_n_35539), .b(n_35526), .o(n_36018) );
na02f80 g753179 ( .a(n_27204), .b(n_25777), .o(n_27420) );
no03m80 g762823 ( .a(n_17726), .b(n_17683), .c(n_17684), .o(n_17727) );
no02f80 g775733 ( .a(n_5300), .b(FE_OCP_RBN2626_n_3848), .o(n_5340) );
in01f80 FE_OCP_RBC2561_n_29819 ( .a(n_29819), .o(FE_OCP_RBN2561_n_29819) );
in01f80 g738663 ( .a(n_41387), .o(n_41425) );
in01f80 newInst_2660 ( .a(newNet_142), .o(newNet_2660) );
no02f80 g772853 ( .a(n_8002), .b(n_8069), .o(n_8070) );
oa12f80 g746742 ( .a(n_32925), .b(n_33066), .c(n_32967), .o(n_33145) );
ao22s80 FE_RC_1255_0 ( .a(n_4968), .b(FE_OCP_RBN2875_n_5082), .c(n_5082), .d(n_4969), .o(n_5221) );
in01f80 FE_OCP_RBC3596_FE_OCPN1243_n_44460 ( .a(FE_OCPN1243_n_44460), .o(FE_OCP_RBN3596_FE_OCPN1243_n_44460) );
no02f80 g767753 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_), .o(n_13204) );
na02f80 g749472 ( .a(n_30455), .b(n_30469), .o(n_30534) );
in01f80 newInst_2195 ( .a(newNet_2194), .o(newNet_2195) );
no02f80 g756414 ( .a(n_23657), .b(n_23775), .o(n_23776) );
na02f80 g773058 ( .a(n_7656), .b(n_7685), .o(n_7754) );
na02f80 g748686 ( .a(n_31207), .b(n_31206), .o(n_31208) );
in01f80 g749251 ( .a(n_30904), .o(n_30926) );
in01f80 g743610 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_18_), .o(n_36503) );
na02f80 g766500 ( .a(n_14060), .b(n_13391), .o(n_14144) );
in01f80 g779514 ( .a(n_1719), .o(n_1720) );
no02f80 g741902 ( .a(n_38172), .b(n_38091), .o(n_38244) );
na02f80 g769882 ( .a(n_11249), .b(n_11152), .o(n_11259) );
na02f80 g749297 ( .a(n_30817), .b(n_30621), .o(n_30841) );
no02f80 g741037 ( .a(n_38966), .b(n_38833), .o(n_39221) );
in01f80 newInst_476 ( .a(newNet_475), .o(newNet_476) );
no02f80 g754819 ( .a(n_25247), .b(n_25246), .o(n_25248) );
oa12f80 g774252 ( .a(n_6624), .b(n_6828), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n_6829) );
na02f80 g741323 ( .a(FE_OCP_RBN3582_n_44944), .b(n_38601), .o(n_39123) );
in01f80 g738962 ( .a(n_41194), .o(n_41215) );
in01f80 newInst_2709 ( .a(newNet_2708), .o(newNet_2709) );
in01f80 newInst_136 ( .a(newNet_135), .o(newNet_136) );
no02f80 g756640 ( .a(n_23558), .b(n_23557), .o(n_23559) );
na02f80 g777723 ( .a(n_3296), .b(n_2566), .o(n_3337) );
in01f80 newInst_1136 ( .a(newNet_1064), .o(newNet_1136) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_8_ ( .ck(newNet_3272), .d(n_31470), .o(delay_add_ln22_unr20_stage8_stallmux_q_8_) );
no02f80 g773179 ( .a(FE_OCP_RBN2228_n_7598), .b(n_7683), .o(n_7684) );
na02f80 g764252 ( .a(n_16393), .b(n_16400), .o(n_16490) );
no02f80 g770967 ( .a(n_9463), .b(n_9582), .o(n_9583) );
in01f80 g771083 ( .a(n_9763), .o(n_9845) );
in01f80 g739964 ( .a(n_39961), .o(n_39962) );
in01f80 g780890 ( .a(n_444), .o(n_445) );
na02f80 g738414 ( .a(n_41699), .b(n_41698), .o(n_41700) );
oa12f80 g778460 ( .a(n_2345), .b(n_2344), .c(n_2343), .o(n_2446) );
oa12f80 g738902 ( .a(n_41271), .b(n_41270), .c(n_41269), .o(n_41299) );
na02f80 g763248 ( .a(n_16918), .b(n_16834), .o(n_17008) );
na02f80 g760252 ( .a(n_20249), .b(n_19262), .o(n_20473) );
no02f80 g746773 ( .a(n_32960), .b(FE_OCP_RBN2167_n_32892), .o(n_32998) );
in01f80 g755792 ( .a(n_25006), .o(n_25007) );
oa22f80 g740120 ( .a(FE_OCP_RBN3056_n_39913), .b(n_39800), .c(FE_OCP_RBN3719_n_39913), .d(n_39817), .o(n_40322) );
na02f80 g741250 ( .a(FE_OCP_RBN2638_n_38806), .b(n_38494), .o(n_38983) );
na02f80 g738950 ( .a(n_41169), .b(n_41168), .o(n_41170) );
in01f80 FE_OCP_DRV_C1557_n_19590 ( .a(n_19590), .o(FE_OCP_DRV_N1557_n_19590) );
oa12f80 g746509 ( .a(n_35159), .b(n_34666), .c(n_34889), .o(n_35508) );
na02f80 g753803 ( .a(n_26374), .b(n_26410), .o(n_26529) );
na02f80 g770878 ( .a(n_9968), .b(n_9716), .o(n_10092) );
in01f80 g740096 ( .a(n_40326), .o(n_40327) );
na02f80 g776995 ( .a(n_3810), .b(n_3886), .o(n_3909) );
oa12f80 g741772 ( .a(n_38424), .b(n_38423), .c(n_38422), .o(n_38907) );
oa12f80 g749891 ( .a(n_31042), .b(n_31065), .c(n_31041), .o(n_31416) );
no02f80 g756159 ( .a(n_24177), .b(n_24203), .o(n_24288) );
in01f80 g742054 ( .a(n_37895), .o(n_37896) );
in01f80 FE_OCP_RBC2793_n_10106 ( .a(n_10106), .o(FE_OCP_RBN2793_n_10106) );
no02f80 g768263 ( .a(n_12673), .b(n_12672), .o(n_12695) );
oa12f80 g736452 ( .a(n_314), .b(n_43724), .c(FE_OFN2_n_43918), .o(n_43767) );
ao12f80 g768843 ( .a(n_12056), .b(n_45685), .c(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .o(n_12456) );
in01f80 newInst_250 ( .a(newNet_249), .o(newNet_250) );
na02f80 g744859 ( .a(n_35034), .b(n_35056), .o(n_35145) );
no02f80 g760968 ( .a(n_19185), .b(FE_OCPN1458_n_18426), .o(n_19280) );
in01f80 g770868 ( .a(n_9898), .o(n_9910) );
oa22f80 g763862 ( .a(n_16699), .b(n_17336), .c(n_16681), .d(n_16339), .o(n_16747) );
oa12f80 g742151 ( .a(FE_OCP_RBN3451_n_37945), .b(n_37556), .c(n_37551), .o(n_38217) );
in01f80 g758198 ( .a(n_22041), .o(n_22042) );
in01f80 newInst_280 ( .a(newNet_279), .o(newNet_280) );
in01f80 g756233 ( .a(n_24742), .o(n_24743) );
in01f80 g760290 ( .a(n_20245), .o(n_20275) );
no02f80 g779603 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .o(n_1703) );
na02f80 g771449 ( .a(n_9186), .b(FE_OCPN901_n_44593), .o(n_9376) );
no02f80 g764199 ( .a(n_16471), .b(FE_OCP_RBN2653_n_14684), .o(n_16535) );
in01f80 newInst_2297 ( .a(newNet_861), .o(newNet_2297) );
in01f80 newInst_61 ( .a(newNet_47), .o(newNet_61) );
na02f80 g753285 ( .a(FE_OCPN964_n_27287), .b(n_26492), .o(n_27409) );
in01f80 g753535 ( .a(n_26788), .o(n_26732) );
no02f80 g755680 ( .a(n_24500), .b(n_23921), .o(n_24566) );
in01f80 g777415 ( .a(n_3705), .o(n_3690) );
na02f80 g776631 ( .a(n_4235), .b(n_4208), .o(n_4355) );
oa22f80 g753860 ( .a(n_27035), .b(n_26575), .c(n_27051), .d(n_26574), .o(n_27092) );
in01f80 g755107 ( .a(n_25205), .o(n_25229) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_29_ ( .ck(newNet_3023), .d(n_1124), .o(delay_add_ln22_unr2_stage2_stallmux_q_29_) );
na02f80 g740733 ( .a(n_39518), .b(n_39537), .o(n_40009) );
na02f80 g736900 ( .a(n_43293), .b(n_43483), .o(n_43581) );
oa12f80 g755185 ( .a(n_25194), .b(n_25660), .c(n_25052), .o(n_25717) );
oa12f80 g755608 ( .a(n_24503), .b(n_24471), .c(n_24502), .o(n_24508) );
oa12f80 g738160 ( .a(n_42002), .b(n_42003), .c(n_42001), .o(n_42542) );
no02f80 g743852 ( .a(n_35832), .b(n_35621), .o(n_35920) );
in01f80 g744945 ( .a(n_35001), .o(n_35684) );
oa22f80 g738616 ( .a(n_41716), .b(n_41124), .c(n_41713), .d(n_41501), .o(n_41893) );
na02f80 g741202 ( .a(n_38870), .b(FE_OCP_RBN2370_n_38545), .o(n_39098) );
in01f80 g742933 ( .a(n_37063), .o(n_37064) );
oa12f80 g762633 ( .a(n_18019), .b(n_18020), .c(n_18018), .o(n_18106) );
na02f80 g759894 ( .a(n_21138), .b(n_21137), .o(n_21139) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_7_ ( .ck(newNet_146), .d(n_46371), .o(delay_xor_ln22_unr9_stage4_stallmux_q_7_) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_13_ ( .ck(newNet_2787), .d(n_16601), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_13_) );
no02f80 g775930 ( .a(n_5085), .b(n_3814), .o(n_5184) );
in01f80 g758440 ( .a(n_23353), .o(n_23466) );
in01f80 FE_OCP_DRV_C1594_n_34494 ( .a(FE_OCP_DRV_N1593_n_34494), .o(FE_OCP_DRV_N1594_n_34494) );
in01f80 newInst_458 ( .a(newNet_63), .o(newNet_458) );
in01f80 FE_OCPC1776_n_18263 ( .a(FE_OCPN1775_n_18263), .o(FE_OCPN1776_n_18263) );
in01f80 g758681 ( .a(n_21962), .o(n_21963) );
in01f80 newInst_1133 ( .a(newNet_1132), .o(newNet_1133) );
in01f80 newInst_1144 ( .a(newNet_1143), .o(newNet_1144) );
in01f80 g775400 ( .a(n_5743), .o(n_5744) );
ao12f80 g763857 ( .a(n_17363), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_15_), .o(n_17989) );
ao22s80 g774635 ( .a(n_6480), .b(n_6308), .c(n_6485), .d(n_6309), .o(n_6557) );
oa22f80 g751626 ( .a(n_28335), .b(n_28265), .c(n_28373), .d(n_28266), .o(n_29571) );
no02f80 g738566 ( .a(n_41685), .b(n_41722), .o(n_41723) );
na02f80 g778978 ( .a(n_2205), .b(n_1126), .o(n_2264) );
na02f80 g781206 ( .a(n_121), .b(n_158), .o(n_159) );
in01f80 fopt783925 ( .a(n_30302), .o(n_45631) );
in01f80 FE_OCPC1030_n_28423 ( .a(FE_OCPN1029_n_28423), .o(FE_OCPN1030_n_28423) );
in01f80 newInst_3675 ( .a(newNet_3674), .o(newNet_3675) );
in01f80 g746437 ( .a(n_33331), .o(n_33429) );
na02f80 g777143 ( .a(n_3653), .b(n_3570), .o(n_3654) );
in01f80 g774126 ( .a(n_6627), .o(n_6589) );
ao12f80 g738199 ( .a(n_41967), .b(n_41966), .c(n_41965), .o(n_41991) );
na02f80 g775008 ( .a(n_6112), .b(n_5897), .o(n_6129) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_20_ ( .ck(newNet_2473), .d(n_32325), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_20_) );
in01f80 fopt782713 ( .a(n_44102), .o(n_44112) );
oa12f80 g749647 ( .a(n_29989), .b(n_30080), .c(n_29962), .o(n_30180) );
na03f80 FE_RC_1261_0 ( .a(n_39061), .b(n_38951), .c(n_39060), .o(n_39062) );
in01f80 g746486 ( .a(n_34553), .o(n_34554) );
na02f80 g773816 ( .a(n_7144), .b(n_7138), .o(n_7139) );
in01f80 g756473 ( .a(n_23790), .o(n_23791) );
in01f80 newInst_1685 ( .a(newNet_1684), .o(newNet_1685) );
na02f80 g756021 ( .a(n_25139), .b(n_25136), .o(n_25254) );
oa12f80 g767707 ( .a(n_13014), .b(n_12823), .c(n_13013), .o(n_13028) );
no02f80 g749203 ( .a(n_30771), .b(n_30681), .o(n_30772) );
no02f80 FE_RC_3957_0 ( .a(FE_RN_1714_0), .b(n_24042), .o(n_24080) );
in01f80 g755838 ( .a(n_24395), .o(n_24422) );
in01f80 FE_RC_1036_0 ( .a(n_23046), .o(FE_RN_298_0) );
no02f80 g784409 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_), .o(n_46221) );
no02f80 g738040 ( .a(n_42137), .b(n_42570), .o(n_42136) );
in01f80 g755458 ( .a(n_24870), .o(n_24850) );
na02f80 g777891 ( .a(n_3117), .b(n_3115), .o(n_4761) );
in01f80 g779491 ( .a(n_1876), .o(n_1877) );
na02f80 g778664 ( .a(n_2235), .b(n_2237), .o(n_2238) );
na02f80 g754509 ( .a(n_26814), .b(n_26832), .o(n_26829) );
no02f80 FE_RC_2054_0 ( .a(FE_RN_694_0), .b(n_27086), .o(n_27276) );
in01f80 FE_OCP_RBC3252_delay_xor_ln22_unr6_stage3_stallmux_q_0_ ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_0_), .o(FE_OCP_RBN3252_delay_xor_ln22_unr6_stage3_stallmux_q_0_) );
in01f80 newInst_2522 ( .a(newNet_690), .o(newNet_2522) );
in01f80 newInst_1998 ( .a(newNet_1997), .o(newNet_1998) );
oa12f80 g772764 ( .a(n_8039), .b(n_8084), .c(n_8140), .o(n_8204) );
in01f80 g778469 ( .a(n_2640), .o(n_2641) );
na02f80 g753002 ( .a(n_27347), .b(FE_OCPN964_n_27287), .o(n_27469) );
no02f80 g760651 ( .a(n_19771), .b(n_19740), .o(n_19878) );
in01f80 FE_OCP_RBC2415_n_8219 ( .a(n_8219), .o(FE_OCP_RBN2415_n_8219) );
oa22f80 g748352 ( .a(FE_OCPN1052_n_31674), .b(n_30350), .c(FE_OCP_RBN3089_FE_OCPN1052_n_31674), .d(n_30324), .o(n_31914) );
in01f80 g765392 ( .a(n_15371), .o(n_15372) );
in01f80 g767980 ( .a(n_12786), .o(n_12787) );
in01f80 FE_OCP_RBC2908_n_26173 ( .a(n_26173), .o(FE_OCP_RBN2908_n_26173) );
in01f80 FE_RC_3686_0 ( .a(n_12393), .o(FE_RN_1619_0) );
na02f80 g745323 ( .a(n_35723), .b(n_35722), .o(n_35807) );
na02f80 g766939 ( .a(n_14487), .b(n_14561), .o(n_15209) );
na02f80 g736491 ( .a(n_43664), .b(n_43333), .o(n_43717) );
in01f80 FE_OCPUNCOC3145_n_21058 ( .a(n_21058), .o(FE_OCPUNCON3145_n_21058) );
in01f80 g778812 ( .a(n_3615), .o(n_3106) );
no02f80 g768043 ( .a(n_12739), .b(n_12256), .o(n_12781) );
no02f80 g784702 ( .a(n_7332), .b(n_47179), .o(n_47180) );
na02f80 g761337 ( .a(n_19983), .b(n_19649), .o(n_19846) );
in01f80 g745082 ( .a(n_34947), .o(n_34919) );
no02f80 g773158 ( .a(FE_OCP_RBN2227_n_7598), .b(n_7702), .o(n_7645) );
in01f80 FE_OCP_RBC2315_n_41420 ( .a(FE_OCP_RBN2313_n_41420), .o(FE_OCP_RBN2315_n_41420) );
no02f80 g755887 ( .a(n_25436), .b(n_25086), .o(n_25493) );
no02f80 g763794 ( .a(n_17363), .b(n_17362), .o(n_17364) );
no02f80 g743095 ( .a(n_36564), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37099) );
no02f80 g780794 ( .a(n_528), .b(n_358), .o(n_425) );
na02f80 g754107 ( .a(n_26077), .b(FE_OCPN1494_n_23398), .o(n_26117) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_9_ ( .ck(newNet_427), .d(n_27843), .o(delay_xor_ln22_unr18_stage7_stallmux_q_9_) );
in01f80 FE_RC_2755_0 ( .a(n_2636), .o(FE_RN_1172_0) );
na02f80 g749941 ( .a(n_30213), .b(FE_OCP_RBN2328_n_29378), .o(n_30242) );
in01f80 g767266 ( .a(n_13570), .o(n_13589) );
in01f80 g738696 ( .a(n_41536), .o(n_41558) );
in01f80 newInst_1479 ( .a(newNet_1478), .o(newNet_1479) );
na02f80 g779339 ( .a(n_1623), .b(n_1622), .o(n_1694) );
in01f80 g777456 ( .a(n_3604), .o(n_3637) );
ao22s80 FE_RC_3770_0 ( .a(FE_RN_1654_0), .b(FE_OCP_RBN2461_n_14273), .c(FE_OCP_RBN2253_n_13017), .d(n_14273), .o(n_14468) );
no02f80 g765560 ( .a(FE_OCPN1054_n_14098), .b(n_15105), .o(n_15127) );
oa12f80 g768707 ( .a(n_12175), .b(n_12174), .c(n_12173), .o(n_13095) );
na02f80 g766541 ( .a(n_13957), .b(FE_OCPN1466_n_13014), .o(n_13997) );
no02f80 g764374 ( .a(n_16231), .b(FE_OCPN3775_n_14730), .o(n_16232) );
in01f80 FE_RC_2741_0 ( .a(n_37662), .o(FE_RN_1163_0) );
in01f80 g753220 ( .a(n_27222), .o(n_27667) );
no02f80 g746092 ( .a(n_35190), .b(n_35160), .o(n_35161) );
no02f80 g738080 ( .a(n_42062), .b(n_42061), .o(n_42063) );
no02f80 g755483 ( .a(n_24694), .b(n_24691), .o(n_24692) );
no02f80 g757206 ( .a(n_44068), .b(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .o(n_23378) );
in01f80 newInst_3643 ( .a(newNet_2995), .o(newNet_3643) );
na02f80 g748413 ( .a(FE_OCPN1052_n_31674), .b(n_30731), .o(n_31760) );
in01f80 g752013 ( .a(n_28877), .o(n_28958) );
no02f80 g780378 ( .a(n_955), .b(n_46055), .o(n_901) );
oa12f80 g773985 ( .a(n_6847), .b(n_6973), .c(n_6910), .o(n_7000) );
in01f80 FE_OCPC851_n_694 ( .a(n_694), .o(FE_OCPN851_n_694) );
na02f80 g757027 ( .a(n_23803), .b(n_23804), .o(n_23833) );
no02f80 g778335 ( .a(n_2604), .b(n_3039), .o(n_2605) );
oa12f80 g742548 ( .a(n_37155), .b(n_37467), .c(n_37350), .o(n_37513) );
na02f80 g743585 ( .a(n_36457), .b(n_36033), .o(n_36471) );
na02f80 g749191 ( .a(n_30738), .b(n_27131), .o(n_30774) );
in01f80 g765108 ( .a(n_16308), .o(n_16309) );
in01f80 g758599 ( .a(n_21950), .o(n_21965) );
no02f80 g779084 ( .a(n_2009), .b(n_2008), .o(n_2010) );
in01f80 g771608 ( .a(n_10296), .o(n_10297) );
na03f80 g746746 ( .a(n_33672), .b(n_34174), .c(n_33653), .o(n_34231) );
in01f80 g770723 ( .a(n_10521), .o(n_10522) );
no02f80 g765210 ( .a(n_15265), .b(n_15339), .o(n_15416) );
na02f80 g781047 ( .a(sin_out_10), .b(FE_OFN3_n_43918), .o(n_327) );
in01f80 newInst_1182 ( .a(newNet_1181), .o(newNet_1182) );
in01f80 g740525 ( .a(n_39689), .o(n_39760) );
ao12f80 g773601 ( .a(n_7329), .b(n_7347), .c(n_7328), .o(n_7402) );
na02f80 g752126 ( .a(FE_OCPN878_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_12_), .o(n_28044) );
oa12f80 g741795 ( .a(n_44031), .b(n_38420), .c(n_38139), .o(n_38446) );
no02f80 g744723 ( .a(n_35123), .b(n_35122), .o(n_35184) );
ao12f80 g774204 ( .a(n_6880), .b(n_6872), .c(delay_xor_ln21_unr6_stage3_stallmux_q_11_), .o(n_7042) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_3_ ( .ck(newNet_1474), .d(n_31689), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_) );
no02f80 g746038 ( .a(n_33878), .b(n_33877), .o(n_33879) );
no02f80 g765301 ( .a(n_15745), .b(n_15873), .o(n_16543) );
in01f80 newInst_2631 ( .a(newNet_1596), .o(newNet_2631) );
in01f80 g752156 ( .a(n_28088), .o(n_28089) );
no02f80 g771930 ( .a(n_8955), .b(n_8925), .o(n_9110) );
in01f80 g772619 ( .a(n_8355), .o(n_8323) );
na02f80 g771661 ( .a(n_8971), .b(n_8920), .o(n_9025) );
na02f80 g736461 ( .a(n_43716), .b(n_43368), .o(n_43764) );
in01f80 g778353 ( .a(n_2647), .o(n_2642) );
ao12f80 g779069 ( .a(n_2014), .b(n_2023), .c(n_2013), .o(n_2056) );
ao12f80 g771479 ( .a(n_7744), .b(n_8878), .c(n_7738), .o(n_8941) );
in01f80 g754674 ( .a(n_27014), .o(n_30584) );
ao22s80 FE_RC_554_0 ( .a(n_30599), .b(n_30220), .c(n_30600), .d(n_30221), .o(n_30697) );
na02f80 g754235 ( .a(n_26909), .b(n_26908), .o(n_26910) );
no02f80 g741004 ( .a(n_39054), .b(n_38973), .o(n_39163) );
in01f80 g742944 ( .a(n_37058), .o(n_37187) );
no02f80 g757605 ( .a(FE_OCP_RBN3823_n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_5_), .o(n_22889) );
in01f80 g769954 ( .a(n_11096), .o(n_11097) );
in01f80 newInst_1439 ( .a(newNet_1159), .o(newNet_1439) );
no02f80 g759759 ( .a(n_20272), .b(n_20237), .o(n_20320) );
in01f80 g776134 ( .a(n_4581), .o(n_4624) );
in01f80 g753164 ( .a(n_27480), .o(n_27481) );
in01f80 g765297 ( .a(n_15923), .o(n_16021) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_13_ ( .ck(newNet_1764), .d(n_22118), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_) );
na02f80 g763830 ( .a(n_17157), .b(n_17257), .o(n_17371) );
in01f80 g761531 ( .a(n_18829), .o(n_18868) );
in01f80 g742860 ( .a(n_37214), .o(n_37195) );
na02f80 g775833 ( .a(n_47002), .b(n_5447), .o(n_5547) );
oa12f80 g772591 ( .a(n_7831), .b(n_8305), .c(n_7858), .o(n_8645) );
ao22s80 g761391 ( .a(n_20086), .b(n_20136), .c(n_19980), .d(n_20135), .o(n_20200) );
no02f80 g761806 ( .a(n_18380), .b(n_18411), .o(n_18564) );
in01f80 g740877 ( .a(n_39237), .o(n_39291) );
ao22s80 g778190 ( .a(n_2756), .b(n_3217), .c(n_2792), .d(n_3178), .o(n_2899) );
no02f80 g767724 ( .a(n_13066), .b(n_13210), .o(n_13284) );
oa12f80 g743177 ( .a(n_36877), .b(n_36876), .c(n_36875), .o(n_37655) );
in01f80 g772309 ( .a(n_8632), .o(n_8653) );
na02f80 g739147 ( .a(n_40990), .b(n_40712), .o(n_40991) );
no02f80 g768809 ( .a(n_11916), .b(n_11560), .o(n_11982) );
no02f80 g756871 ( .a(n_23990), .b(n_23701), .o(n_23866) );
na02f80 g772846 ( .a(n_7970), .b(n_7330), .o(n_8023) );
in01f80 g774495 ( .a(n_6877), .o(n_6939) );
ao12f80 g737483 ( .a(n_42566), .b(n_42554), .c(n_42378), .o(n_42600) );
na02f80 g765888 ( .a(n_13659), .b(n_14829), .o(n_14927) );
no02f80 g779742 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_18_), .o(n_1629) );
na02f80 g738413 ( .a(n_41579), .b(n_41583), .o(n_41845) );
in01f80 g773272 ( .a(n_7802), .o(n_7817) );
in01f80 g739444 ( .a(n_40850), .o(n_40719) );
na02f80 g741309 ( .a(FE_OCP_RBN2548_n_44944), .b(n_38498), .o(n_38902) );
in01f80 g754768 ( .a(FE_OCP_RBN2961_n_26231), .o(n_26856) );
in01f80 g738770 ( .a(n_41369), .o(n_42181) );
in01f80 g751728 ( .a(n_28357), .o(n_28358) );
in01f80 g767860 ( .a(n_13084), .o(n_13069) );
oa12f80 g759725 ( .a(n_21671), .b(n_21599), .c(n_21691), .o(n_21827) );
na02f80 g762927 ( .a(n_17762), .b(delay_add_ln22_unr11_stage5_stallmux_q_7_), .o(n_17865) );
no02f80 FE_RC_2922_0 ( .a(n_27549), .b(n_27598), .o(FE_RN_1271_0) );
in01f80 g737651 ( .a(n_42758), .o(n_42759) );
in01f80 g764473 ( .a(n_16316), .o(n_16361) );
in01f80 newInst_2303 ( .a(newNet_2302), .o(newNet_2303) );
in01f80 g763619 ( .a(n_17502), .o(n_17576) );
in01f80 FE_RC_1615_0 ( .a(n_30345), .o(FE_RN_450_0) );
in01f80 g744615 ( .a(n_35360), .o(n_35361) );
oa22f80 g757784 ( .a(n_22479), .b(n_20231), .c(n_22443), .d(n_22580), .o(n_22535) );
in01f80 g779489 ( .a(n_1472), .o(n_1473) );
oa12f80 g742731 ( .a(n_37440), .b(n_37439), .c(n_37438), .o(n_37912) );
in01f80 g771956 ( .a(n_9308), .o(n_9283) );
in01f80 g746623 ( .a(n_34544), .o(n_34640) );
na02f80 g743013 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n_37074) );
no02f80 g755852 ( .a(n_24251), .b(n_23848), .o(n_24271) );
na02f80 g752494 ( .a(n_27638), .b(n_27561), .o(n_27688) );
na02f80 g778689 ( .a(FE_OCP_RBN2294_n_2438), .b(n_2644), .o(n_2745) );
in01f80 newInst_1026 ( .a(newNet_654), .o(newNet_1026) );
in01f80 newInst_604 ( .a(newNet_385), .o(newNet_604) );
no02f80 g753245 ( .a(n_27083), .b(n_25598), .o(n_27152) );
oa12f80 g781137 ( .a(n_212), .b(n_211), .c(n_210), .o(n_393) );
in01f80 g780264 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_17_), .o(n_1083) );
na02f80 g770983 ( .a(n_9503), .b(n_9363), .o(n_9507) );
no02f80 g776200 ( .a(n_4506), .b(n_4563), .o(n_4611) );
in01f80 newInst_3183 ( .a(newNet_3182), .o(newNet_3183) );
in01f80 FE_OCPC3750_n_44222 ( .a(n_44222), .o(FE_OCPN3750_n_44222) );
na02f80 g764160 ( .a(n_16527), .b(n_16486), .o(n_16559) );
in01f80 drc784098 ( .a(n_45844), .o(n_45845) );
in01f80 g759348 ( .a(n_20919), .o(n_20920) );
na02f80 FE_RC_1709_0 ( .a(n_15648), .b(n_15727), .o(FE_RN_471_0) );
in01f80 FE_OCP_RBC1681_n_33491 ( .a(FE_OCP_RBN1680_n_33491), .o(FE_OCP_RBN1681_n_33491) );
na02f80 g750279 ( .a(n_29785), .b(n_29828), .o(n_29873) );
no02f80 g761282 ( .a(n_19011), .b(FE_OCP_DRV_N1552_n_19010), .o(n_19081) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_20_ ( .ck(newNet_172), .d(n_46347), .o(delay_xor_ln22_unr9_stage4_stallmux_q_20_) );
in01f80 g773196 ( .a(n_7739), .o(n_7807) );
no02f80 g760118 ( .a(FE_OCP_RBN3849_n_20290), .b(n_20125), .o(n_20316) );
oa22f80 FE_RC_762_0 ( .a(FE_OCP_RBN2304_n_7817), .b(FE_OCP_RBN2472_n_8664), .c(FE_OCP_RBN3473_n_7886), .d(n_8664), .o(n_8803) );
no02f80 g761656 ( .a(n_19524), .b(n_19523), .o(n_19525) );
in01f80 FE_OCP_RBC2444_n_42051 ( .a(n_42051), .o(FE_OCP_RBN2444_n_42051) );
na02f80 g779366 ( .a(n_1589), .b(n_1446), .o(n_1592) );
no02f80 g764238 ( .a(n_16493), .b(FE_OCP_RBN1184_n_14638), .o(n_16516) );
na02f80 g771072 ( .a(n_9741), .b(n_9740), .o(n_9800) );
na02f80 g769354 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .o(n_11798) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_13_ ( .ck(newNet_1648), .d(n_27093), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_) );
na02f80 g766261 ( .a(n_14363), .b(n_14376), .o(n_14442) );
no02f80 g778969 ( .a(n_2148), .b(n_1747), .o(n_2151) );
na02f80 g749183 ( .a(n_30801), .b(FE_OCP_RBN2376_n_29480), .o(n_30855) );
in01f80 g781202 ( .a(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_17427) );
no02f80 g757999 ( .a(n_22099), .b(FE_OCP_RBN1724_n_21004), .o(n_22133) );
na02f80 g753760 ( .a(n_44325), .b(n_26409), .o(n_26501) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_31_ ( .ck(newNet_2819), .d(n_12240), .o(delay_add_ln22_unr8_stage4_stallmux_q_31_) );
na02f80 g759907 ( .a(n_21051), .b(n_21819), .o(n_21171) );
in01f80 g769993 ( .a(n_10948), .o(n_11003) );
no02f80 FE_RC_2226_0 ( .a(n_37030), .b(n_37029), .o(FE_RN_808_0) );
in01f80 g772561 ( .a(n_8374), .o(n_8400) );
no02f80 g752511 ( .a(n_27691), .b(n_27667), .o(n_27668) );
no02f80 g771423 ( .a(FE_OCP_RBN2530_n_9044), .b(n_8309), .o(n_9118) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_23_ ( .ck(newNet_714), .d(n_46187), .o(delay_xor_ln21_unr6_stage3_stallmux_q_23_) );
in01f80 g739857 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n_40467) );
no02f80 g784414 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n_46226) );
in01f80 fopt783249 ( .a(n_1863), .o(n_44812) );
in01f80 newInst_2254 ( .a(newNet_2253), .o(newNet_2254) );
no02f80 g752531 ( .a(n_27603), .b(n_27295), .o(n_27624) );
no02f80 g766895 ( .a(n_13878), .b(n_14210), .o(n_14426) );
ao12f80 g766340 ( .a(n_14146), .b(n_14228), .c(n_14230), .o(n_14365) );
in01f80 FE_RC_2048_0 ( .a(n_25625), .o(FE_RN_690_0) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_9_ ( .ck(newNet_2985), .d(n_1129), .o(delay_add_ln22_unr2_stage2_stallmux_q_9_) );
no02f80 g738111 ( .a(n_42059), .b(n_41735), .o(n_42096) );
no02f80 g775120 ( .a(n_5964), .b(n_5925), .o(n_6038) );
no02f80 g738045 ( .a(n_42109), .b(n_42118), .o(n_42151) );
na02f80 g758286 ( .a(FE_OCP_RBN1846_n_22068), .b(n_20555), .o(n_22150) );
na02f80 g773640 ( .a(n_47181), .b(n_6895), .o(n_7393) );
in01f80 FE_OCP_RBC1209_n_16814 ( .a(FE_OCP_RBN1207_n_16814), .o(FE_OCP_RBN1209_n_16814) );
na02f80 g777872 ( .a(n_3220), .b(n_47023), .o(n_3263) );
na02f80 g737374 ( .a(n_42807), .b(n_42626), .o(n_42828) );
na02f80 g738988 ( .a(n_41161), .b(n_41160), .o(n_41162) );
no02f80 g748256 ( .a(FE_OCP_RBN3083_n_31819), .b(n_30465), .o(n_32055) );
na02f80 g743919 ( .a(n_35651), .b(n_35707), .o(n_35708) );
na02f80 g775064 ( .a(n_6049), .b(n_6053), .o(n_6146) );
oa22f80 FE_RC_3367_0 ( .a(n_30708), .b(n_31081), .c(n_27131), .d(n_31026), .o(n_31099) );
ao12f80 g756946 ( .a(n_23933), .b(n_24188), .c(n_23399), .o(n_24414) );
in01f80 newInst_1345 ( .a(newNet_1024), .o(newNet_1345) );
ao12f80 g778745 ( .a(n_1415), .b(n_2225), .c(n_1479), .o(n_2251) );
oa22f80 g759825 ( .a(n_21714), .b(n_21819), .c(n_21691), .d(n_20198), .o(n_21884) );
na02f80 g778268 ( .a(n_2575), .b(n_2325), .o(n_2619) );
no02f80 FE_RC_2746_0 ( .a(n_38927), .b(n_38928), .o(FE_RN_1166_0) );
in01f80 g774863 ( .a(n_6240), .o(n_6222) );
na02f80 g754467 ( .a(n_26938), .b(n_26937), .o(n_26939) );
in01f80 newInst_1409 ( .a(newNet_687), .o(newNet_1409) );
in01f80 g763323 ( .a(n_17382), .o(n_17383) );
in01f80 FE_RC_2826_0 ( .a(n_29494), .o(FE_RN_1213_0) );
in01f80 g745401 ( .a(n_35561), .o(n_35562) );
oa12f80 g765774 ( .a(n_15094), .b(n_15093), .c(n_15092), .o(n_15168) );
in01f80 g738716 ( .a(n_41445), .o(n_41418) );
no02f80 g743288 ( .a(n_36742), .b(n_36710), .o(n_36757) );
in01f80 newInst_272 ( .a(newNet_271), .o(newNet_272) );
no02f80 g745063 ( .a(n_34858), .b(n_34562), .o(n_34860) );
na02f80 g773106 ( .a(n_8031), .b(n_8030), .o(n_8032) );
no02f80 g748077 ( .a(n_32865), .b(n_32864), .o(n_32866) );
na02f80 g778473 ( .a(n_2628), .b(delay_add_ln22_unr2_stage2_stallmux_q_25_), .o(n_2656) );
no02f80 g764590 ( .a(n_15816), .b(FE_OCP_RBN2803_n_15706), .o(n_16866) );
no02f80 g765852 ( .a(n_14883), .b(n_14858), .o(n_14978) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_17_ ( .ck(newNet_180), .d(n_46352), .o(delay_xor_ln22_unr9_stage4_stallmux_q_17_) );
oa12f80 g759435 ( .a(n_21699), .b(n_21714), .c(n_21819), .o(n_21888) );
oa12f80 g778007 ( .a(n_2970), .b(n_2969), .c(n_3013), .o(n_3580) );
oa12f80 g748946 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32586) );
no02f80 g746713 ( .a(n_34252), .b(n_34251), .o(n_34253) );
in01f80 newInst_400 ( .a(newNet_399), .o(newNet_400) );
no02f80 g749837 ( .a(FE_OCP_RBN3012_n_31117), .b(n_31171), .o(n_31224) );
in01f80 newInst_1009 ( .a(newNet_1008), .o(newNet_1009) );
ao22s80 g767659 ( .a(n_12865), .b(n_12800), .c(n_12754), .d(n_14003), .o(n_12949) );
no02f80 g772516 ( .a(n_8431), .b(n_8430), .o(n_8432) );
no02f80 g763902 ( .a(n_16591), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17106) );
in01f80 newInst_3692 ( .a(newNet_3691), .o(newNet_3692) );
na02f80 g748215 ( .a(n_32750), .b(n_32533), .o(n_32768) );
oa12f80 g754472 ( .a(n_25323), .b(n_25566), .c(n_25231), .o(n_25632) );
na02f80 FE_RC_2547_0 ( .a(FE_RN_1043_0), .b(FE_RN_1039_0), .o(n_39290) );
in01f80 g768813 ( .a(n_12060), .o(n_12131) );
na02f80 g774870 ( .a(n_6178), .b(n_6119), .o(n_6224) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_4_ ( .ck(newNet_1689), .d(n_21931), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_4_) );
in01f80 g758953 ( .a(n_21361), .o(n_21362) );
na02f80 g761865 ( .a(n_18373), .b(n_18372), .o(n_18407) );
no02f80 g750863 ( .a(n_29063), .b(n_28683), .o(n_29092) );
na02f80 g747838 ( .a(n_33571), .b(n_33720), .o(n_33738) );
no02f80 g766476 ( .a(n_14030), .b(n_14067), .o(n_14149) );
na02f80 g771156 ( .a(n_9793), .b(n_9464), .o(n_9883) );
na02f80 FE_RC_2774_0 ( .a(FE_RN_1181_0), .b(n_8953), .o(FE_RN_1182_0) );
in01f80 FE_RC_3642_0 ( .a(n_31082), .o(FE_RN_1598_0) );
in01f80 g742011 ( .a(n_38183), .o(n_38184) );
in01f80 FE_OCP_RBC3114_n_6379 ( .a(n_6379), .o(FE_OCP_RBN3114_n_6379) );
na03f80 g743230 ( .a(n_38022), .b(n_38093), .c(n_38020), .o(n_38094) );
ao12f80 g757181 ( .a(n_23169), .b(n_23189), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n_23216) );
no02f80 FE_RC_2059_0 ( .a(n_24992), .b(FE_RN_697_0), .o(n_25042) );
in01f80 FE_OCPC887_n_42367 ( .a(FE_OCPN886_n_42367), .o(FE_OCPN887_n_42367) );
na02f80 g743870 ( .a(n_35627), .b(n_35519), .o(n_35673) );
in01f80 newInst_557 ( .a(newNet_556), .o(newNet_557) );
ao12f80 g766839 ( .a(n_13043), .b(n_13633), .c(n_13015), .o(n_13645) );
in01f80 g778132 ( .a(n_2957), .o(n_2958) );
oa12f80 g762056 ( .a(n_18114), .b(n_18196), .c(n_18078), .o(n_18248) );
in01f80 FE_OCP_RBC1367_n_20763 ( .a(n_20763), .o(FE_OCP_RBN1367_n_20763) );
in01f80 g745824 ( .a(n_34201), .o(n_34176) );
ao12f80 g746732 ( .a(n_34173), .b(n_34172), .c(n_34171), .o(n_34738) );
in01f80 newInst_2945 ( .a(newNet_2944), .o(newNet_2945) );
in01f80 newInst_990 ( .a(newNet_989), .o(newNet_990) );
no02f80 g761275 ( .a(n_20036), .b(n_19845), .o(n_19984) );
in01f80 g738647 ( .a(FE_OCP_RBN2313_n_41420), .o(n_41582) );
in01f80 newInst_2459 ( .a(newNet_2111), .o(newNet_2459) );
in01f80 newInst_3752 ( .a(newNet_2918), .o(newNet_3752) );
na02f80 g761925 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n_18511) );
no02f80 g736860 ( .a(n_43504), .b(n_43449), .o(n_43615) );
na02f80 g763669 ( .a(n_17614), .b(n_17468), .o(n_17539) );
na02f80 g769611 ( .a(n_11363), .b(n_11236), .o(n_11408) );
oa12f80 g780734 ( .a(n_606), .b(n_605), .c(n_604), .o(n_773) );
na02f80 g770541 ( .a(n_10359), .b(n_10396), .o(n_10494) );
no02f80 FE_RC_2794_0 ( .a(FE_RN_1193_0), .b(n_14096), .o(FE_RN_1194_0) );
no02f80 g743308 ( .a(n_36673), .b(n_36750), .o(n_36742) );
no02f80 g744297 ( .a(FE_OCP_RBN2902_n_44174), .b(n_34999), .o(n_35900) );
no02f80 g745166 ( .a(n_34542), .b(n_34193), .o(n_34604) );
in01f80 newInst_3529 ( .a(newNet_769), .o(newNet_3529) );
no02f80 g751696 ( .a(n_28391), .b(n_28369), .o(n_28370) );
no02f80 g764831 ( .a(n_15561), .b(n_15099), .o(n_15625) );
oa12f80 g784610 ( .a(n_42904), .b(n_42881), .c(n_42760), .o(n_46938) );
no02f80 g736660 ( .a(n_43372), .b(n_43166), .o(n_43373) );
no02f80 FE_RC_2854_0 ( .a(FE_RN_1228_0), .b(FE_RN_1229_0), .o(n_14286) );
oa12f80 g756367 ( .a(n_23796), .b(n_23795), .c(n_23794), .o(n_23890) );
in01f80 g761724 ( .a(n_19369), .o(n_19370) );
no02f80 g768131 ( .a(n_12663), .b(n_12281), .o(n_12679) );
oa12f80 g777856 ( .a(n_2413), .b(n_3120), .c(FE_OCP_RBN2319_n_2367), .o(n_3222) );
in01f80 newInst_859 ( .a(newNet_560), .o(newNet_859) );
no02f80 g745626 ( .a(n_34286), .b(FE_OCP_RBN2262_n_33691), .o(n_34531) );
oa12f80 g753332 ( .a(n_26907), .b(n_27613), .c(n_26856), .o(n_27627) );
in01f80 newInst_890 ( .a(newNet_371), .o(newNet_890) );
na02f80 g764581 ( .a(n_16544), .b(n_16543), .o(n_16545) );
no02f80 g759084 ( .a(n_21388), .b(n_21423), .o(n_21571) );
in01f80 g762429 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_18_), .o(n_18008) );
no02f80 FE_RC_2697_0 ( .a(FE_RN_1130_0), .b(n_8774), .o(FE_RN_1131_0) );
oa12f80 g759153 ( .a(n_21417), .b(n_21416), .c(n_21415), .o(n_21486) );
na02f80 g760668 ( .a(n_20277), .b(n_19829), .o(n_20301) );
in01f80 g738345 ( .a(n_41816), .o(n_41862) );
no02f80 g750685 ( .a(n_29232), .b(n_28672), .o(n_29281) );
in01f80 g752847 ( .a(n_27058), .o(n_27076) );
no02f80 g741726 ( .a(n_38907), .b(n_38908), .o(n_38518) );
no02f80 g742497 ( .a(n_37563), .b(n_36938), .o(n_37609) );
in01f80 g745386 ( .a(n_36080), .o(n_36081) );
no02f80 g759777 ( .a(n_21795), .b(n_21298), .o(n_22179) );
na02f80 g751783 ( .a(n_28254), .b(n_27917), .o(n_28309) );
in01f80 newInst_2116 ( .a(newNet_1767), .o(newNet_2116) );
ao12f80 g770706 ( .a(n_9933), .b(FE_OCP_RBN2791_n_9910), .c(n_10017), .o(n_10062) );
na02f80 g737558 ( .a(n_42400), .b(n_42412), .o(n_42453) );
oa12f80 g758604 ( .a(n_21692), .b(n_22431), .c(n_21748), .o(n_22527) );
in01f80 g771787 ( .a(n_8891), .o(n_8934) );
na03f80 FE_RC_349_0 ( .a(FE_RN_32_0), .b(n_11695), .c(n_12026), .o(n_12106) );
no02f80 g776549 ( .a(n_4131), .b(n_4073), .o(n_4074) );
na02f80 g780605 ( .a(n_694), .b(n_701), .o(n_710) );
na02f80 g737529 ( .a(n_42337), .b(n_42253), .o(n_42379) );
no02f80 g757047 ( .a(n_23616), .b(n_22882), .o(n_23703) );
no02f80 g765905 ( .a(n_14753), .b(n_14606), .o(n_14891) );
in01f80 newInst_507 ( .a(newNet_506), .o(newNet_507) );
in01f80 g768953 ( .a(n_11778), .o(n_11725) );
no02f80 FE_RC_1783_0 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_15_), .b(n_28025), .o(FE_RN_521_0) );
no02f80 g777178 ( .a(n_4622), .b(n_4921), .o(n_5665) );
no02f80 g757741 ( .a(n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_0_), .o(n_22560) );
ao12f80 g758158 ( .a(n_22697), .b(FE_OCP_RBN2047_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n_23091) );
in01f80 FE_OCP_RBC2960_n_26231 ( .a(FE_OCP_RBN2956_n_26231), .o(FE_OCP_RBN2960_n_26231) );
no02f80 g761911 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_29_), .o(n_18820) );
in01f80 g763178 ( .a(FE_OCPN1456_n_18860), .o(n_18919) );
na02f80 g740899 ( .a(n_44309), .b(n_39361), .o(n_39428) );
na02f80 g748182 ( .a(n_47274), .b(n_32017), .o(n_32124) );
in01f80 g767073 ( .a(n_13669), .o(n_13670) );
in01f80 g740576 ( .a(n_39643), .o(n_39644) );
oa12f80 g754351 ( .a(n_26942), .b(n_26941), .c(n_26940), .o(n_26999) );
in01f80 FE_OCP_RBC2506_n_13896 ( .a(FE_OCP_RBN2501_n_13896), .o(FE_OCP_RBN2506_n_13896) );
in01f80 g754140 ( .a(n_26068), .o(n_26028) );
na02f80 g765415 ( .a(n_15181), .b(n_15143), .o(n_15294) );
no02f80 g778240 ( .a(n_47025), .b(n_2766), .o(n_2777) );
no02f80 g744468 ( .a(n_35483), .b(FE_OCP_DRV_N1580_n_35482), .o(n_35490) );
ao12f80 g773598 ( .a(n_7394), .b(n_7393), .c(n_7392), .o(n_7923) );
in01f80 FE_OCPC1424_delay_sub_ln23_0_unr21_stage8_stallmux_q ( .a(FE_OCPN1423_delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q) );
na02f80 g763843 ( .a(n_16645), .b(FE_OCP_RBN3608_n_14905), .o(n_16708) );
na02f80 g778571 ( .a(n_2422), .b(n_3245), .o(n_2503) );
in01f80 g761292 ( .a(n_20010), .o(n_20051) );
in01f80 FE_OCP_RBC2525_n_24902 ( .a(n_24902), .o(FE_OCP_RBN2525_n_24902) );
ao12f80 g780720 ( .a(n_441), .b(n_619), .c(n_567), .o(n_622) );
na02f80 g748300 ( .a(n_31824), .b(n_31897), .o(n_31919) );
no02f80 g768845 ( .a(n_11823), .b(n_11915), .o(n_11916) );
in01f80 newInst_2191 ( .a(newNet_2190), .o(newNet_2191) );
na02f80 g778215 ( .a(n_2772), .b(n_2726), .o(n_2864) );
no02f80 g770939 ( .a(n_9890), .b(n_9685), .o(n_10013) );
na02f80 g752824 ( .a(n_27400), .b(FE_OCP_RBN2853_n_26169), .o(n_27432) );
no02f80 g749686 ( .a(n_31191), .b(n_31114), .o(n_31259) );
oa22f80 FE_RC_1550_0 ( .a(n_41997), .b(n_41779), .c(n_41780), .d(n_41996), .o(n_42051) );
in01f80 g751260 ( .a(n_29800), .o(n_29782) );
no02f80 g778728 ( .a(n_2215), .b(n_2250), .o(n_2269) );
na02f80 g768885 ( .a(n_11787), .b(n_11543), .o(n_11929) );
in01f80 g750280 ( .a(n_29826), .o(n_29827) );
in01f80 newInst_3405 ( .a(newNet_1768), .o(newNet_3405) );
in01f80 g739094 ( .a(n_41447), .o(n_41062) );
no02f80 g756340 ( .a(n_24455), .b(n_24454), .o(n_24456) );
in01f80 g774249 ( .a(n_7077), .o(n_7078) );
oa22f80 FE_RC_1258_0 ( .a(FE_OCP_RBN2820_n_4872), .b(n_5122), .c(n_5121), .d(n_4900), .o(n_5300) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_9_ ( .ck(newNet_2504), .d(n_27029), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_9_) );
no02f80 g740408 ( .a(FE_OCP_RBN3027_n_39942), .b(n_39989), .o(n_40057) );
in01f80 newInst_744 ( .a(newNet_743), .o(newNet_744) );
no02f80 g743056 ( .a(n_36152), .b(n_46254), .o(n_37014) );
na02f80 g759977 ( .a(n_21102), .b(n_21101), .o(n_21103) );
in01f80 g767048 ( .a(n_13895), .o(n_13876) );
in01f80 newInst_2324 ( .a(newNet_2323), .o(newNet_2324) );
na02f80 g778604 ( .a(n_2701), .b(n_2643), .o(n_3305) );
no02f80 FE_RC_2649_0 ( .a(n_12097), .b(FE_RN_1105_0), .o(n_12292) );
ao12f80 g739258 ( .a(n_40750), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n_41099) );
in01f80 g753914 ( .a(n_26291), .o(n_27210) );
in01f80 newInst_441 ( .a(newNet_440), .o(newNet_441) );
in01f80 g740390 ( .a(n_39934), .o(n_40313) );
in01f80 newInst_1162 ( .a(newNet_146), .o(newNet_1162) );
in01f80 g779398 ( .a(n_1662), .o(n_1604) );
ao22s80 FE_RC_4067_0 ( .a(FE_RN_1769_0), .b(n_26516), .c(n_26564), .d(FE_RN_1770_0), .o(n_26721) );
no02f80 g739999 ( .a(n_40255), .b(n_40104), .o(n_40295) );
in01f80 FE_OCP_RBC1379_n_20732 ( .a(n_20732), .o(FE_OCP_RBN1379_n_20732) );
oa12f80 g738327 ( .a(n_41819), .b(n_41818), .c(n_41817), .o(n_41915) );
no02f80 g754492 ( .a(n_26611), .b(n_26577), .o(n_26645) );
in01f80 newInst_1527 ( .a(newNet_1526), .o(newNet_1527) );
na02f80 g769980 ( .a(n_11019), .b(n_10926), .o(n_11126) );
na02f80 g777786 ( .a(n_3293), .b(n_3105), .o(n_3294) );
na02f80 g771710 ( .a(n_9327), .b(n_9228), .o(n_9387) );
na03f80 FE_RC_1911_0 ( .a(n_33216), .b(n_33609), .c(n_33610), .o(n_33636) );
na02f80 g743038 ( .a(n_37096), .b(n_37095), .o(n_37521) );
in01f80 newInst_627 ( .a(newNet_434), .o(newNet_627) );
na02f80 g771819 ( .a(n_9431), .b(n_9480), .o(n_9481) );
no02f80 g764428 ( .a(n_16197), .b(n_14524), .o(n_16199) );
na02f80 g779276 ( .a(n_1728), .b(delay_add_ln22_unr2_stage2_stallmux_q_6_), .o(n_1815) );
in01f80 newInst_1384 ( .a(newNet_1383), .o(newNet_1384) );
ao12f80 g777737 ( .a(n_3319), .b(n_3318), .c(n_3317), .o(n_3320) );
in01f80 newInst_2055 ( .a(newNet_623), .o(newNet_2055) );
na02f80 g770072 ( .a(n_10792), .b(n_10763), .o(n_10831) );
no02f80 g777063 ( .a(n_5191), .b(n_5188), .o(n_5356) );
in01f80 g759000 ( .a(n_21605), .o(n_21700) );
na02f80 g751726 ( .a(n_28334), .b(n_28043), .o(n_28359) );
no02f80 g766085 ( .a(n_14631), .b(n_14604), .o(n_14709) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_9_ ( .ck(newNet_687), .d(n_46152), .o(delay_xor_ln21_unr6_stage3_stallmux_q_9_) );
in01f80 g772406 ( .a(n_8521), .o(n_8522) );
no02f80 g754526 ( .a(n_26573), .b(n_26541), .o(n_26714) );
in01f80 g737956 ( .a(n_42187), .o(n_42205) );
na02f80 g778207 ( .a(n_2856), .b(n_2799), .o(n_2861) );
oa12f80 g739050 ( .a(n_41132), .b(n_41131), .c(n_41130), .o(n_41175) );
no02f80 g755133 ( .a(n_25373), .b(n_24451), .o(n_25535) );
oa22f80 g740118 ( .a(FE_OCP_RBN3718_n_39913), .b(n_39550), .c(FE_OCP_RBN3719_n_39913), .d(n_39551), .o(n_40221) );
na02f80 g742196 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38251), .o(n_38253) );
in01f80 g778752 ( .a(n_2473), .o(n_3023) );
in01f80 newInst_171 ( .a(newNet_170), .o(newNet_171) );
na02f80 g768794 ( .a(n_12062), .b(n_12061), .o(n_12179) );
na02f80 g762343 ( .a(n_18421), .b(n_18418), .o(n_18451) );
in01f80 g770344 ( .a(n_10746), .o(n_10747) );
in01f80 g777440 ( .a(n_3912), .o(n_3951) );
na02f80 g739664 ( .a(n_40537), .b(n_40249), .o(n_40557) );
na02f80 g761207 ( .a(n_19832), .b(n_19876), .o(n_20353) );
na02f80 g775047 ( .a(n_6077), .b(n_5930), .o(n_6147) );
in01f80 g774307 ( .a(n_6560), .o(n_6876) );
in01f80 FE_OCP_RBC1171_n_13858 ( .a(n_13858), .o(FE_OCP_RBN1171_n_13858) );
na02f80 g746274 ( .a(n_33589), .b(n_33588), .o(n_33590) );
oa22f80 g772425 ( .a(n_8449), .b(FE_OCP_RBN2373_n_8221), .c(FE_OCP_RBN2374_n_8221), .d(n_8448), .o(n_8571) );
in01f80 FE_OCP_RBC1706_n_20616 ( .a(n_20616), .o(FE_OCP_RBN1706_n_20616) );
in01f80 g780535 ( .a(n_1059), .o(n_1060) );
in01f80 newInst_1629 ( .a(newNet_200), .o(newNet_1629) );
na02f80 g767379 ( .a(n_13585), .b(n_13584), .o(n_13586) );
oa12f80 g757768 ( .a(n_23093), .b(n_23092), .c(n_23091), .o(n_23800) );
no02f80 g777276 ( .a(n_4875), .b(FE_OFN825_n_5067), .o(n_5111) );
ao12f80 g761856 ( .a(n_18995), .b(n_18994), .c(n_18993), .o(n_19677) );
in01f80 g762709 ( .a(n_18231), .o(n_18232) );
in01f80 g765987 ( .a(n_14746), .o(n_14747) );
na03f80 FE_RC_3245_0 ( .a(n_10665), .b(n_10624), .c(n_10598), .o(n_10666) );
no02f80 g737747 ( .a(n_42284), .b(n_42277), .o(n_42330) );
in01f80 g758173 ( .a(n_22153), .o(n_22196) );
no02f80 g758935 ( .a(n_21394), .b(n_45026), .o(n_21429) );
no02f80 g776293 ( .a(n_4568), .b(n_4468), .o(n_4536) );
na02f80 g751473 ( .a(n_28491), .b(n_28547), .o(n_28569) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_30_ ( .ck(newNet_3013), .d(FE_OFN27_n_1142), .o(delay_add_ln22_unr2_stage2_stallmux_q_30_) );
na02f80 g753583 ( .a(n_26697), .b(n_26301), .o(n_26756) );
oa12f80 g756427 ( .a(n_24115), .b(n_24114), .c(n_24113), .o(n_24957) );
in01f80 g759384 ( .a(n_20804), .o(n_20862) );
no02f80 g769718 ( .a(n_11201), .b(n_11230), .o(n_11231) );
in01f80 g741197 ( .a(n_38985), .o(n_39103) );
in01f80 FE_RC_4250_0 ( .a(n_26824), .o(FE_RN_1870_0) );
no02f80 g761327 ( .a(n_20197), .b(n_20234), .o(n_20927) );
in01f80 newInst_2772 ( .a(newNet_2771), .o(newNet_2772) );
in01f80 newInst_643 ( .a(newNet_642), .o(newNet_643) );
na02f80 g745518 ( .a(n_34651), .b(n_34650), .o(n_34652) );
na02f80 g744932 ( .a(n_34835), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34883) );
in01f80 newInst_145 ( .a(newNet_144), .o(newNet_145) );
na02f80 g742980 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_10_), .o(n_37006) );
na02f80 g744152 ( .a(n_35856), .b(n_35897), .o(n_35898) );
in01f80 g749965 ( .a(n_30012), .o(n_30013) );
in01f80 newInst_2407 ( .a(newNet_2406), .o(newNet_2407) );
in01f80 g778261 ( .a(n_2918), .o(n_2919) );
na02f80 g753239 ( .a(n_27110), .b(n_27217), .o(n_27218) );
no02f80 g772681 ( .a(FE_OCP_RBN2383_n_8342), .b(n_8300), .o(n_8315) );
oa22f80 FE_RC_3316_0 ( .a(n_17869), .b(n_17907), .c(FE_RN_1459_0), .d(n_17908), .o(n_18038) );
oa12f80 g762954 ( .a(n_17960), .b(n_17959), .c(n_17958), .o(n_18688) );
oa12f80 g745149 ( .a(n_34605), .b(n_34604), .c(n_34603), .o(n_34677) );
in01f80 newInst_1397 ( .a(newNet_1396), .o(newNet_1397) );
in01f80 g759770 ( .a(n_20754), .o(n_20755) );
no02f80 FE_RC_3001_0 ( .a(FE_RN_1313_0), .b(FE_OCP_RBN3094_n_11475), .o(n_11560) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_10_ ( .ck(newNet_760), .d(n_46160), .o(delay_xor_ln21_unr6_stage3_stallmux_q_10_) );
oa22f80 g745787 ( .a(n_44112), .b(n_34206), .c(n_44102), .d(n_34224), .o(n_34445) );
no02f80 g761700 ( .a(n_18714), .b(n_18605), .o(n_18750) );
na02f80 g755139 ( .a(n_25373), .b(n_24555), .o(n_25582) );
in01f80 newInst_3354 ( .a(newNet_3353), .o(newNet_3354) );
in01f80 newInst_3631 ( .a(newNet_3630), .o(newNet_3631) );
no02f80 g738976 ( .a(n_41155), .b(n_40993), .o(n_41244) );
ao12f80 g741501 ( .a(n_38757), .b(n_38756), .c(n_38755), .o(n_38786) );
in01f80 g747245 ( .a(n_32695), .o(n_32696) );
na02f80 g753859 ( .a(n_27054), .b(n_27066), .o(n_27093) );
in01f80 newInst_1233 ( .a(newNet_652), .o(newNet_1233) );
na02f80 g762903 ( .a(FE_OCPN1506_n_17680), .b(n_17624), .o(n_17801) );
na02f80 g770678 ( .a(n_10072), .b(n_44464), .o(n_10264) );
in01f80 FE_OCP_RBC2571_n_29922 ( .a(n_29857), .o(FE_OCP_RBN2571_n_29922) );
na02f80 g738030 ( .a(n_42160), .b(n_42569), .o(n_42161) );
in01f80 g739674 ( .a(n_40593), .o(n_40584) );
na02f80 g750401 ( .a(n_29609), .b(n_29633), .o(n_29687) );
na02f80 g752540 ( .a(n_27620), .b(n_27509), .o(n_27638) );
in01f80 g769579 ( .a(n_11494), .o(n_11463) );
in01f80 FE_RC_3997_0 ( .a(FE_RN_1734_0), .o(FE_RN_1733_0) );
in01f80 g750129 ( .a(n_30421), .o(n_30422) );
na02f80 FE_RC_2918_0 ( .a(n_24446), .b(n_24373), .o(FE_RN_1270_0) );
no02f80 g758164 ( .a(n_44267), .b(n_21339), .o(n_22221) );
in01f80 newInst_247 ( .a(newNet_246), .o(newNet_247) );
na02f80 g738945 ( .a(n_41246), .b(n_41026), .o(n_41283) );
oa12f80 g782644 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_36991), .c(n_36951), .o(n_44038) );
in01f80 g755083 ( .a(n_25691), .o(n_25692) );
no02f80 g744470 ( .a(n_35448), .b(n_35283), .o(n_35468) );
in01f80 FE_RC_3859_0 ( .a(n_31103), .o(FE_RN_1685_0) );
in01f80 g770334 ( .a(n_10748), .o(n_10749) );
ao12f80 g774273 ( .a(n_6391), .b(n_44711), .c(n_6291), .o(n_6503) );
na02f80 g736882 ( .a(n_43430), .b(n_43499), .o(n_43599) );
in01f80 g738109 ( .a(n_42158), .o(n_42124) );
in01f80 newInst_1037 ( .a(newNet_1036), .o(newNet_1037) );
no02f80 g776382 ( .a(n_4543), .b(n_4445), .o(n_4604) );
no02f80 g772492 ( .a(n_8649), .b(n_8648), .o(n_8650) );
in01f80 g736326 ( .a(n_43885), .o(n_43871) );
oa22f80 g784548 ( .a(n_11490), .b(FE_OFN801_n_46285), .c(n_11409), .d(FE_OCP_RBN3043_n_46337), .o(n_46369) );
oa12f80 g751805 ( .a(n_28946), .b(n_28882), .c(n_28836), .o(n_28960) );
oa22f80 FE_RC_443_0 ( .a(n_17584), .b(n_17723), .c(n_17753), .d(n_45472), .o(n_17770) );
oa12f80 g749055 ( .a(n_31387), .b(n_32227), .c(n_31411), .o(n_32272) );
oa12f80 g747857 ( .a(n_33315), .b(n_33310), .c(n_33281), .o(n_33334) );
in01f80 g758470 ( .a(FE_OFN738_n_22641), .o(n_25824) );
na02f80 g764734 ( .a(n_15800), .b(n_15763), .o(n_15895) );
in01f80 g780673 ( .a(n_679), .o(n_694) );
in01f80 FE_RC_1878_0 ( .a(delay_xor_ln22_unr9_stage4_stallmux_q_3_), .o(FE_RN_582_0) );
in01f80 g746473 ( .a(n_35187), .o(n_35188) );
no03m80 g774081 ( .a(n_6708), .b(n_6734), .c(n_6600), .o(n_6760) );
na02f80 g741174 ( .a(n_38847), .b(n_38507), .o(n_38951) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_3_ ( .ck(newNet_886), .d(n_32288), .o(delay_xor_ln21_unr21_stage8_stallmux_q_3_) );
in01f80 g769044 ( .a(n_11693), .o(n_11955) );
in01f80 newInst_2984 ( .a(newNet_2983), .o(newNet_2984) );
in01f80 g754214 ( .a(n_26004), .o(n_25971) );
na02f80 g767925 ( .a(n_12818), .b(n_12496), .o(n_12921) );
ao22s80 FE_RC_546_0 ( .a(n_23844), .b(n_24308), .c(n_23845), .d(n_24307), .o(n_24421) );
in01f80 g741512 ( .a(n_38734), .o(n_38735) );
in01f80 g759787 ( .a(n_21776), .o(n_21777) );
in01f80 FE_OCP_RBC2690_FE_OCPN843_n_3912 ( .a(FE_OCPN843_n_3912), .o(FE_OCP_RBN2690_FE_OCPN843_n_3912) );
in01f80 g738499 ( .a(n_41786), .o(n_41787) );
in01f80 g753652 ( .a(n_26652), .o(n_26653) );
in01f80 g763909 ( .a(n_17359), .o(n_17300) );
no02f80 g772882 ( .a(n_7894), .b(n_7941), .o(n_7942) );
in01f80 newInst_2959 ( .a(newNet_2958), .o(newNet_2959) );
na02f80 g741812 ( .a(n_38508), .b(n_38429), .o(n_38509) );
na02f80 g775531 ( .a(n_5663), .b(n_5451), .o(n_5770) );
in01f80 g777124 ( .a(n_3873), .o(n_3874) );
no02f80 g779102 ( .a(n_2038), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .o(n_2059) );
oa12f80 g784643 ( .a(n_16999), .b(n_16938), .c(n_16753), .o(n_46973) );
na02f80 g741754 ( .a(n_38491), .b(n_38490), .o(n_38492) );
in01f80 g750364 ( .a(n_29671), .o(n_29681) );
in01f80 FE_OCPC1010_n_7802 ( .a(n_7802), .o(FE_OCPN1010_n_7802) );
no02f80 FE_RC_3397_0 ( .a(FE_RN_1471_0), .b(n_16589), .o(n_46978) );
ao12f80 g742760 ( .a(n_37388), .b(n_37387), .c(n_37386), .o(n_38235) );
oa12f80 g750150 ( .a(n_29869), .b(n_30111), .c(n_29296), .o(n_30295) );
in01f80 g741293 ( .a(n_38939), .o(n_39045) );
na02f80 g741158 ( .a(FE_OCP_RBN2635_n_38806), .b(n_38061), .o(n_38864) );
no02f80 g768827 ( .a(n_11876), .b(n_11686), .o(n_12034) );
in01f80 newInst_3235 ( .a(newNet_3234), .o(newNet_3235) );
na02f80 g774182 ( .a(n_6546), .b(n_6607), .o(n_6639) );
in01f80 g762180 ( .a(n_46972), .o(n_18208) );
in01f80 newInst_357 ( .a(newNet_356), .o(newNet_357) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_5_ ( .ck(newNet_295), .d(n_1316), .o(delay_xor_ln22_unr3_stage2_stallmux_q_5_) );
no02f80 g741693 ( .a(n_38523), .b(n_38182), .o(n_38524) );
na02f80 g757777 ( .a(n_23089), .b(n_23087), .o(n_23158) );
oa12f80 g743472 ( .a(n_37635), .b(n_37634), .c(n_46240), .o(n_37730) );
in01f80 newInst_2288 ( .a(newNet_2287), .o(newNet_2288) );
in01f80 g765628 ( .a(n_14944), .o(n_14964) );
in01f80 FE_RC_3602_0 ( .a(n_45008), .o(FE_RN_1574_0) );
in01f80 g781121 ( .a(n_225), .o(n_226) );
no02f80 g762258 ( .a(n_18584), .b(n_18583), .o(n_18619) );
na02f80 g742066 ( .a(n_38007), .b(n_37948), .o(n_38033) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_11_ ( .ck(newNet_2321), .d(n_40404), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_11_) );
ao22s80 FE_RC_4200_0 ( .a(n_23923), .b(n_24327), .c(n_23924), .d(n_24348), .o(n_24451) );
na02f80 g768785 ( .a(n_11765), .b(n_11917), .o(n_11967) );
no02f80 g760361 ( .a(n_18949), .b(n_20164), .o(n_20214) );
in01f80 newInst_2968 ( .a(newNet_2967), .o(newNet_2968) );
ao22s80 FE_RC_3891_0 ( .a(n_18545), .b(n_19003), .c(n_18544), .d(n_19002), .o(n_19148) );
no02f80 g764935 ( .a(n_15612), .b(n_15536), .o(n_15613) );
in01f80 g746990 ( .a(n_34081), .o(n_34082) );
no02f80 g751766 ( .a(n_28341), .b(n_28317), .o(n_28454) );
in01f80 FE_OCP_RBC2498_n_8835 ( .a(FE_OCP_RBN2497_n_8835), .o(FE_OCP_RBN2498_n_8835) );
in01f80 g742082 ( .a(n_38237), .o(n_38238) );
no02f80 g772600 ( .a(n_8445), .b(n_8444), .o(n_8482) );
ao12f80 g744006 ( .a(n_35535), .b(n_35537), .c(n_35536), .o(n_35538) );
na02f80 g749679 ( .a(n_30057), .b(n_30025), .o(n_30026) );
na02f80 g741934 ( .a(n_38064), .b(n_38122), .o(n_38123) );
na02f80 g762732 ( .a(n_17827), .b(n_17779), .o(n_17828) );
in01f80 newInst_2149 ( .a(newNet_2148), .o(newNet_2149) );
in01f80 g743374 ( .a(n_36705), .o(n_36720) );
ao12f80 g774267 ( .a(n_6342), .b(n_44711), .c(n_6383), .o(n_6502) );
in01f80 g769911 ( .a(n_11048), .o(n_11078) );
oa22f80 g771730 ( .a(FE_OCP_RBN3543_n_44575), .b(FE_OCP_RBN2567_n_8904), .c(FE_OCP_RBN3551_n_44575), .d(n_8904), .o(n_9165) );
in01f80 FE_OCP_RBC3393_n_37557 ( .a(n_37557), .o(FE_OCP_RBN3393_n_37557) );
na02f80 g749706 ( .a(n_31228), .b(n_31227), .o(n_31229) );
no02f80 g766439 ( .a(n_14154), .b(n_14153), .o(n_14155) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_13_ ( .ck(newNet_2315), .d(n_40421), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_) );
na02f80 g746781 ( .a(n_32934), .b(n_32942), .o(n_32976) );
no03m80 FE_RC_3943_0 ( .a(FE_RN_437_0), .b(n_28039), .c(FE_OCP_RBN2165_n_28249), .o(n_28319) );
na02f80 g773622 ( .a(n_7390), .b(n_7049), .o(n_7456) );
no02f80 g763441 ( .a(n_16836), .b(n_15949), .o(n_17042) );
in01f80 g752929 ( .a(n_28053), .o(n_27901) );
in01f80 newInst_2428 ( .a(newNet_2427), .o(newNet_2428) );
no02f80 g764751 ( .a(n_46981), .b(n_15935), .o(n_16067) );
no02f80 g740215 ( .a(n_39916), .b(n_39973), .o(n_39974) );
in01f80 g741926 ( .a(n_38124), .o(n_38145) );
in01f80 g747340 ( .a(n_32575), .o(n_32576) );
no02f80 g778065 ( .a(n_3024), .b(n_3023), .o(n_3038) );
in01f80 g756900 ( .a(n_23330), .o(n_23331) );
no02f80 g745997 ( .a(n_34427), .b(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_34036) );
no02f80 g746463 ( .a(n_33330), .b(n_33143), .o(n_33382) );
no02f80 FE_RC_1305_0 ( .a(FE_RN_381_0), .b(FE_RN_382_0), .o(FE_RN_383_0) );
na02f80 g776303 ( .a(n_4388), .b(n_3029), .o(n_4521) );
na02f80 g738015 ( .a(n_42149), .b(n_42196), .o(n_42167) );
ao12f80 g764205 ( .a(n_16022), .b(n_16798), .c(n_15880), .o(n_16822) );
in01f80 g779195 ( .a(n_1965), .o(n_2302) );
in01f80 g756862 ( .a(n_23753), .o(n_23754) );
na02f80 g778123 ( .a(n_2845), .b(n_2844), .o(n_2846) );
in01f80 newInst_2398 ( .a(newNet_2271), .o(newNet_2398) );
ao12f80 g739262 ( .a(n_40932), .b(n_45155), .c(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n_40952) );
in01f80 g751531 ( .a(n_28471), .o(n_28472) );
na02f80 g757978 ( .a(n_22311), .b(n_22046), .o(n_22312) );
in01f80 g740133 ( .a(n_39866), .o(n_39902) );
in01f80 newInst_2496 ( .a(newNet_1734), .o(newNet_2496) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_20_ ( .ck(newNet_3317), .d(n_32192), .o(delay_add_ln22_unr20_stage8_stallmux_q_20_) );
in01f80 g770226 ( .a(n_10755), .o(n_10756) );
no02f80 g759931 ( .a(n_21374), .b(n_21373), .o(n_21403) );
no02f80 FE_RC_1356_0 ( .a(n_30712), .b(FE_RN_404_0), .o(n_46957) );
in01f80 g776144 ( .a(n_5077), .o(n_5114) );
in01f80 g740554 ( .a(n_39672), .o(n_39655) );
in01f80 g769947 ( .a(n_11102), .o(n_11103) );
na02f80 g739555 ( .a(n_40653), .b(n_40642), .o(n_40660) );
na02f80 g749794 ( .a(n_31338), .b(n_31569), .o(n_31625) );
oa12f80 g764718 ( .a(n_15258), .b(n_15804), .c(n_15180), .o(n_15805) );
in01f80 g780257 ( .a(n_1087), .o(n_1129) );
na02f80 g775765 ( .a(n_5305), .b(n_5125), .o(n_5426) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_2_ ( .ck(newNet_3605), .d(n_15221), .o(delay_add_ln22_unr11_stage5_stallmux_q_2_) );
na02f80 g762075 ( .a(FE_OCP_RBN2205_n_18242), .b(n_18329), .o(n_18354) );
in01f80 g775504 ( .a(n_5844), .o(n_5845) );
no02f80 g763920 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_), .o(n_17355) );
oa22f80 FE_RC_356_0 ( .a(n_15908), .b(n_15601), .c(n_15602), .d(n_15909), .o(n_16088) );
na02f80 g736926 ( .a(n_43038), .b(n_42668), .o(n_43111) );
oa12f80 g763167 ( .a(n_17172), .b(n_17287), .c(n_16839), .o(n_17344) );
in01f80 g744925 ( .a(n_35003), .o(n_35027) );
ao12f80 g773543 ( .a(n_7451), .b(n_7450), .c(n_7449), .o(n_7915) );
no02f80 g740424 ( .a(FE_OCP_RBN3029_n_39942), .b(n_39590), .o(n_40168) );
ao12f80 g763700 ( .a(n_17533), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_), .o(n_17706) );
na02f80 g768017 ( .a(FE_OCP_RBN2225_n_12729), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_), .o(n_12848) );
in01f80 g740156 ( .a(n_40218), .o(n_40219) );
no02f80 g776161 ( .a(n_4653), .b(n_3029), .o(n_4840) );
na02f80 g776804 ( .a(n_4281), .b(n_4280), .o(n_4334) );
na02f80 g762619 ( .a(n_17999), .b(n_17953), .o(n_18057) );
ao22s80 FE_RC_1394_0 ( .a(n_36481), .b(FE_OCPN3791_n_36069), .c(n_36070), .d(n_36514), .o(n_36545) );
in01f80 FE_OCP_RBC2647_n_47014 ( .a(FE_OCP_RBN3590_n_47014), .o(FE_OCP_RBN2647_n_47014) );
in01f80 g757125 ( .a(n_24188), .o(n_24350) );
no02f80 g753119 ( .a(n_27213), .b(n_27464), .o(n_27504) );
in01f80 FE_RC_856_0 ( .a(n_43071), .o(FE_RN_256_0) );
no02f80 g764622 ( .a(n_15862), .b(n_14650), .o(n_15950) );
in01f80 g774513 ( .a(n_6658), .o(n_6705) );
na02f80 g754031 ( .a(n_26369), .b(FE_OCP_DRV_N1542_n_26125), .o(n_26127) );
na02f80 g779160 ( .a(n_2487), .b(FE_OFN812_n_2405), .o(n_1933) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_30_ ( .ck(newNet_3384), .d(n_27804), .o(delay_add_ln22_unr17_stage7_stallmux_q_30_) );
in01f80 g768618 ( .a(n_12212), .o(n_12194) );
no02f80 g750616 ( .a(n_29514), .b(n_29513), .o(n_29515) );
na02f80 g774074 ( .a(n_6762), .b(n_6761), .o(n_6763) );
in01f80 g775470 ( .a(n_5469), .o(n_5523) );
na02f80 g738362 ( .a(n_41518), .b(n_41517), .o(n_41519) );
in01f80 g778761 ( .a(n_2455), .o(n_2434) );
na02f80 g742843 ( .a(n_37195), .b(n_37079), .o(n_37221) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_6_ ( .ck(newNet_1281), .d(n_791), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_) );
no03m80 FE_RC_610_0 ( .a(n_38088), .b(n_38111), .c(n_38112), .o(n_38113) );
no02f80 g759313 ( .a(n_46968), .b(n_21212), .o(n_21259) );
no02f80 g747546 ( .a(n_34074), .b(n_33603), .o(n_33672) );
na02f80 g777112 ( .a(n_3989), .b(n_3912), .o(n_4128) );
in01f80 newInst_3370 ( .a(newNet_3369), .o(newNet_3370) );
in01f80 g766749 ( .a(n_15788), .o(n_14112) );
in01f80 newInst_725 ( .a(newNet_724), .o(newNet_725) );
na02f80 g770751 ( .a(FE_OCP_RBN3654_n_10100), .b(n_10183), .o(n_10592) );
oa12f80 g775487 ( .a(n_5274), .b(n_5624), .c(n_5353), .o(n_5721) );
in01f80 newInst_1452 ( .a(newNet_1451), .o(newNet_1452) );
in01f80 g764895 ( .a(n_15561), .o(n_15588) );
no02f80 g749479 ( .a(n_30508), .b(n_30200), .o(n_30556) );
in01f80 g739818 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_12_), .o(n_40454) );
in01f80 g754207 ( .a(n_26039), .o(n_26077) );
na02f80 g760397 ( .a(n_20146), .b(n_20145), .o(n_20147) );
in01f80 newInst_1981 ( .a(newNet_1980), .o(newNet_1981) );
in01f80 fopt783149 ( .a(n_1282), .o(n_44659) );
in01f80 FE_OCP_DRV_C1540_n_35427 ( .a(FE_OCP_DRV_N1539_n_35427), .o(FE_OCP_DRV_N1540_n_35427) );
in01f80 g750526 ( .a(FE_OCP_RBN2376_n_29480), .o(n_29523) );
na02f80 g784777 ( .a(FE_OCP_RBN3666_n_10106), .b(n_10226), .o(n_47263) );
no02f80 g755403 ( .a(n_24852), .b(n_24892), .o(n_24941) );
oa12f80 g738448 ( .a(n_41416), .b(FE_OCPN953_n_41540), .c(n_41407), .o(n_41838) );
no02f80 g739322 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_25_), .o(n_40861) );
na02f80 g763782 ( .a(n_16648), .b(n_16629), .o(n_16739) );
na02f80 g771053 ( .a(n_9361), .b(n_8232), .o(n_9503) );
in01f80 newInst_2931 ( .a(newNet_2930), .o(newNet_2931) );
in01f80 newInst_589 ( .a(newNet_91), .o(newNet_589) );
no02f80 g763010 ( .a(n_17590), .b(n_17589), .o(n_17622) );
na02f80 g778425 ( .a(n_2428), .b(n_2427), .o(n_2429) );
in01f80 FE_RC_2740_0 ( .a(n_37661), .o(FE_RN_1162_0) );
na02f80 g741752 ( .a(n_38516), .b(n_38467), .o(n_38517) );
na02f80 g736760 ( .a(n_43054), .b(n_46943), .o(n_43045) );
in01f80 newInst_2351 ( .a(newNet_2350), .o(newNet_2351) );
oa22f80 g743599 ( .a(n_36412), .b(n_36257), .c(n_36413), .d(n_36256), .o(n_36460) );
in01f80 g759333 ( .a(n_21177), .o(n_21178) );
na02f80 g754008 ( .a(n_26104), .b(n_26084), .o(n_26159) );
na02f80 g757043 ( .a(n_23743), .b(n_23901), .o(n_23932) );
in01f80 newInst_2162 ( .a(newNet_2161), .o(newNet_2162) );
na02f80 g775349 ( .a(n_5807), .b(n_5660), .o(n_5880) );
na02f80 g774463 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .o(n_6938) );
na02f80 g770471 ( .a(n_10500), .b(n_10403), .o(n_10550) );
in01f80 FE_RC_78_0 ( .a(n_17741), .o(FE_RN_21_0) );
ao22s80 FE_RC_3461_0 ( .a(n_30320), .b(n_30670), .c(n_30321), .d(n_30698), .o(n_30820) );
in01f80 g755849 ( .a(n_24438), .o(n_24458) );
in01f80 FE_OFC804_n_46196 ( .a(n_46195), .o(FE_OFN804_n_46196) );
in01f80 fopt782975 ( .a(n_25507), .o(n_44441) );
ao12f80 g762177 ( .a(n_18627), .b(n_18626), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_19608) );
in01f80 newInst_798 ( .a(newNet_733), .o(newNet_798) );
no02f80 FE_RC_1342_0 ( .a(FE_RN_399_0), .b(FE_RN_400_0), .o(FE_RN_401_0) );
oa22f80 g764229 ( .a(n_16741), .b(n_15872), .c(n_16768), .d(n_15871), .o(n_16847) );
oa22f80 g755937 ( .a(n_25188), .b(n_24153), .c(n_25139), .d(n_24131), .o(n_25256) );
no02f80 g757451 ( .a(n_44066), .b(delay_xor_ln21_unr15_stage6_stallmux_q_11_), .o(n_23391) );
in01f80 newInst_2643 ( .a(newNet_2642), .o(newNet_2643) );
in01f80 g776338 ( .a(n_4667), .o(n_4668) );
in01f80 newInst_2215 ( .a(newNet_2214), .o(newNet_2215) );
in01f80 g762362 ( .a(n_18616), .o(n_18577) );
no03m80 FE_RC_2604_0 ( .a(FE_RN_1081_0), .b(n_17971), .c(n_17975), .o(n_18096) );
ao12f80 g747204 ( .a(n_33802), .b(n_33801), .c(n_33800), .o(n_34582) );
no02f80 g780417 ( .a(n_888), .b(n_887), .o(n_889) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_6_ ( .ck(newNet_2612), .d(n_21541), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_6_) );
in01f80 newInst_294 ( .a(newNet_153), .o(newNet_294) );
no02f80 g777650 ( .a(n_3423), .b(n_3397), .o(n_3398) );
no02f80 g766757 ( .a(n_13789), .b(n_13788), .o(n_13829) );
no02f80 g762399 ( .a(n_18421), .b(n_18419), .o(n_18498) );
ao12f80 g750661 ( .a(n_25738), .b(n_29262), .c(n_29327), .o(n_29328) );
na02f80 g759302 ( .a(n_22076), .b(n_45024), .o(n_21180) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_28_ ( .ck(newNet_2541), .d(n_27755), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_8_ ( .ck(newNet_288), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_8_) );
in01f80 g766397 ( .a(n_14359), .o(n_14397) );
no02f80 g746978 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n_33098) );
in01f80 g756534 ( .a(n_23962), .o(n_23963) );
na02f80 g762410 ( .a(FE_OFN750_n_45003), .b(n_18574), .o(n_18840) );
na02f80 g739840 ( .a(n_40431), .b(n_40226), .o(n_40442) );
na02f80 g747795 ( .a(n_33372), .b(n_33573), .o(n_33653) );
na02f80 g769134 ( .a(n_11586), .b(n_11651), .o(n_11739) );
in01f80 g758664 ( .a(n_22485), .o(n_22486) );
no02f80 g750803 ( .a(n_29212), .b(n_29186), .o(n_29318) );
no02f80 g769373 ( .a(n_45659), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_27_), .o(n_12077) );
na02f80 g775043 ( .a(n_6010), .b(n_5725), .o(n_6056) );
no02f80 g780845 ( .a(n_401), .b(n_416), .o(n_568) );
in01f80 newInst_3721 ( .a(newNet_3720), .o(newNet_3721) );
in01f80 g771177 ( .a(n_9704), .o(n_9705) );
in01f80 newInst_563 ( .a(newNet_562), .o(newNet_563) );
in01f80 g779790 ( .a(n_1431), .o(n_1432) );
in01f80 FE_OCP_RBC2729_n_4219 ( .a(FE_OCP_RBN2726_n_4219), .o(FE_OCP_RBN2729_n_4219) );
na02f80 g760420 ( .a(n_20079), .b(n_19973), .o(n_20098) );
in01f80 newInst_3419 ( .a(newNet_3418), .o(newNet_3419) );
oa12f80 g747167 ( .a(n_33932), .b(n_33931), .c(n_33930), .o(n_34547) );
ao12f80 g742659 ( .a(n_37196), .b(n_37380), .c(n_36963), .o(n_37432) );
in01f80 g745810 ( .a(n_34144), .o(n_34145) );
na02f80 g750299 ( .a(n_29778), .b(FE_OCP_DRV_N1570_n_29777), .o(n_29828) );
in01f80 FE_OCP_RBC1332_n_20249 ( .a(n_20249), .o(FE_OCP_RBN1332_n_20249) );
no02f80 g778253 ( .a(n_2763), .b(n_2565), .o(n_2829) );
in01f80 g780556 ( .a(n_761), .o(n_816) );
in01f80 g777204 ( .a(n_3677), .o(n_3706) );
in01f80 newInst_2230 ( .a(newNet_2229), .o(newNet_2230) );
in01f80 g764039 ( .a(n_19170), .o(n_19218) );
no02f80 FE_RC_3189_0 ( .a(FE_RN_1415_0), .b(FE_RN_1416_0), .o(FE_RN_1417_0) );
no02f80 g744392 ( .a(n_35485), .b(n_35502), .o(n_35577) );
na02f80 g751981 ( .a(n_28749), .b(n_27957), .o(n_28812) );
in01f80 g769123 ( .a(n_11731), .o(n_11682) );
na02f80 g756994 ( .a(n_23290), .b(n_23289), .o(n_23291) );
in01f80 g771725 ( .a(n_8923), .o(n_8983) );
no02f80 g763391 ( .a(n_16912), .b(FE_OCPN973_n_15900), .o(n_17036) );
in01f80 newInst_2863 ( .a(newNet_2862), .o(newNet_2863) );
ao12f80 g780639 ( .a(n_745), .b(n_906), .c(n_905), .o(n_865) );
na02f80 g771132 ( .a(n_9546), .b(FE_OCPN903_n_44581), .o(n_9624) );
in01f80 newInst_513 ( .a(newNet_280), .o(newNet_513) );
na02f80 g749116 ( .a(n_30904), .b(n_30936), .o(n_30941) );
in01f80 g762797 ( .a(n_17868), .o(n_17869) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_0_ ( .ck(newNet_3355), .d(n_30734), .o(delay_add_ln22_unr20_stage8_stallmux_q_0_) );
in01f80 g780342 ( .a(n_924), .o(n_981) );
in01f80 g775691 ( .a(n_5627), .o(n_5628) );
oa22f80 FE_RC_3917_0 ( .a(n_32277), .b(n_32133), .c(n_32132), .d(n_32278), .o(n_32384) );
in01f80 g780939 ( .a(n_285), .o(n_286) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_18_ ( .ck(newNet_2296), .d(n_40464), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_) );
na02f80 g765340 ( .a(FE_OCP_RBN3621_n_15135), .b(n_14265), .o(n_15571) );
na02f80 g767579 ( .a(n_13190), .b(n_13101), .o(n_13240) );
in01f80 FE_OCP_RBC2442_n_8402 ( .a(FE_OCP_RBN2441_n_8402), .o(FE_OCP_RBN2442_n_8402) );
no02f80 g740258 ( .a(n_40033), .b(n_40032), .o(n_40061) );
in01f80 newInst_463 ( .a(newNet_409), .o(newNet_463) );
ao22s80 FE_RC_518_0 ( .a(n_24085), .b(n_23732), .c(n_23731), .d(n_24084), .o(n_24165) );
na02f80 g758860 ( .a(n_21764), .b(n_21763), .o(n_21842) );
oa22f80 g748093 ( .a(n_31785), .b(n_31774), .c(n_31784), .d(n_31775), .o(n_31878) );
na02f80 g773950 ( .a(n_6991), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .o(n_7062) );
na02f80 g756761 ( .a(n_23425), .b(n_23412), .o(n_23502) );
na02f80 g779063 ( .a(n_2104), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_15_), .o(n_2111) );
na02f80 g740454 ( .a(n_39757), .b(n_39775), .o(n_39790) );
no02f80 g757449 ( .a(n_44066), .b(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .o(n_23461) );
in01f80 newInst_3657 ( .a(newNet_3656), .o(newNet_3657) );
na03f80 g747306 ( .a(FE_OCP_RBN2102_n_44962), .b(n_32690), .c(n_32688), .o(n_32691) );
ao12f80 g747860 ( .a(n_33173), .b(n_33172), .c(n_33171), .o(n_33227) );
in01f80 g777048 ( .a(n_3761), .o(n_3762) );
in01f80 newInst_1919 ( .a(newNet_1918), .o(newNet_1919) );
in01f80 g744607 ( .a(n_35330), .o(n_35331) );
no02f80 g745382 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35842), .o(n_35844) );
in01f80 newInst_666 ( .a(newNet_665), .o(newNet_666) );
in01f80 FE_OCP_RBC2467_n_8767 ( .a(n_8767), .o(FE_OCP_RBN2467_n_8767) );
in01f80 g752040 ( .a(n_28166), .o(n_28167) );
na02f80 g760700 ( .a(n_19689), .b(n_18112), .o(n_19770) );
na02f80 g745596 ( .a(n_34315), .b(n_34314), .o(n_34339) );
no02f80 g748625 ( .a(n_31423), .b(n_31194), .o(n_31465) );
no02f80 g760713 ( .a(n_19694), .b(n_19659), .o(n_19802) );
na02f80 g763529 ( .a(FE_OCP_RBN3079_n_16977), .b(FE_OCP_RBN2780_n_15595), .o(n_17114) );
na02f80 g741071 ( .a(n_39184), .b(FE_OCP_RBN3582_n_44944), .o(n_39233) );
oa12f80 g762225 ( .a(n_18134), .b(n_18135), .c(n_18133), .o(n_18188) );
oa12f80 g763309 ( .a(n_17025), .b(n_17125), .c(n_17226), .o(n_17472) );
na02f80 g778431 ( .a(n_2735), .b(n_2643), .o(n_2687) );
in01f80 g749776 ( .a(n_31629), .o(n_31630) );
no02f80 g758976 ( .a(n_21980), .b(n_21520), .o(n_22030) );
in01f80 g765505 ( .a(n_15826), .o(n_15778) );
ao12f80 g770976 ( .a(n_9555), .b(n_9637), .c(n_9659), .o(n_9762) );
na02f80 g740867 ( .a(n_39222), .b(n_39221), .o(n_39223) );
no02f80 g743951 ( .a(n_35625), .b(n_35648), .o(n_35649) );
no02f80 g744897 ( .a(n_35897), .b(FE_OCPN1794_n_30612), .o(n_35055) );
no02f80 g748748 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n_32507) );
na02f80 g778019 ( .a(n_3019), .b(n_3009), .o(n_3673) );
in01f80 g762641 ( .a(n_17952), .o(n_17953) );
in01f80 g739276 ( .a(n_40986), .o(n_40987) );
in01f80 FE_OCPC1444_n_45050 ( .a(FE_OCPN1443_n_45050), .o(FE_OCPN1444_n_45050) );
in01f80 g737400 ( .a(n_42778), .o(n_42779) );
no02f80 g764508 ( .a(n_16541), .b(n_16019), .o(n_16571) );
no02f80 FE_RC_2720_0 ( .a(n_8440), .b(FE_RN_1148_0), .o(n_8506) );
na02f80 g737763 ( .a(n_42656), .b(n_42607), .o(n_42677) );
oa12f80 g750958 ( .a(n_28815), .b(n_28967), .c(n_28867), .o(n_29015) );
oa12f80 g737223 ( .a(n_42522), .b(n_42902), .c(n_42526), .o(n_42970) );
in01f80 FE_OCP_RBC2411_n_13960 ( .a(n_13960), .o(FE_OCP_RBN2411_n_13960) );
in01f80 g769380 ( .a(n_11933), .o(n_11934) );
na02f80 g740534 ( .a(n_39672), .b(n_39654), .o(n_39685) );
no02f80 g741634 ( .a(FE_OCP_RBN2397_n_38586), .b(FE_OCP_RBN2370_n_38545), .o(n_38612) );
no02f80 g756897 ( .a(n_23313), .b(n_23096), .o(n_23314) );
na02f80 g769658 ( .a(n_11203), .b(n_11227), .o(n_11277) );
in01f80 FE_OCP_RBC2992_n_35539 ( .a(FE_OCP_RBN2989_n_35539), .o(FE_OCP_RBN2992_n_35539) );
in01f80 g774179 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n_6680) );
in01f80 g737672 ( .a(n_42724), .o(n_42725) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_3_ ( .ck(newNet_1905), .d(n_36792), .o(delay_sub_ln22_unr24_stage9_stallmux_q_3_) );
in01f80 g760188 ( .a(n_20400), .o(n_20401) );
ao22s80 FE_RC_620_0 ( .a(n_30219), .b(n_30453), .c(n_30218), .d(n_30454), .o(n_30541) );
no02f80 g743464 ( .a(n_37711), .b(n_46210), .o(n_37747) );
ao12f80 g752836 ( .a(n_28200), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n_28750) );
oa12f80 g775368 ( .a(n_5431), .b(n_5721), .c(n_5372), .o(n_5798) );
oa22f80 g737656 ( .a(FE_OCPN887_n_42367), .b(n_42116), .c(n_42392), .d(n_42101), .o(n_42815) );
no02f80 g747111 ( .a(n_33998), .b(n_33997), .o(n_34043) );
in01f80 g750755 ( .a(n_29232), .o(n_29263) );
in01f80 newInst_318 ( .a(newNet_317), .o(newNet_318) );
no02f80 g757987 ( .a(n_22196), .b(n_22128), .o(n_22307) );
no02f80 g765491 ( .a(n_15514), .b(n_15513), .o(n_15515) );
in01f80 FE_OCPC1007_n_13962 ( .a(FE_OCP_RBN2506_n_13896), .o(FE_OCPN1007_n_13962) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_31_ ( .ck(newNet_3599), .d(n_17834), .o(delay_add_ln22_unr11_stage5_stallmux_q_31_) );
in01f80 g745309 ( .a(n_35767), .o(n_35768) );
in01f80 FE_OCP_RBC1328_n_36489 ( .a(FE_OCP_RBN1327_n_36489), .o(FE_OCP_RBN1328_n_36489) );
in01f80 FE_RC_3772_0 ( .a(FE_RN_1655_0), .o(FE_RN_1654_0) );
ao12f80 g741888 ( .a(n_38357), .b(n_38356), .c(n_38355), .o(n_38430) );
oa12f80 g780171 ( .a(n_1078), .b(n_1077), .c(n_1159), .o(n_1142) );
in01f80 g750975 ( .a(n_28948), .o(n_28949) );
no02f80 g772968 ( .a(n_7785), .b(n_7676), .o(n_7838) );
in01f80 FE_OCP_RBC1988_delay_xor_ln23_unr6_stage3_stallmux_q ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .o(FE_OCP_RBN1988_delay_xor_ln23_unr6_stage3_stallmux_q) );
in01f80 FE_OCP_RBC2587_n_9492 ( .a(n_9492), .o(FE_OCP_RBN2587_n_9492) );
in01f80 g751381 ( .a(n_29817), .o(n_29408) );
in01f80 newInst_1699 ( .a(newNet_1698), .o(newNet_1699) );
no02f80 FE_RC_2182_0 ( .a(FE_OCPN1450_n_20443), .b(n_22066), .o(FE_RN_779_0) );
no02f80 g753139 ( .a(n_27309), .b(n_27386), .o(n_27492) );
ao12f80 g763204 ( .a(n_17335), .b(n_17231), .c(n_16857), .o(n_17481) );
na02f80 FE_RC_648_0 ( .a(FE_RN_204_0), .b(FE_RN_205_0), .o(FE_RN_206_0) );
na02f80 g767273 ( .a(n_13431), .b(n_12890), .o(n_13490) );
na02f80 g754154 ( .a(n_25986), .b(FE_OCPN1494_n_23398), .o(n_26025) );
na02f80 g743222 ( .a(n_36904), .b(n_36903), .o(n_36905) );
no02f80 g755994 ( .a(n_24288), .b(n_21975), .o(n_24289) );
oa12f80 g776261 ( .a(n_4757), .b(n_4786), .c(n_4756), .o(n_4828) );
oa22f80 g743077 ( .a(n_36461), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .d(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n_37456) );
na02f80 FE_RC_2453_0 ( .a(FE_RN_981_0), .b(n_42201), .o(FE_RN_982_0) );
no02f80 g763769 ( .a(n_17107), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17266) );
no02f80 g740498 ( .a(n_39711), .b(n_39686), .o(n_39712) );
no02f80 g755324 ( .a(n_24984), .b(n_25035), .o(n_25107) );
in01f80 g739864 ( .a(n_40417), .o(n_40418) );
in01f80 FE_OCP_RBC2735_n_14985 ( .a(n_14985), .o(FE_OCP_RBN2735_n_14985) );
no02f80 g764435 ( .a(n_16117), .b(FE_OCPN3775_n_14730), .o(n_16163) );
ao22s80 FE_RC_2556_0 ( .a(n_28083), .b(n_28145), .c(FE_RN_529_0), .d(n_28123), .o(n_28207) );
in01f80 g750321 ( .a(n_29808), .o(n_29772) );
in01f80 newInst_544 ( .a(newNet_543), .o(newNet_544) );
in01f80 g741901 ( .a(n_38244), .o(n_38407) );
in01f80 g744096 ( .a(n_35691), .o(n_35692) );
in01f80 g774154 ( .a(n_6734), .o(n_6679) );
in01f80 g779506 ( .a(n_1609), .o(n_1610) );
oa22f80 FE_RC_1390_0 ( .a(n_22295), .b(n_22444), .c(n_22296), .d(n_22475), .o(n_22596) );
na02f80 g780494 ( .a(n_1015), .b(n_1051), .o(n_1057) );
no02f80 g779562 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .o(n_1947) );
in01f80 FE_OCP_RBC2403_n_24638 ( .a(FE_OCP_RBN2402_n_24638), .o(FE_OCP_RBN2403_n_24638) );
no02f80 g772003 ( .a(n_8875), .b(n_8539), .o(n_8876) );
ao22s80 FE_RC_1368_0 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .b(n_39546), .c(n_45840), .d(n_39531), .o(n_39597) );
no02f80 g742611 ( .a(n_37463), .b(n_37448), .o(n_37527) );
in01f80 g757686 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n_22669) );
na02f80 g765935 ( .a(n_14898), .b(n_14869), .o(n_14870) );
na02f80 g750839 ( .a(n_29064), .b(n_29038), .o(n_29167) );
in01f80 g769622 ( .a(n_11411), .o(n_11396) );
oa12f80 g762754 ( .a(n_17261), .b(n_18158), .c(n_17260), .o(n_18183) );
in01f80 g776359 ( .a(n_4595), .o(n_4596) );
no02f80 g747729 ( .a(n_33421), .b(n_33393), .o(n_33794) );
no02f80 g752958 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_), .o(n_28051) );
na02f80 g766744 ( .a(n_13828), .b(n_13801), .o(n_13944) );
in01f80 g779220 ( .a(n_1880), .o(n_2494) );
in01f80 newInst_2677 ( .a(newNet_2676), .o(newNet_2677) );
na02f80 g742185 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38298), .o(n_38300) );
ao12f80 g748776 ( .a(n_32498), .b(n_32481), .c(n_32497), .o(n_32587) );
na02f80 g765522 ( .a(n_15664), .b(n_15747), .o(n_15924) );
no02f80 g751379 ( .a(n_29358), .b(n_29007), .o(n_29487) );
in01f80 g764310 ( .a(n_16431), .o(n_16458) );
no02f80 g774758 ( .a(n_6310), .b(n_6287), .o(n_6398) );
oa22f80 g764136 ( .a(n_16602), .b(n_17584), .c(n_16579), .d(n_16338), .o(n_16633) );
in01f80 FE_OCP_RBC3502_n_38592 ( .a(n_38592), .o(FE_OCP_RBN3502_n_38592) );
no02f80 FE_RC_2240_0 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .b(FE_RN_818_0), .o(FE_RN_819_0) );
na02f80 g773677 ( .a(n_7355), .b(n_7337), .o(n_7365) );
in01f80 FE_OCP_RBC3218_n_21358 ( .a(n_21358), .o(FE_OCP_RBN3218_n_21358) );
ao22s80 g752521 ( .a(n_27645), .b(n_27468), .c(n_27634), .d(n_27467), .o(n_27743) );
in01f80 g780028 ( .a(n_1259), .o(n_1264) );
in01f80 newInst_3081 ( .a(newNet_3080), .o(newNet_3081) );
in01f80 g753962 ( .a(n_26217), .o(n_26253) );
in01f80 FE_OCP_RBC2131_n_32649 ( .a(n_32649), .o(FE_OCP_RBN2131_n_32649) );
oa12f80 g745170 ( .a(n_34477), .b(n_34601), .c(n_34522), .o(n_34576) );
na02f80 g740143 ( .a(n_39781), .b(n_39844), .o(n_39924) );
oa22f80 FE_RC_3160_0 ( .a(n_17336), .b(n_17728), .c(n_16338), .d(n_17682), .o(n_17777) );
oa12f80 g780818 ( .a(n_457), .b(n_480), .c(n_479), .o(n_481) );
in01f80 FE_OCP_RBC2877_n_10354 ( .a(n_10354), .o(FE_OCP_RBN2877_n_10354) );
no02f80 g760063 ( .a(n_20292), .b(n_20314), .o(n_20412) );
in01f80 g745375 ( .a(n_35847), .o(n_35934) );
no02f80 FE_RC_2761_0 ( .a(n_8906), .b(n_8998), .o(FE_RN_1175_0) );
in01f80 g743408 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n_36994) );
na02f80 g739106 ( .a(n_41029), .b(n_40940), .o(n_41293) );
na02f80 g761029 ( .a(n_19243), .b(n_17836), .o(n_19318) );
na02f80 g784760 ( .a(n_18268), .b(n_18368), .o(n_47246) );
in01f80 g736445 ( .a(n_43790), .o(n_43791) );
in01f80 FE_OCP_RBC3460_n_7886 ( .a(n_7886), .o(FE_OCP_RBN3460_n_7886) );
in01f80 g747356 ( .a(n_33768), .o(n_32574) );
in01f80 fopt783671 ( .a(n_45323), .o(n_45322) );
in01f80 fopt784028 ( .a(n_27593), .o(n_45766) );
na02f80 g736998 ( .a(n_43230), .b(n_42954), .o(n_43297) );
ao12f80 g760599 ( .a(n_19811), .b(n_19810), .c(n_19809), .o(n_21639) );
ao12f80 g738171 ( .a(n_41788), .b(n_41995), .c(n_41761), .o(n_42031) );
in01f80 FE_OCP_RBC2226_n_7531 ( .a(n_7531), .o(FE_OCP_RBN2226_n_7531) );
na02f80 g766075 ( .a(n_14641), .b(n_13487), .o(n_14719) );
in01f80 newInst_2223 ( .a(newNet_2222), .o(newNet_2223) );
na02f80 g769178 ( .a(n_11544), .b(n_11601), .o(n_11602) );
na02f80 g745889 ( .a(n_34065), .b(n_34079), .o(n_34138) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_1_ ( .ck(newNet_457), .d(n_27671), .o(delay_xor_ln22_unr18_stage7_stallmux_q_1_) );
in01f80 g752248 ( .a(n_28030), .o(n_28031) );
in01f80 FE_OCP_RBC3313_delay_xor_ln22_unr18_stage7_stallmux_q_2_ ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_2_), .o(FE_OCP_RBN3313_delay_xor_ln22_unr18_stage7_stallmux_q_2_) );
no02f80 g750393 ( .a(n_29643), .b(n_29663), .o(n_29697) );
no02f80 g774345 ( .a(n_6865), .b(n_6940), .o(n_7316) );
na02f80 g751426 ( .a(n_28496), .b(n_28437), .o(n_28532) );
na02f80 g768464 ( .a(n_45659), .b(delay_xor_ln21_unr9_stage4_stallmux_q_22_), .o(n_12434) );
oa22f80 g779870 ( .a(n_44652), .b(n_1127), .c(n_44637), .d(n_1088), .o(n_1338) );
oa12f80 g775029 ( .a(n_5919), .b(n_6019), .c(n_5887), .o(n_6083) );
no02f80 g766603 ( .a(n_14015), .b(n_13944), .o(n_14050) );
na02f80 g736786 ( .a(n_43248), .b(n_42962), .o(n_43268) );
oa12f80 g775992 ( .a(n_4767), .b(n_4942), .c(n_4689), .o(n_5023) );
in01f80 newInst_329 ( .a(newNet_328), .o(newNet_329) );
no02f80 g752193 ( .a(n_28085), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .o(n_28112) );
no02f80 g766268 ( .a(n_14780), .b(n_14756), .o(n_14757) );
in01f80 g771565 ( .a(n_9519), .o(n_9520) );
in01f80 g769804 ( .a(n_46424), .o(n_11142) );
oa12f80 g773114 ( .a(n_8059), .b(n_8232), .c(n_8030), .o(n_8867) );
in01f80 newInst_2062 ( .a(newNet_397), .o(newNet_2062) );
no02f80 FE_RC_2468_0 ( .a(FE_RN_992_0), .b(n_14110), .o(FE_RN_993_0) );
na02f80 g762360 ( .a(FE_OCP_RBN3409_n_45120), .b(n_17883), .o(n_18580) );
na02f80 g754457 ( .a(n_26816), .b(n_26814), .o(n_26817) );
in01f80 newInst_1550 ( .a(newNet_1549), .o(newNet_1550) );
in01f80 g781390 ( .a(beta_24), .o(n_13) );
in01f80 g769945 ( .a(n_11180), .o(n_11154) );
in01f80 g756660 ( .a(n_23599), .o(n_23821) );
oa12f80 g774165 ( .a(n_6561), .b(n_6671), .c(n_6593), .o(n_6966) );
no02f80 g739137 ( .a(n_40964), .b(n_40744), .o(n_40945) );
in01f80 newInst_3014 ( .a(newNet_433), .o(newNet_3014) );
no02f80 g777768 ( .a(n_3281), .b(n_3280), .o(n_3282) );
in01f80 g769987 ( .a(n_11058), .o(n_11059) );
na02f80 FE_RC_479_0 ( .a(FE_RN_141_0), .b(FE_RN_142_0), .o(FE_RN_143_0) );
na02f80 g740413 ( .a(FE_OCP_RBN3027_n_39942), .b(n_39612), .o(n_40267) );
na02f80 g765901 ( .a(n_14851), .b(n_14815), .o(n_14852) );
na02f80 g753410 ( .a(n_27039), .b(n_27023), .o(n_27100) );
no02f80 g771610 ( .a(n_9165), .b(FE_OCP_RBN3543_n_44575), .o(n_9337) );
in01f80 g745630 ( .a(n_34310), .o(n_34311) );
na02f80 g774507 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n_6944) );
in01f80 newInst_2509 ( .a(newNet_2508), .o(newNet_2509) );
in01f80 g753061 ( .a(n_27923), .o(n_27948) );
in01f80 g760844 ( .a(n_19530), .o(n_19531) );
na02f80 g744517 ( .a(n_35366), .b(n_30633), .o(n_35405) );
no02f80 g753435 ( .a(n_26986), .b(n_26354), .o(n_27017) );
in01f80 FE_RC_178_0 ( .a(n_12295), .o(FE_RN_57_0) );
na02f80 g768304 ( .a(n_12516), .b(n_12388), .o(n_12517) );
ms00f80 cos_out_reg_10_ ( .ck(newNet_3754), .d(n_43766), .o(cos_out_10) );
no02f80 g741981 ( .a(n_38036), .b(n_38005), .o(n_38037) );
na02f80 g747613 ( .a(n_32362), .b(n_32276), .o(n_32363) );
in01f80 g736402 ( .a(n_43836), .o(n_43837) );
no02f80 g765576 ( .a(FE_OCP_RBN1222_n_45522), .b(n_15137), .o(n_15226) );
ao12f80 g777919 ( .a(n_3108), .b(n_3111), .c(n_2589), .o(n_3157) );
oa12f80 g736287 ( .a(n_288), .b(n_43857), .c(FE_OFN3_n_43918), .o(n_43889) );
in01f80 newInst_2454 ( .a(newNet_2453), .o(newNet_2454) );
in01f80 g745138 ( .a(n_35613), .o(n_34869) );
in01f80 g781002 ( .a(n_281), .o(n_284) );
na02f80 g762214 ( .a(n_18501), .b(n_18445), .o(n_18703) );
no02f80 g742419 ( .a(n_37762), .b(n_37739), .o(n_37740) );
no02f80 g779583 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_27_), .o(n_2126) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_17_ ( .ck(newNet_2664), .d(n_22540), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_) );
na02f80 g766410 ( .a(n_14156), .b(n_14132), .o(n_14273) );
no02f80 g766727 ( .a(n_13694), .b(n_12870), .o(n_13729) );
na02f80 g749656 ( .a(n_30248), .b(n_30247), .o(n_30249) );
oa12f80 g776151 ( .a(n_4930), .b(n_4929), .c(n_4951), .o(n_4992) );
in01f80 newInst_2923 ( .a(newNet_2922), .o(newNet_2923) );
in01f80 g736789 ( .a(n_43556), .o(n_43557) );
no02f80 g779581 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .o(n_1668) );
na02f80 g780705 ( .a(n_631), .b(n_630), .o(n_632) );
in01f80 g777772 ( .a(n_3368), .o(n_3369) );
na02f80 g770577 ( .a(n_10431), .b(n_10430), .o(n_10432) );
no02f80 FE_RC_1602_0 ( .a(n_27470), .b(FE_RN_449_0), .o(n_27531) );
in01f80 g754984 ( .a(n_25867), .o(n_26546) );
na02f80 g764396 ( .a(n_16127), .b(n_16164), .o(n_16333) );
in01f80 g770922 ( .a(FE_OCP_RBN2784_n_9859), .o(n_11292) );
in01f80 g773962 ( .a(n_6934), .o(n_6935) );
in01f80 g777282 ( .a(n_4361), .o(n_4362) );
na02f80 g776034 ( .a(n_5055), .b(n_4625), .o(n_5123) );
no02f80 g748520 ( .a(n_31446), .b(FE_OCP_DRV_N1606_n_31445), .o(n_31468) );
no02f80 g739328 ( .a(n_45147), .b(delay_add_ln22_unr27_stage10_stallmux_q_10_), .o(n_40738) );
in01f80 g781259 ( .a(n_144), .o(n_145) );
na02f80 g768278 ( .a(n_12550), .b(n_12563), .o(n_12574) );
in01f80 g750768 ( .a(n_29231), .o(n_29260) );
no02f80 g777378 ( .a(n_3674), .b(FE_OCPN1042_n_3673), .o(n_3692) );
no02f80 FE_RC_2855_0 ( .a(n_13280), .b(n_13281), .o(FE_RN_1230_0) );
na02f80 g758018 ( .a(n_22197), .b(n_22187), .o(n_22268) );
in01f80 g775803 ( .a(n_5300), .o(n_5335) );
no02f80 g737608 ( .a(n_42287), .b(n_42286), .o(n_42261) );
no02f80 g748150 ( .a(n_31903), .b(n_32103), .o(n_32136) );
na02f80 g753426 ( .a(n_26768), .b(n_26723), .o(n_26883) );
in01f80 g754299 ( .a(n_25928), .o(n_26113) );
in01f80 g776673 ( .a(n_3992), .o(n_4050) );
na02f80 g740835 ( .a(n_39291), .b(n_39329), .o(n_39382) );
no02f80 FE_RC_1187_0 ( .a(n_13536), .b(FE_RN_359_0), .o(n_13703) );
in01f80 g765745 ( .a(n_14942), .o(n_14959) );
oa22f80 FE_RC_3054_0 ( .a(n_36657), .b(n_36694), .c(n_36631), .d(n_36693), .o(n_36741) );
in01f80 g775192 ( .a(n_6069), .o(n_6187) );
na02f80 g755559 ( .a(n_24573), .b(n_24537), .o(n_24694) );
in01f80 FE_RC_2501_0 ( .a(n_41782), .o(FE_RN_1015_0) );
no02f80 g739372 ( .a(n_40769), .b(FE_RN_1091_0), .o(n_41240) );
in01f80 newInst_1353 ( .a(newNet_1352), .o(newNet_1353) );
in01f80 g773203 ( .a(n_7681), .o(n_7682) );
in01f80 g765677 ( .a(n_15565), .o(n_15664) );
in01f80 newInst_1506 ( .a(newNet_1505), .o(newNet_1506) );
no02f80 g771983 ( .a(FE_OCP_RBN3644_n_44490), .b(n_9587), .o(n_9649) );
na02f80 g744676 ( .a(n_35179), .b(n_35084), .o(n_35239) );
in01f80 g779835 ( .a(n_1377), .o(n_1575) );
no02f80 g776058 ( .a(n_5117), .b(n_5203), .o(n_5405) );
in01f80 g757837 ( .a(n_23009), .o(n_23010) );
in01f80 g759477 ( .a(n_20693), .o(n_20735) );
na02f80 g768292 ( .a(n_12640), .b(n_12621), .o(n_12659) );
in01f80 g739347 ( .a(n_41007), .o(n_41008) );
na02f80 g767932 ( .a(n_12707), .b(n_12706), .o(n_12708) );
in01f80 g748844 ( .a(n_31232), .o(n_31233) );
na02f80 g779321 ( .a(n_1660), .b(delay_add_ln22_unr2_stage2_stallmux_q_4_), .o(n_1724) );
in01f80 FE_OFC782_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN782_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_13_ ( .ck(newNet_1028), .d(n_17832), .o(delay_xor_ln21_unr12_stage5_stallmux_q_13_) );
in01f80 g757036 ( .a(n_23981), .o(n_24024) );
in01f80 FE_RC_2576_0 ( .a(n_2814), .o(FE_RN_1060_0) );
in01f80 g745195 ( .a(n_34707), .o(n_35703) );
na02f80 g781315 ( .a(beta_31), .b(beta_13), .o(n_116) );
no02f80 g741110 ( .a(n_38998), .b(n_38942), .o(n_38999) );
na02f80 g778946 ( .a(n_2229), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .o(n_2300) );
in01f80 FE_RC_3940_0 ( .a(n_16970), .o(FE_RN_1704_0) );
in01f80 newInst_3054 ( .a(newNet_3053), .o(newNet_3054) );
in01f80 FE_OCP_RBC3105_n_6358 ( .a(n_6358), .o(FE_OCP_RBN3105_n_6358) );
in01f80 g760793 ( .a(n_19623), .o(n_19624) );
oa22f80 g781283 ( .a(n_13), .b(n_46055), .c(n_7), .d(beta_24), .o(n_266) );
oa22f80 FE_RC_3784_0 ( .a(n_36748), .b(n_36781), .c(n_36780), .d(n_36749), .o(n_36829) );
in01f80 g777340 ( .a(n_4852), .o(n_4921) );
in01f80 g749862 ( .a(n_31526), .o(n_31527) );
na02f80 g776684 ( .a(n_4042), .b(n_3953), .o(n_4225) );
in01f80 g772303 ( .a(n_8562), .o(n_8610) );
in01f80 g743869 ( .a(n_35673), .o(n_35674) );
no02f80 g780865 ( .a(n_354), .b(beta_2), .o(n_371) );
in01f80 fopt782724 ( .a(n_44133), .o(n_44102) );
na02f80 g770622 ( .a(n_10022), .b(n_10065), .o(n_10150) );
in01f80 newInst_1592 ( .a(newNet_1591), .o(newNet_1592) );
in01f80 g774662 ( .a(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_7172) );
na02f80 g749607 ( .a(n_30375), .b(n_29982), .o(n_30374) );
in01f80 g748437 ( .a(n_31550), .o(n_31551) );
in01f80 newInst_869 ( .a(newNet_868), .o(newNet_869) );
in01f80 g779311 ( .a(n_1727), .o(n_1728) );
na02f80 FE_RC_1852_0 ( .a(n_27194), .b(n_27026), .o(n_27362) );
na02f80 g751042 ( .a(n_29974), .b(n_29997), .o(n_29998) );
na02f80 g755092 ( .a(n_25074), .b(n_25018), .o(n_25076) );
in01f80 FE_OFC814_n_18287 ( .a(FE_OFN832_n_18287), .o(FE_OFN814_n_18287) );
oa12f80 g777977 ( .a(n_2832), .b(n_3057), .c(n_2741), .o(n_3138) );
na02f80 FE_RC_3846_0 ( .a(n_23445), .b(FE_RN_1677_0), .o(FE_RN_1678_0) );
in01f80 g738121 ( .a(n_42041), .o(n_42042) );
oa12f80 g743476 ( .a(n_37678), .b(n_37713), .c(n_46241), .o(n_37725) );
na02f80 g756924 ( .a(n_24024), .b(n_23986), .o(n_24479) );
oa22f80 g768711 ( .a(n_44450), .b(n_12049), .c(n_44451), .d(n_12048), .o(n_12720) );
no02f80 g755628 ( .a(n_24614), .b(n_24613), .o(n_24636) );
na02f80 g742872 ( .a(n_37104), .b(n_37183), .o(n_37343) );
no02f80 FE_RC_3498_0 ( .a(n_31664), .b(n_31605), .o(FE_RN_1509_0) );
in01f80 g741599 ( .a(n_38652), .o(n_38630) );
no02f80 g756727 ( .a(n_23939), .b(n_23813), .o(n_24190) );
no02f80 g779804 ( .a(n_1377), .b(n_1193), .o(n_1669) );
ao12f80 g779427 ( .a(n_1668), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_12_), .o(n_1688) );
na02f80 g767338 ( .a(n_13408), .b(n_13416), .o(n_13511) );
na02f80 g781082 ( .a(n_255), .b(n_254), .o(n_256) );
no02f80 g756339 ( .a(n_23930), .b(n_23894), .o(n_23895) );
no02f80 g760194 ( .a(n_20899), .b(n_20898), .o(n_20900) );
no02f80 g758233 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_5_), .o(n_22697) );
na02f80 FE_RC_2333_0 ( .a(FE_RN_891_0), .b(n_6966), .o(n_6762) );
na02f80 g768471 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_18_), .o(n_12374) );
in01f80 newInst_823 ( .a(newNet_822), .o(newNet_823) );
in01f80 g765706 ( .a(FE_OFN766_n_15670), .o(n_16339) );
na02f80 g765003 ( .a(n_15385), .b(n_15427), .o(n_15503) );
in01f80 newInst_1594 ( .a(newNet_1593), .o(newNet_1594) );
in01f80 FE_OCP_RBC3394_n_12504 ( .a(n_12504), .o(FE_OCP_RBN3394_n_12504) );
na02f80 g746407 ( .a(n_35020), .b(n_35019), .o(n_35021) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_14_ ( .ck(newNet_1872), .d(n_16721), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_14_) );
na02f80 g742973 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_22_), .o(n_36974) );
na02f80 g780321 ( .a(n_848), .b(n_755), .o(n_849) );
no02f80 g758245 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_17_), .o(n_22844) );
oa22f80 g758523 ( .a(n_21919), .b(n_21813), .c(n_21918), .d(n_21814), .o(n_21969) );
in01f80 g759071 ( .a(n_21197), .o(n_21198) );
in01f80 FE_OCP_RBC2983_n_26767 ( .a(FE_OCP_RBN2982_n_26767), .o(FE_OCP_RBN2983_n_26767) );
no02f80 g748160 ( .a(n_31846), .b(n_30608), .o(n_31905) );
in01f80 newInst_1690 ( .a(newNet_475), .o(newNet_1690) );
na02f80 g738420 ( .a(n_41730), .b(n_41696), .o(n_41998) );
na02f80 g766800 ( .a(n_13745), .b(FE_OCP_RBN2348_n_13702), .o(n_13746) );
no02f80 g755754 ( .a(n_24445), .b(n_23999), .o(n_24463) );
na02f80 g740973 ( .a(n_39163), .b(n_38975), .o(n_39164) );
no02f80 g752728 ( .a(n_27549), .b(n_27292), .o(n_27551) );
no02f80 g753497 ( .a(n_26871), .b(n_26824), .o(n_26961) );
oa12f80 g761385 ( .a(n_18863), .b(n_18862), .c(n_18948), .o(n_18980) );
no02f80 g749118 ( .a(n_30882), .b(n_30345), .o(n_30884) );
na02f80 g773670 ( .a(n_7237), .b(n_6167), .o(n_7326) );
in01f80 g781089 ( .a(n_424), .o(n_260) );
in01f80 g745338 ( .a(n_36161), .o(n_36162) );
in01f80 g738526 ( .a(n_41622), .o(n_41623) );
in01f80 FE_OCP_RBC1137_n_11779 ( .a(n_11779), .o(FE_OCP_RBN1137_n_11779) );
ao12f80 g784657 ( .a(n_11080), .b(n_11045), .c(n_10989), .o(n_46987) );
na02f80 g737604 ( .a(n_42254), .b(n_42253), .o(n_42262) );
na02f80 g748689 ( .a(n_31204), .b(n_31203), .o(n_31205) );
na02f80 g750464 ( .a(n_29546), .b(FE_OFN788_n_25834), .o(n_29616) );
in01f80 g781366 ( .a(beta_31), .o(n_1) );
no02f80 g755591 ( .a(n_24450), .b(n_24529), .o(n_24531) );
na02f80 g736336 ( .a(n_43833), .b(n_43432), .o(n_43859) );
na02f80 g767434 ( .a(n_13338), .b(n_13360), .o(n_13401) );
ms00f80 delay_sub_ln23_0_unr18_stage7_stallmux_q_reg ( .ck(newNet_1670), .d(n_25160), .o(n_25834) );
na02f80 g742125 ( .a(n_37861), .b(n_37274), .o(n_37906) );
na02f80 g773470 ( .a(n_7522), .b(n_7521), .o(n_7559) );
in01f80 FE_RC_4036_0 ( .a(n_23486), .o(FE_RN_1753_0) );
na02f80 g753835 ( .a(n_26426), .b(n_26425), .o(n_26427) );
in01f80 g780899 ( .a(n_395), .o(n_396) );
na02f80 g738522 ( .a(FE_OCP_RBN2312_n_41420), .b(n_41542), .o(n_41583) );
no02f80 g737318 ( .a(n_42848), .b(n_42612), .o(n_42874) );
no02f80 g775174 ( .a(n_5750), .b(n_4875), .o(n_5769) );
no02f80 g747691 ( .a(n_33812), .b(n_33989), .o(n_34441) );
no02f80 g750113 ( .a(FE_OCP_RBN3566_n_29857), .b(n_29292), .o(n_30050) );
in01f80 g750432 ( .a(n_29592), .o(n_29593) );
in01f80 newInst_1673 ( .a(newNet_1672), .o(newNet_1673) );
ao12f80 g745555 ( .a(n_34402), .b(FE_OCPN1732_n_34369), .c(n_33564), .o(n_34854) );
in01f80 g767383 ( .a(n_13343), .o(n_13344) );
na02f80 g773871 ( .a(n_7044), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .o(n_7102) );
na02f80 g767371 ( .a(n_13587), .b(n_13164), .o(n_13638) );
ms00f80 mux_while_ln12_psv_q_reg_1_ ( .ck(newNet_126), .d(n_98), .o(mux_while_ln12_psv_q_1_) );
ao12f80 g746449 ( .a(n_33252), .b(n_33291), .c(n_33210), .o(n_33307) );
ao22s80 FE_RC_3530_0 ( .a(FE_RN_1526_0), .b(FE_OCP_RBN2007_n_45209), .c(n_45209), .d(n_45224), .o(n_11760) );
oa22f80 FE_RC_1645_0 ( .a(n_19033), .b(n_19518), .c(n_20307), .d(n_19475), .o(n_19666) );
na02f80 g756396 ( .a(n_23694), .b(n_23693), .o(n_23695) );
na02f80 g769825 ( .a(n_11129), .b(n_11015), .o(n_11216) );
in01f80 FE_OCP_RBC2809_n_35285 ( .a(FE_OCP_RBN2808_n_35285), .o(FE_OCP_RBN2809_n_35285) );
no02f80 g768886 ( .a(n_11835), .b(n_11834), .o(n_11836) );
no02f80 g747423 ( .a(FE_OCP_RBN2103_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_7_), .o(n_32634) );
na02f80 g778916 ( .a(n_2246), .b(delay_add_ln22_unr2_stage2_stallmux_q_20_), .o(n_2271) );
oa12f80 g770788 ( .a(n_10140), .b(n_10182), .c(n_10139), .o(n_10222) );
na02f80 g746203 ( .a(n_33622), .b(n_33157), .o(n_33648) );
in01f80 newInst_1174 ( .a(newNet_1173), .o(newNet_1174) );
na02f80 g743195 ( .a(n_36887), .b(n_36886), .o(n_36909) );
oa12f80 g742158 ( .a(n_37846), .b(n_37853), .c(n_37845), .o(n_38799) );
in01f80 newInst_2757 ( .a(newNet_2756), .o(newNet_2757) );
ao12f80 g772830 ( .a(n_8065), .b(n_8064), .c(n_8063), .o(n_9642) );
ao12f80 g743901 ( .a(n_36927), .b(n_36942), .c(n_46237), .o(n_37020) );
ao12f80 g757931 ( .a(n_23057), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n_23647) );
in01f80 newInst_2974 ( .a(newNet_2973), .o(newNet_2974) );
no02f80 g755807 ( .a(n_24274), .b(n_23926), .o(n_24272) );
no02f80 g755540 ( .a(n_24616), .b(n_24092), .o(n_24720) );
in01f80 g780300 ( .a(n_998), .o(n_1048) );
na02f80 g763940 ( .a(n_16625), .b(n_16598), .o(n_16663) );
in01f80 g751714 ( .a(n_28383), .o(n_28384) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_11_ ( .ck(newNet_3082), .d(n_1163), .o(delay_add_ln22_unr2_stage2_stallmux_q_11_) );
in01f80 g738689 ( .a(n_41826), .o(n_41827) );
no02f80 g748691 ( .a(n_31380), .b(n_29843), .o(n_31462) );
in01f80 g743998 ( .a(n_36194), .o(n_36195) );
no02f80 g759128 ( .a(n_21459), .b(FE_OCP_DRV_N1596_n_21458), .o(n_21487) );
in01f80 g745581 ( .a(n_34318), .o(n_34405) );
oa12f80 g762007 ( .a(n_18846), .b(n_18847), .c(n_18845), .o(n_18935) );
oa22f80 FE_RC_1682_0 ( .a(n_18639), .b(n_19108), .c(n_18640), .d(n_19107), .o(n_19241) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_14_ ( .ck(newNet_258), .d(n_46151), .o(delay_xor_ln22_unr6_stage3_stallmux_q_14_) );
in01f80 g769105 ( .a(n_11806), .o(n_11807) );
na02f80 g768551 ( .a(n_12276), .b(n_12309), .o(n_12508) );
oa22f80 g744813 ( .a(n_36450), .b(n_36175), .c(n_36451), .d(n_36174), .o(n_36496) );
na02f80 g746810 ( .a(n_33305), .b(n_33851), .o(n_33321) );
na02f80 g763733 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .o(n_17536) );
in01f80 newInst_3072 ( .a(newNet_3071), .o(newNet_3072) );
na02f80 g776787 ( .a(n_5629), .b(n_3938), .o(n_4024) );
na02f80 g747157 ( .a(n_32720), .b(n_32701), .o(n_32875) );
oa22f80 g776878 ( .a(n_3681), .b(n_2918), .c(n_3655), .d(n_2919), .o(n_3848) );
oa22f80 g784563 ( .a(FE_OFN800_n_46285), .b(n_10739), .c(FE_OCP_RBN3709_n_46337), .d(n_10721), .o(n_46384) );
oa22f80 g751858 ( .a(n_28161), .b(n_28146), .c(n_28162), .d(n_28192), .o(n_29391) );
no02f80 g763822 ( .a(n_17464), .b(n_17463), .o(n_17992) );
in01f80 g772794 ( .a(n_8182), .o(n_8183) );
in01f80 g742695 ( .a(n_37871), .o(n_37884) );
na02f80 g770896 ( .a(n_9762), .b(n_9740), .o(n_9908) );
ao12f80 g738666 ( .a(n_41360), .b(n_41367), .c(n_41372), .o(n_41381) );
in01f80 g772053 ( .a(n_45503), .o(n_8700) );
na02f80 g781039 ( .a(cos_out_14), .b(FE_OFN2_n_43918), .o(n_344) );
ao12f80 g747972 ( .a(n_33086), .b(n_33085), .c(n_33084), .o(n_33354) );
na02f80 g766160 ( .a(n_14462), .b(n_13469), .o(n_14550) );
no02f80 g771205 ( .a(FE_RN_1198_0), .b(n_9468), .o(n_9569) );
no02f80 g769395 ( .a(n_11403), .b(n_10292), .o(n_11418) );
no02f80 g746822 ( .a(n_33158), .b(n_33137), .o(n_33196) );
na02f80 g748835 ( .a(n_31262), .b(n_31261), .o(n_31263) );
ao12f80 g745113 ( .a(n_34464), .b(n_34749), .c(n_34460), .o(n_34855) );
ao12f80 g746561 ( .a(n_34607), .b(n_34810), .c(n_33865), .o(n_35162) );
na02f80 g753313 ( .a(n_27110), .b(n_26471), .o(n_27326) );
in01f80 g778503 ( .a(n_2520), .o(n_2458) );
no02f80 g784112 ( .a(n_45858), .b(n_6819), .o(n_45863) );
na02f80 g769892 ( .a(n_11033), .b(n_11051), .o(n_11132) );
na02f80 g779756 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .o(n_1681) );
in01f80 g751207 ( .a(n_28830), .o(n_28831) );
na02f80 g768400 ( .a(n_12491), .b(n_12439), .o(n_12500) );
no02f80 g775957 ( .a(n_4978), .b(n_4958), .o(n_5065) );
in01f80 FE_OCP_RBC2245_n_13017 ( .a(FE_OCP_RBN2243_n_13017), .o(FE_OCP_RBN2245_n_13017) );
in01f80 g746502 ( .a(n_35559), .o(n_35583) );
na02f80 g777148 ( .a(n_5001), .b(n_5069), .o(n_5113) );
no02f80 g740791 ( .a(n_39293), .b(n_39104), .o(n_39295) );
in01f80 g741668 ( .a(n_38594), .o(n_38595) );
na02f80 g779274 ( .a(n_1754), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_), .o(n_1833) );
in01f80 newInst_2900 ( .a(newNet_2899), .o(newNet_2900) );
in01f80 newInst_1850 ( .a(newNet_1849), .o(newNet_1850) );
na02f80 g750130 ( .a(FE_OCPN1786_n_30134), .b(n_30399), .o(n_30421) );
in01f80 g773046 ( .a(n_7713), .o(n_7718) );
na02f80 g738496 ( .a(n_41540), .b(n_41345), .o(n_41745) );
na02f80 g769904 ( .a(n_10978), .b(n_44498), .o(n_11051) );
in01f80 newInst_238 ( .a(newNet_37), .o(newNet_238) );
in01f80 g738354 ( .a(n_42241), .o(n_42335) );
ao12f80 g762979 ( .a(n_17684), .b(n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_7_), .o(n_17592) );
in01f80 newInst_1761 ( .a(newNet_1221), .o(newNet_1761) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_12_ ( .ck(newNet_3562), .d(n_22016), .o(delay_add_ln22_unr14_stage6_stallmux_q_12_) );
ao12f80 g739183 ( .a(n_40867), .b(n_44804), .c(n_40767), .o(n_40894) );
oa12f80 g756085 ( .a(n_23767), .b(n_24147), .c(n_23736), .o(n_24148) );
in01f80 g740928 ( .a(n_39306), .o(n_39307) );
in01f80 g769115 ( .a(n_11801), .o(n_11802) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_15_ ( .ck(newNet_3437), .d(n_27534), .o(delay_add_ln22_unr17_stage7_stallmux_q_15_) );
no02f80 g750709 ( .a(n_29197), .b(n_28736), .o(n_29273) );
in01f80 FE_OCPC1457_n_18426 ( .a(n_18426), .o(FE_OCPN1457_n_18426) );
no02f80 g740270 ( .a(n_40131), .b(FE_OCP_RBN2871_n_39542), .o(n_40099) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_11_ ( .ck(newNet_1429), .d(n_36452), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_11_) );
no02f80 g742416 ( .a(n_37742), .b(n_37741), .o(n_37757) );
oa12f80 g764659 ( .a(n_15578), .b(n_15812), .c(n_15810), .o(n_15857) );
no02f80 g758750 ( .a(n_21558), .b(n_21661), .o(n_21662) );
na02f80 g746558 ( .a(n_34912), .b(n_34760), .o(n_35019) );
no02f80 g748601 ( .a(n_31306), .b(n_31156), .o(n_31364) );
in01f80 g757369 ( .a(n_23438), .o(n_23468) );
in01f80 newInst_1281 ( .a(newNet_1280), .o(newNet_1281) );
in01f80 FE_OCPC1053_n_14098 ( .a(n_14098), .o(FE_OCPN1053_n_14098) );
no02f80 g770274 ( .a(n_10485), .b(n_10484), .o(n_10486) );
in01f80 FE_OCPC3772_n_15371 ( .a(n_15371), .o(FE_OCPN3772_n_15371) );
na03f80 g737726 ( .a(n_42343), .b(n_42417), .c(n_42416), .o(n_42440) );
na02f80 g763367 ( .a(n_16811), .b(n_16785), .o(n_16840) );
oa12f80 g744762 ( .a(n_35970), .b(n_36464), .c(n_35938), .o(n_36498) );
in01f80 newInst_2129 ( .a(newNet_2128), .o(newNet_2129) );
no02f80 g743838 ( .a(n_35714), .b(n_35576), .o(n_35878) );
in01f80 newInst_3299 ( .a(newNet_3298), .o(newNet_3299) );
in01f80 newInst_212 ( .a(newNet_211), .o(newNet_212) );
na02f80 g768073 ( .a(n_13004), .b(n_12222), .o(n_12815) );
in01f80 newInst_3508 ( .a(newNet_2761), .o(newNet_3508) );
in01f80 newInst_1370 ( .a(newNet_1369), .o(newNet_1370) );
no02f80 FE_RC_3475_0 ( .a(FE_RN_1493_0), .b(n_40050), .o(n_40124) );
oa22f80 g739779 ( .a(n_40444), .b(n_40062), .c(n_40445), .d(n_40061), .o(n_40487) );
na03f80 FE_RC_3474_0 ( .a(n_39924), .b(n_39866), .c(n_39925), .o(FE_RN_1493_0) );
no02f80 g755687 ( .a(FE_OCP_RBN2364_n_24372), .b(n_22089), .o(n_24434) );
na02f80 g762264 ( .a(n_18522), .b(n_18581), .o(n_19520) );
in01f80 g739227 ( .a(n_40906), .o(n_40907) );
no02f80 g745717 ( .a(n_34202), .b(n_44104), .o(n_34244) );
na02f80 g766865 ( .a(n_13599), .b(n_13567), .o(n_13629) );
in01f80 FE_OCP_RBC3642_n_44490 ( .a(FE_OCP_RBN3638_n_44490), .o(FE_OCP_RBN3642_n_44490) );
in01f80 newInst_3163 ( .a(newNet_2939), .o(newNet_3163) );
na02f80 g758880 ( .a(n_21399), .b(n_21287), .o(n_21477) );
in01f80 g774331 ( .a(n_6924), .o(n_6925) );
oa12f80 g773928 ( .a(n_7278), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .o(n_7292) );
ao22s80 FE_RC_207_0 ( .a(n_17409), .b(FE_OCP_RBN3211_n_44365), .c(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .d(FE_OCP_RBN3213_n_44365), .o(n_17485) );
in01f80 newInst_957 ( .a(newNet_956), .o(newNet_957) );
in01f80 FE_RC_2525_0 ( .a(n_22910), .o(FE_RN_1029_0) );
in01f80 FE_OCP_RBC2382_n_3502 ( .a(FE_OCP_RBN2381_n_3502), .o(FE_OCP_RBN2382_n_3502) );
in01f80 g753104 ( .a(n_27396), .o(n_27397) );
na02f80 g751469 ( .a(n_28843), .b(n_28887), .o(n_28914) );
in01f80 g758302 ( .a(FE_OCPN3184_n_22294), .o(n_22415) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_13_ ( .ck(newNet_263), .d(n_46175), .o(delay_xor_ln22_unr6_stage3_stallmux_q_13_) );
in01f80 newInst_3448 ( .a(newNet_3447), .o(newNet_3448) );
in01f80 newInst_1075 ( .a(newNet_738), .o(newNet_1075) );
no02f80 FE_RC_3963_0 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .b(n_23599), .o(FE_RN_1716_0) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_4_ ( .ck(newNet_1180), .d(n_4380), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_4_) );
in01f80 g751139 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_30587) );
na02f80 g751545 ( .a(n_28438), .b(n_28473), .o(n_28528) );
no02f80 g778921 ( .a(n_2246), .b(delay_add_ln22_unr2_stage2_stallmux_q_20_), .o(n_2313) );
in01f80 g754514 ( .a(n_25544), .o(n_25566) );
na02f80 g774972 ( .a(n_6180), .b(n_6117), .o(n_6207) );
in01f80 newInst_2001 ( .a(newNet_2000), .o(newNet_2001) );
ao22s80 g746866 ( .a(n_33108), .b(n_32335), .c(FE_OCP_RBN3387_n_33108), .d(delay_add_ln22_unr20_stage8_stallmux_q_31_), .o(n_33447) );
na02f80 g743730 ( .a(n_36272), .b(n_35918), .o(n_36346) );
in01f80 g769594 ( .a(n_11388), .o(n_11389) );
ao12f80 g762046 ( .a(n_18505), .b(n_18355), .c(delay_add_ln22_unr11_stage5_stallmux_q_27_), .o(n_18539) );
in01f80 g774933 ( .a(n_6266), .o(n_6259) );
in01f80 newInst_3437 ( .a(newNet_3436), .o(newNet_3437) );
in01f80 FE_OCP_RBC2766_n_4376 ( .a(n_4376), .o(FE_OCP_RBN2766_n_4376) );
no02f80 g757081 ( .a(n_23569), .b(n_23568), .o(n_23570) );
in01f80 g745044 ( .a(n_34923), .o(n_34946) );
oa22f80 FE_RC_756_0 ( .a(n_10263), .b(n_10441), .c(n_10262), .d(n_10440), .o(n_10570) );
na02f80 g757652 ( .a(n_23244), .b(n_22763), .o(n_23276) );
oa12f80 g760074 ( .a(n_21024), .b(n_21023), .c(n_21022), .o(n_21626) );
in01f80 newInst_1153 ( .a(newNet_336), .o(newNet_1153) );
na02f80 g778058 ( .a(n_2914), .b(n_2280), .o(n_2915) );
in01f80 FE_RC_2115_0 ( .a(n_24142), .o(FE_RN_733_0) );
na02f80 g779162 ( .a(n_1908), .b(FE_OFN810_n_1941), .o(n_1940) );
in01f80 newInst_2913 ( .a(newNet_2912), .o(newNet_2913) );
in01f80 g765912 ( .a(n_14916), .o(n_15139) );
in01f80 FE_RC_359_0 ( .a(n_17390), .o(FE_RN_106_0) );
no02f80 g775167 ( .a(n_5818), .b(n_4556), .o(n_5819) );
in01f80 newInst_1615 ( .a(newNet_1614), .o(newNet_1615) );
no02f80 g747216 ( .a(n_32829), .b(delay_add_ln22_unr20_stage8_stallmux_q_4_), .o(n_32846) );
na02f80 g750355 ( .a(n_29617), .b(n_29596), .o(n_29672) );
no02f80 g761321 ( .a(n_19822), .b(n_19820), .o(n_19910) );
in01f80 FE_RC_1970_0 ( .a(n_25293), .o(FE_RN_638_0) );
in01f80 g755067 ( .a(n_25378), .o(n_25379) );
na02f80 g774773 ( .a(n_6340), .b(n_6353), .o(n_6447) );
na02f80 g740606 ( .a(n_39635), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39662) );
oa12f80 g751513 ( .a(n_28528), .b(n_28460), .c(n_28473), .o(n_28865) );
ao12f80 g753826 ( .a(n_26302), .b(n_26224), .c(FE_OCPN1748_n_23354), .o(n_26340) );
no02f80 g759602 ( .a(n_20877), .b(n_20876), .o(n_20841) );
oa12f80 g773655 ( .a(n_7299), .b(n_7298), .c(n_7297), .o(n_7848) );
in01f80 FE_OCP_RBC2709_n_15135 ( .a(FE_OCP_RBN3622_n_15135), .o(FE_OCP_RBN2709_n_15135) );
na02f80 g769020 ( .a(n_11499), .b(n_11440), .o(n_11698) );
na02f80 g746785 ( .a(n_33326), .b(n_33325), .o(n_33327) );
oa12f80 g747891 ( .a(n_33126), .b(n_33125), .c(n_33124), .o(n_33626) );
na02f80 g770811 ( .a(n_10071), .b(n_9854), .o(n_10141) );
in01f80 g763891 ( .a(n_17353), .o(n_17497) );
oa12f80 g739687 ( .a(n_40376), .b(n_40524), .c(n_40112), .o(n_40536) );
na02f80 g765012 ( .a(n_15641), .b(n_15640), .o(n_15642) );
in01f80 g744101 ( .a(n_36034), .o(n_35947) );
ms00f80 delay_sub_ln23_0_unr26_stage9_stallmux_q_reg_2_ ( .ck(newNet_1445), .d(n_34666), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_) );
no02f80 g748312 ( .a(n_31763), .b(n_32168), .o(n_31802) );
no02f80 g779593 ( .a(n_1363), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1400) );
na02f80 g776831 ( .a(n_4139), .b(n_4084), .o(n_4085) );
in01f80 FE_OCP_RBC1218_n_21088 ( .a(n_21088), .o(FE_OCP_RBN1218_n_21088) );
no02f80 g768249 ( .a(n_12565), .b(delay_add_ln22_unr8_stage4_stallmux_q_17_), .o(n_12619) );
no02f80 g780875 ( .a(n_403), .b(n_399), .o(n_414) );
oa22f80 g743357 ( .a(n_36751), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .c(n_36701), .d(n_36750), .o(n_36763) );
in01f80 newInst_3614 ( .a(newNet_2372), .o(newNet_3614) );
in01f80 g737870 ( .a(n_42574), .o(n_42575) );
na02f80 g762133 ( .a(n_18243), .b(n_18220), .o(n_18259) );
ao22s80 FE_RC_3833_0 ( .a(n_30140), .b(n_30388), .c(n_30139), .d(n_30379), .o(n_30451) );
in01f80 FE_OCPC890_n_7802 ( .a(FE_OCPN889_n_7802), .o(FE_OCPN890_n_7802) );
in01f80 newInst_2889 ( .a(newNet_1948), .o(newNet_2889) );
in01f80 g751418 ( .a(n_28478), .o(n_28441) );
na02f80 g746831 ( .a(n_33077), .b(n_33055), .o(n_33343) );
ao12f80 g758737 ( .a(n_21676), .b(n_21794), .c(n_21727), .o(n_21818) );
in01f80 g743784 ( .a(n_36108), .o(n_36109) );
no02f80 g760941 ( .a(n_19449), .b(n_19350), .o(n_19625) );
in01f80 g759845 ( .a(n_22484), .o(n_24691) );
na02f80 g768752 ( .a(n_12093), .b(n_12179), .o(n_12249) );
in01f80 FE_OCP_RBC1183_n_14638 ( .a(n_14638), .o(FE_OCP_RBN1183_n_14638) );
in01f80 g749084 ( .a(n_30834), .o(n_30863) );
in01f80 newInst_2221 ( .a(newNet_2220), .o(newNet_2221) );
in01f80 g742142 ( .a(n_37939), .o(n_37940) );
na02f80 g771090 ( .a(n_9674), .b(n_9670), .o(n_9718) );
na02f80 g736800 ( .a(n_43247), .b(n_43315), .o(n_43347) );
no02f80 g748340 ( .a(n_31791), .b(n_31664), .o(n_31893) );
in01f80 g778935 ( .a(n_2297), .o(n_2298) );
na02f80 g765042 ( .a(n_15281), .b(FE_OCPN1007_n_13962), .o(n_15427) );
in01f80 g767687 ( .a(n_13132), .o(n_13133) );
in01f80 g770152 ( .a(n_10760), .o(n_10761) );
in01f80 newInst_538 ( .a(newNet_537), .o(newNet_538) );
na02f80 g753209 ( .a(n_27204), .b(n_26107), .o(n_27342) );
no02f80 g758216 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n_22877) );
na02f80 g763597 ( .a(n_17610), .b(n_17609), .o(n_18326) );
oa12f80 g736420 ( .a(n_43649), .b(n_43768), .c(n_43390), .o(n_43798) );
no02f80 g771775 ( .a(FE_OCP_RBN3547_n_44575), .b(n_9020), .o(n_9236) );
no02f80 g746981 ( .a(n_32994), .b(n_32970), .o(n_32971) );
na02f80 g748735 ( .a(n_31266), .b(n_31299), .o(n_31379) );
in01f80 g751991 ( .a(n_28858), .o(n_28859) );
in01f80 g779800 ( .a(n_1722), .o(n_1723) );
in01f80 FE_RC_3658_0 ( .a(n_21621), .o(FE_RN_1606_0) );
in01f80 newInst_2680 ( .a(newNet_2679), .o(newNet_2680) );
in01f80 g749516 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n_31887) );
in01f80 FE_OCP_RBC2780_n_15595 ( .a(FE_OCP_RBN2778_n_15595), .o(FE_OCP_RBN2780_n_15595) );
in01f80 g767289 ( .a(n_13517), .o(n_13518) );
no02f80 g756430 ( .a(n_24238), .b(n_24237), .o(n_24239) );
no02f80 g742670 ( .a(n_37380), .b(n_37188), .o(n_37403) );
in01f80 g743491 ( .a(n_36667), .o(n_36668) );
oa12f80 g736256 ( .a(n_295), .b(n_43907), .c(FE_OFN5_n_43918), .o(n_43916) );
na02f80 g777153 ( .a(n_4746), .b(n_4745), .o(n_4819) );
no02f80 g763893 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_), .o(n_17309) );
na02f80 g737062 ( .a(n_43082), .b(n_42911), .o(n_43260) );
in01f80 g738709 ( .a(n_41875), .o(n_41876) );
in01f80 g749729 ( .a(n_31147), .o(n_31228) );
in01f80 newInst_230 ( .a(tau_clk), .o(newNet_230) );
in01f80 newInst_3453 ( .a(newNet_3452), .o(newNet_3453) );
na02f80 g779269 ( .a(n_1745), .b(n_1744), .o(n_1873) );
in01f80 g743801 ( .a(n_46253), .o(n_37283) );
no02f80 g778413 ( .a(n_2684), .b(n_2683), .o(n_2751) );
ao12f80 g767508 ( .a(n_13355), .b(n_13382), .c(n_13354), .o(n_13893) );
na02f80 g742216 ( .a(n_44877), .b(n_37967), .o(n_37968) );
in01f80 g747243 ( .a(n_32668), .o(n_32669) );
no02f80 g772725 ( .a(n_8266), .b(n_7743), .o(n_8267) );
ao12f80 g771305 ( .a(n_9308), .b(n_9780), .c(n_9380), .o(n_9881) );
oa12f80 g746864 ( .a(n_32905), .b(n_32994), .c(n_32868), .o(n_33066) );
in01f80 g774803 ( .a(n_6334), .o(n_6335) );
no02f80 g773062 ( .a(n_7667), .b(n_167), .o(n_7679) );
oa22f80 g748563 ( .a(n_31335), .b(n_31331), .c(n_31334), .d(n_31330), .o(n_31405) );
na02f80 g742384 ( .a(n_37780), .b(n_37753), .o(n_37782) );
no02f80 g774934 ( .a(n_6161), .b(n_5331), .o(n_6266) );
in01f80 g754797 ( .a(n_26160), .o(n_26231) );
in01f80 g763140 ( .a(delay_xor_ln21_unr12_stage5_stallmux_q_6_), .o(n_17409) );
na02f80 g777358 ( .a(n_4759), .b(n_4777), .o(n_4999) );
in01f80 g781347 ( .a(beta_27), .o(n_47) );
in01f80 g779285 ( .a(n_2463), .o(n_2492) );
no02f80 g766686 ( .a(n_13813), .b(n_13781), .o(n_13782) );
na02f80 g742591 ( .a(n_37507), .b(n_37506), .o(n_37508) );
in01f80 g753551 ( .a(n_26785), .o(n_26758) );
na02f80 g742539 ( .a(n_37513), .b(n_37536), .o(n_37597) );
no02f80 g746692 ( .a(n_33163), .b(n_32997), .o(n_33205) );
in01f80 newInst_2554 ( .a(newNet_2553), .o(newNet_2554) );
no02f80 g779254 ( .a(n_1786), .b(n_1544), .o(n_1812) );
no02f80 g779326 ( .a(n_1660), .b(delay_add_ln22_unr2_stage2_stallmux_q_4_), .o(n_1678) );
ao12f80 g781264 ( .a(n_68), .b(n_46055), .c(beta_16), .o(n_125) );
in01f80 FE_OCP_RBC3670_n_46982 ( .a(FE_OCP_RBN3669_n_46982), .o(FE_OCP_RBN3670_n_46982) );
ao12f80 g756623 ( .a(n_23418), .b(n_23579), .c(n_23455), .o(n_23666) );
ao22s80 g779169 ( .a(n_1934), .b(n_1717), .c(n_1959), .d(n_1718), .o(n_2015) );
in01f80 g756855 ( .a(n_47245), .o(n_23460) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_0_ ( .ck(newNet_531), .d(n_22424), .o(delay_xor_ln22_unr15_stage6_stallmux_q_0_) );
in01f80 newInst_1821 ( .a(newNet_1342), .o(newNet_1821) );
no02f80 g779249 ( .a(n_1853), .b(n_1595), .o(n_1889) );
in01f80 g736909 ( .a(n_43632), .o(n_43633) );
in01f80 FE_RC_1341_0 ( .a(n_4363), .o(FE_RN_400_0) );
no02f80 g751465 ( .a(n_28785), .b(n_28828), .o(n_28849) );
ao12f80 g777015 ( .a(n_3659), .b(n_3689), .c(n_3029), .o(n_3811) );
na02f80 g741247 ( .a(FE_OCP_RBN2636_n_38806), .b(n_38517), .o(n_39010) );
in01f80 g741044 ( .a(n_39329), .o(n_39330) );
in01f80 g768268 ( .a(n_12569), .o(n_12597) );
na02f80 g779345 ( .a(n_1593), .b(n_1178), .o(n_1667) );
no02f80 g750720 ( .a(n_29319), .b(n_29342), .o(n_29440) );
oa12f80 g781122 ( .a(n_42), .b(n_222), .c(n_109), .o(n_225) );
no02f80 g740017 ( .a(n_39952), .b(FE_OCP_RBN3055_n_39913), .o(n_40020) );
na02f80 g769796 ( .a(n_11216), .b(n_11189), .o(n_11307) );
in01f80 g741336 ( .a(n_38973), .o(n_39021) );
in01f80 g746192 ( .a(FE_OCP_RBN2283_n_33846), .o(n_33895) );
ao12f80 g747287 ( .a(n_32685), .b(n_32770), .c(n_32686), .o(n_32848) );
in01f80 g754873 ( .a(n_25948), .o(n_25949) );
na02f80 g736626 ( .a(n_43193), .b(n_43192), .o(n_43194) );
in01f80 g751054 ( .a(n_30062), .o(n_30129) );
no02f80 g764674 ( .a(n_15845), .b(n_15905), .o(n_16001) );
ao22s80 g743534 ( .a(n_36472), .b(n_36139), .c(n_36444), .d(n_36140), .o(n_36515) );
na02f80 g761507 ( .a(n_18867), .b(n_18858), .o(n_18945) );
no02f80 g774114 ( .a(n_6966), .b(n_6965), .o(n_6967) );
in01f80 newInst_2687 ( .a(newNet_2686), .o(newNet_2687) );
in01f80 g777743 ( .a(n_3403), .o(n_3404) );
na02f80 g753568 ( .a(n_26756), .b(n_26520), .o(n_26778) );
no02f80 g764369 ( .a(n_16288), .b(n_16188), .o(n_16322) );
oa12f80 g768379 ( .a(n_12441), .b(n_12467), .c(n_12440), .o(n_13495) );
in01f80 g743119 ( .a(n_37102), .o(n_37043) );
in01f80 g767747 ( .a(n_13126), .o(n_13127) );
in01f80 g737649 ( .a(n_42728), .o(n_42729) );
na02f80 g770783 ( .a(FE_OCP_RBN3653_n_10100), .b(n_9155), .o(n_10253) );
na02f80 g754133 ( .a(n_26001), .b(n_25976), .o(n_26087) );
in01f80 newInst_3431 ( .a(newNet_3430), .o(newNet_3431) );
na02f80 g750468 ( .a(n_30549), .b(n_30548), .o(n_30550) );
oa12f80 g744822 ( .a(n_35969), .b(n_36463), .c(n_35940), .o(n_36476) );
na02f80 g737199 ( .a(n_42970), .b(n_42826), .o(n_42987) );
oa12f80 g757415 ( .a(n_23094), .b(n_23033), .c(FE_OCPN930_n_44083), .o(n_23326) );
no02f80 g779730 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n_1570) );
na02f80 g759279 ( .a(n_20802), .b(n_20578), .o(n_20831) );
no02f80 g740030 ( .a(n_40252), .b(FE_OCP_RBN3029_n_39942), .o(n_40332) );
no02f80 g740092 ( .a(n_40251), .b(FE_OCP_RBN2896_n_39575), .o(n_40252) );
na02f80 g781069 ( .a(cos_out_24), .b(FE_OFN1_n_43918), .o(n_291) );
in01f80 g778862 ( .a(n_2759), .o(n_2913) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_23_ ( .ck(newNet_2184), .d(n_1165), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_23_) );
na02f80 g777784 ( .a(n_3255), .b(n_3101), .o(n_3345) );
na02f80 g758322 ( .a(n_22066), .b(FE_OCPN1450_n_20443), .o(n_22154) );
no02f80 g757251 ( .a(n_23189), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n_23208) );
na02f80 g765941 ( .a(n_14754), .b(n_14724), .o(n_14755) );
in01f80 FE_RC_3977_0 ( .a(n_29566), .o(FE_RN_1723_0) );
na02f80 g749792 ( .a(n_31254), .b(n_31281), .o(n_31255) );
na02f80 g751445 ( .a(n_28484), .b(n_28549), .o(n_28609) );
na02f80 g753864 ( .a(n_26264), .b(FE_OCPN1048_n_24819), .o(n_26335) );
in01f80 newInst_700 ( .a(newNet_58), .o(newNet_700) );
ao12f80 g773657 ( .a(n_7317), .b(n_7332), .c(n_7316), .o(n_7888) );
na02f80 g748925 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32403) );
in01f80 newInst_647 ( .a(newNet_646), .o(newNet_647) );
in01f80 fopt783281 ( .a(n_11980), .o(n_44857) );
no02f80 g748003 ( .a(n_33003), .b(n_32459), .o(n_33006) );
no02f80 g755786 ( .a(n_24273), .b(n_24296), .o(n_24369) );
in01f80 g743457 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n_36540) );
no02f80 g778277 ( .a(n_2625), .b(n_2636), .o(n_2853) );
ao22s80 g780358 ( .a(n_806), .b(n_856), .c(n_855), .d(n_420), .o(n_910) );
ao12f80 g779136 ( .a(n_1920), .b(n_1921), .c(n_1919), .o(n_2702) );
in01f80 g774244 ( .a(n_6601), .o(n_6602) );
in01f80 newInst_10 ( .a(newNet_9), .o(newNet_10) );
in01f80 g753344 ( .a(n_27207), .o(n_27204) );
na02f80 FE_RC_1933_0 ( .a(FE_RN_614_0), .b(n_19210), .o(n_19246) );
na02f80 g760286 ( .a(FE_OCPN1261_n_20242), .b(n_19317), .o(n_20426) );
in01f80 g760278 ( .a(n_20404), .o(n_20387) );
in01f80 FE_OCP_RBC3846_FE_RN_1242_0 ( .a(FE_OCP_RBN3845_FE_RN_1242_0), .o(FE_OCP_RBN3846_FE_RN_1242_0) );
no02f80 g764173 ( .a(n_16583), .b(n_16561), .o(n_16598) );
in01f80 g767387 ( .a(n_13433), .o(n_13446) );
in01f80 newInst_3206 ( .a(newNet_3205), .o(newNet_3206) );
in01f80 g764213 ( .a(n_16816), .o(n_16817) );
no02f80 g753627 ( .a(n_26664), .b(n_26663), .o(n_26665) );
no02f80 g764953 ( .a(n_15319), .b(FE_OCP_RBN2507_n_13896), .o(n_15354) );
in01f80 g769281 ( .a(n_11580), .o(n_11617) );
in01f80 g756151 ( .a(n_24178), .o(n_24204) );
in01f80 g744122 ( .a(n_36065), .o(n_36066) );
in01f80 g753718 ( .a(n_26658), .o(n_26560) );
in01f80 newInst_340 ( .a(newNet_339), .o(newNet_340) );
oa12f80 g775160 ( .a(n_5991), .b(n_5994), .c(n_5990), .o(n_6042) );
na02f80 g743241 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .b(delay_add_ln22_unr23_stage9_stallmux_q_1_), .o(n_36802) );
na02f80 g754911 ( .a(n_25270), .b(n_24457), .o(n_25486) );
in01f80 g744150 ( .a(n_36139), .o(n_36140) );
in01f80 g764624 ( .a(n_16504), .o(n_16544) );
in01f80 g744591 ( .a(n_36662), .o(n_36678) );
in01f80 FE_OCP_RBC3821_n_44061 ( .a(n_44061), .o(FE_OCP_RBN3821_n_44061) );
no02f80 g748433 ( .a(FE_OCP_RBN3088_FE_OCPN1052_n_31674), .b(n_31017), .o(n_31786) );
no02f80 g769576 ( .a(n_11352), .b(FE_OCP_RBN3063_n_11325), .o(n_11410) );
ao12f80 g776003 ( .a(n_5060), .b(n_5059), .c(n_5058), .o(n_5196) );
in01f80 FE_OCPC889_n_7802 ( .a(n_7802), .o(FE_OCPN889_n_7802) );
no02f80 g781293 ( .a(beta_31), .b(beta_22), .o(n_93) );
no02f80 g768642 ( .a(n_12140), .b(n_12139), .o(n_12141) );
in01f80 FE_OCP_RBC1140_n_25816 ( .a(n_25816), .o(FE_OCP_RBN1140_n_25816) );
in01f80 g748522 ( .a(n_31497), .o(n_31498) );
no02f80 g749480 ( .a(n_30530), .b(n_30201), .o(n_30532) );
na02f80 g751635 ( .a(n_28390), .b(FE_OCPN1034_n_28420), .o(n_28660) );
in01f80 g779442 ( .a(n_1917), .o(n_1918) );
no02f80 g750336 ( .a(n_29648), .b(n_29702), .o(n_29703) );
in01f80 g751492 ( .a(n_28766), .o(n_28767) );
oa22f80 FE_RC_3213_0 ( .a(n_1169), .b(n_44659), .c(n_1158), .d(n_44623), .o(n_1322) );
ao12f80 g739263 ( .a(n_44797), .b(n_40823), .c(n_40573), .o(n_40824) );
in01f80 g738912 ( .a(n_41252), .o(n_41253) );
na02f80 g755689 ( .a(n_24369), .b(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24411) );
in01f80 g762266 ( .a(n_18818), .o(n_18695) );
no02f80 g737789 ( .a(n_42199), .b(n_42234), .o(n_42200) );
oa12f80 g741825 ( .a(n_38417), .b(n_38416), .c(n_38415), .o(n_38510) );
no02f80 g777846 ( .a(n_3262), .b(FE_OCPN1042_n_3673), .o(n_3295) );
in01f80 FE_RC_3003_0 ( .a(n_15196), .o(FE_RN_1314_0) );
na02f80 g781204 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_1_), .o(n_168) );
in01f80 FE_RC_4037_0 ( .a(FE_RN_1754_0), .o(n_26591) );
no02f80 g741557 ( .a(n_38689), .b(n_38688), .o(n_38732) );
no02f80 g744648 ( .a(n_36558), .b(n_36228), .o(n_36577) );
no02f80 g760293 ( .a(n_20154), .b(n_19945), .o(n_20194) );
no02f80 FE_RC_2936_0 ( .a(FE_RN_1279_0), .b(n_14921), .o(FE_RN_1280_0) );
na02f80 g766602 ( .a(n_13890), .b(FE_OFN747_n_13889), .o(n_13994) );
in01f80 newInst_3409 ( .a(newNet_3408), .o(newNet_3409) );
no02f80 g774511 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_28_), .o(n_6764) );
in01f80 g752536 ( .a(n_27672), .o(n_27648) );
na02f80 g745461 ( .a(n_34346), .b(n_34297), .o(n_34433) );
in01f80 g769121 ( .a(n_11745), .o(n_11746) );
no02f80 g772002 ( .a(FE_OCP_RBN3544_n_44575), .b(n_7861), .o(n_9219) );
no02f80 g758375 ( .a(n_22249), .b(n_21431), .o(n_22667) );
no02f80 g780877 ( .a(n_457), .b(n_493), .o(n_645) );
no02f80 g759416 ( .a(n_21030), .b(n_20993), .o(n_21061) );
oa12f80 g742891 ( .a(n_37144), .b(n_37204), .c(n_37030), .o(n_37237) );
in01f80 g738258 ( .a(n_41921), .o(n_41922) );
na02f80 g737031 ( .a(n_43030), .b(n_43052), .o(n_43192) );
na02f80 FE_RC_2429_0 ( .a(FE_RN_958_0), .b(FE_RN_965_0), .o(n_7332) );
in01f80 FE_RC_41_0 ( .a(n_2929), .o(FE_RN_9_0) );
na02f80 FE_RC_2885_0 ( .a(FE_RN_1248_0), .b(n_20094), .o(n_20123) );
no02f80 FE_RC_2231_0 ( .a(n_17359), .b(n_17360), .o(FE_RN_812_0) );
na02f80 g748884 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_), .o(n_32416) );
na02f80 g749254 ( .a(n_30759), .b(n_27131), .o(n_30805) );
in01f80 newInst_2135 ( .a(newNet_2134), .o(newNet_2135) );
ao12f80 g749732 ( .a(n_29906), .b(n_29905), .c(n_29904), .o(n_31445) );
no02f80 g757025 ( .a(n_23743), .b(n_23670), .o(n_23905) );
in01f80 newInst_2890 ( .a(newNet_2889), .o(newNet_2890) );
in01f80 FE_OCP_RBC2578_n_47017 ( .a(FE_OCP_RBN2577_n_47017), .o(FE_OCP_RBN2578_n_47017) );
oa12f80 g784077 ( .a(n_7285), .b(n_7284), .c(n_7283), .o(n_45820) );
in01f80 g759315 ( .a(n_21801), .o(n_21891) );
in01f80 newInst_3620 ( .a(newNet_1948), .o(newNet_3620) );
in01f80 g763176 ( .a(n_17250), .o(n_17251) );
ms00f80 sin_out_reg_13_ ( .ck(newNet_81), .d(n_43804), .o(sin_out_13) );
no02f80 g750696 ( .a(n_30338), .b(n_29886), .o(n_30419) );
no02f80 g760744 ( .a(n_19621), .b(n_19618), .o(n_19691) );
no02f80 g753218 ( .a(n_27207), .b(FE_OCP_RBN2782_n_25997), .o(n_27386) );
na02f80 g771178 ( .a(n_9572), .b(n_9538), .o(n_9704) );
in01f80 newInst_1564 ( .a(newNet_1563), .o(newNet_1564) );
no02f80 g750314 ( .a(n_30719), .b(n_30160), .o(n_30812) );
na02f80 g763256 ( .a(n_17088), .b(n_17002), .o(n_17287) );
na02f80 g766679 ( .a(n_13806), .b(n_13381), .o(n_13839) );
in01f80 g775175 ( .a(n_5870), .o(n_5827) );
no02f80 g777338 ( .a(FE_OCP_RBN2692_FE_OCPN843_n_3912), .b(n_4142), .o(n_4216) );
no02f80 g770821 ( .a(n_10215), .b(n_10214), .o(n_10342) );
in01f80 g740257 ( .a(n_40061), .o(n_40062) );
na02f80 g740538 ( .a(n_39658), .b(n_39667), .o(n_39698) );
in01f80 newInst_281 ( .a(newNet_149), .o(newNet_281) );
na02f80 g778593 ( .a(n_2326), .b(n_2325), .o(n_2574) );
in01f80 g751977 ( .a(n_28988), .o(n_28957) );
oa22f80 FE_RC_1371_0 ( .a(n_25583), .b(n_25925), .c(n_25926), .d(n_25584), .o(n_26045) );
no02f80 g773468 ( .a(n_7543), .b(n_7158), .o(n_7583) );
na02f80 g755238 ( .a(n_25095), .b(n_23890), .o(n_25145) );
in01f80 FE_RC_362_0 ( .a(n_375), .o(FE_RN_108_0) );
in01f80 g764646 ( .a(n_15817), .o(n_15816) );
ao12f80 g736403 ( .a(n_43683), .b(n_43822), .c(n_43466), .o(n_43836) );
na02f80 g764494 ( .a(n_16038), .b(n_14805), .o(n_16092) );
in01f80 g758915 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_6_), .o(n_23192) );
in01f80 newInst_2344 ( .a(newNet_1427), .o(newNet_2344) );
in01f80 g771270 ( .a(n_9424), .o(n_9468) );
na02f80 g777079 ( .a(n_3900), .b(FE_OCP_RBN2582_n_3734), .o(n_4070) );
na02f80 FE_RC_837_0 ( .a(FE_RN_249_0), .b(FE_RN_250_0), .o(FE_RN_251_0) );
oa22f80 g748354 ( .a(FE_OCPN1052_n_31674), .b(n_30527), .c(FE_OCP_RBN3090_FE_OCPN1052_n_31674), .d(n_30506), .o(n_31912) );
na02f80 g767946 ( .a(n_13075), .b(n_13115), .o(n_13255) );
in01f80 newInst_1063 ( .a(newNet_1062), .o(newNet_1063) );
in01f80 g741887 ( .a(n_38430), .o(n_38431) );
in01f80 g779759 ( .a(n_1569), .o(n_1514) );
oa12f80 g742162 ( .a(n_38295), .b(FE_OCP_RBN2241_n_44881), .c(n_38293), .o(n_38437) );
na02f80 g740213 ( .a(n_39838), .b(n_39803), .o(n_39897) );
oa12f80 g766512 ( .a(n_13883), .b(n_13930), .c(FE_OCP_RBN2246_n_13017), .o(n_14032) );
na02f80 g771461 ( .a(n_9606), .b(n_9605), .o(n_9607) );
na02f80 g760746 ( .a(n_19637), .b(n_19534), .o(n_19638) );
oa22f80 g747441 ( .a(n_32339), .b(n_32287), .c(n_44434), .d(n_28336), .o(n_32370) );
oa12f80 g749806 ( .a(n_31185), .b(n_31530), .c(n_31189), .o(n_31532) );
no02f80 g747814 ( .a(n_33372), .b(n_33371), .o(n_33462) );
ao12f80 g738181 ( .a(n_41970), .b(n_41969), .c(n_41968), .o(n_42304) );
no02f80 g764434 ( .a(n_16086), .b(n_14524), .o(n_16126) );
oa12f80 g779657 ( .a(n_1731), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_2183) );
na02f80 g758234 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_13_), .o(n_22920) );
no02f80 g782663 ( .a(n_8532), .b(n_8634), .o(n_44057) );
na02f80 g754546 ( .a(n_26383), .b(n_26346), .o(n_26384) );
in01f80 FE_RC_3797_0 ( .a(FE_RN_1256_0), .o(FE_RN_1659_0) );
in01f80 g771703 ( .a(n_9284), .o(n_9285) );
in01f80 g736338 ( .a(n_43846), .o(n_43854) );
in01f80 newInst_2210 ( .a(newNet_2209), .o(newNet_2210) );
no02f80 g774044 ( .a(n_6885), .b(n_6825), .o(n_6946) );
no03m80 g755571 ( .a(n_24560), .b(n_24566), .c(n_23942), .o(n_24600) );
no02f80 g757909 ( .a(n_22854), .b(n_22813), .o(n_22814) );
ao22s80 g736430 ( .a(n_43750), .b(n_43310), .c(n_43751), .d(n_43309), .o(n_43793) );
ao12f80 g770436 ( .a(n_10349), .b(n_10572), .c(n_10423), .o(n_10659) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_7_ ( .ck(newNet_1166), .d(n_4775), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_) );
na02f80 g774116 ( .a(n_6859), .b(n_6829), .o(n_6904) );
no02f80 g772719 ( .a(n_9304), .b(n_7802), .o(n_8132) );
no02f80 g740406 ( .a(n_39942), .b(n_39544), .o(n_40060) );
in01f80 g752754 ( .a(n_27128), .o(n_27161) );
ao12f80 g780700 ( .a(n_510), .b(n_635), .c(n_492), .o(n_647) );
ms00f80 cos_out_reg_3_ ( .ck(newNet_3688), .d(n_43693), .o(cos_out_3) );
in01f80 newInst_3737 ( .a(newNet_3736), .o(newNet_3737) );
in01f80 g775893 ( .a(n_5363), .o(n_5324) );
in01f80 newInst_3521 ( .a(newNet_3520), .o(newNet_3521) );
na02f80 g777616 ( .a(n_3505), .b(FE_OCP_RBN2487_n_3338), .o(n_3530) );
no02f80 g768084 ( .a(n_12914), .b(n_12326), .o(n_13200) );
no02f80 g762226 ( .a(n_18115), .b(n_18023), .o(n_18116) );
no02f80 g753423 ( .a(n_26967), .b(n_26966), .o(n_26989) );
ao12f80 g761858 ( .a(n_19021), .b(n_19020), .c(n_19019), .o(n_20135) );
in01f80 g765698 ( .a(FE_OFN766_n_15670), .o(n_16338) );
in01f80 newInst_1307 ( .a(newNet_1306), .o(newNet_1307) );
in01f80 newInst_1143 ( .a(newNet_1142), .o(newNet_1143) );
na02f80 g741647 ( .a(n_38557), .b(n_38576), .o(n_38616) );
ao12f80 g760769 ( .a(n_19593), .b(n_19592), .c(n_19602), .o(n_21458) );
in01f80 g745958 ( .a(n_35335), .o(n_35800) );
ao12f80 g758527 ( .a(n_21738), .b(n_21900), .c(n_21792), .o(n_21951) );
ao12f80 g737075 ( .a(n_43038), .b(n_43061), .c(n_43037), .o(n_43152) );
in01f80 newInst_2499 ( .a(newNet_1019), .o(newNet_2499) );
in01f80 newInst_2694 ( .a(newNet_2693), .o(newNet_2694) );
in01f80 FE_OFC1_n_43918 ( .a(FE_OFN0_n_43918), .o(FE_OFN1_n_43918) );
na02f80 FE_RC_146_0 ( .a(FE_RN_42_0), .b(FE_RN_43_0), .o(FE_RN_44_0) );
ms00f80 delay_xor_ln23_unr6_stage3_stallmux_q_reg ( .ck(newNet_127), .d(FE_OCP_RBN3075_FE_OFN807_n_46195), .o(delay_xor_ln23_unr6_stage3_stallmux_q) );
in01f80 newInst_1134 ( .a(newNet_948), .o(newNet_1134) );
in01f80 g760546 ( .a(n_20106), .o(n_19945) );
in01f80 g771919 ( .a(n_9034), .o(n_9062) );
in01f80 g746405 ( .a(n_34778), .o(n_34779) );
na02f80 g762259 ( .a(n_18617), .b(n_18616), .o(n_18618) );
na02f80 g749680 ( .a(n_31458), .b(n_31481), .o(n_31459) );
na02f80 g770728 ( .a(n_10179), .b(FE_OCP_RBN2856_n_10176), .o(n_10259) );
oa12f80 g744815 ( .a(n_35764), .b(n_36463), .c(n_36123), .o(n_36477) );
in01f80 newInst_1195 ( .a(newNet_1194), .o(newNet_1195) );
in01f80 g740736 ( .a(n_39553), .o(n_39552) );
no03m80 g743896 ( .a(n_37022), .b(n_36925), .c(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .o(n_37023) );
in01f80 newInst_133 ( .a(newNet_32), .o(newNet_133) );
na02f80 g756867 ( .a(n_24061), .b(n_24044), .o(n_24062) );
oa12f80 g747235 ( .a(n_32812), .b(n_32811), .c(n_32810), .o(n_33588) );
no02f80 g777929 ( .a(n_3122), .b(n_2785), .o(n_3216) );
no02f80 g772324 ( .a(n_8332), .b(n_8507), .o(n_8576) );
oa22f80 g748855 ( .a(n_32314), .b(n_31635), .c(n_32315), .d(n_31636), .o(n_32378) );
oa22f80 g738617 ( .a(n_41716), .b(n_41050), .c(n_41713), .d(n_41444), .o(n_41832) );
in01f80 g763841 ( .a(n_16646), .o(n_16669) );
in01f80 g754341 ( .a(n_25826), .o(n_25825) );
in01f80 g745792 ( .a(n_34303), .o(n_34365) );
na02f80 g779128 ( .a(n_1955), .b(delay_add_ln22_unr2_stage2_stallmux_q_12_), .o(n_2005) );
no02f80 g746205 ( .a(n_33753), .b(n_33340), .o(n_33807) );
in01f80 g749120 ( .a(n_30996), .o(n_30940) );
in01f80 newInst_190 ( .a(newNet_189), .o(newNet_190) );
oa12f80 g745771 ( .a(n_34163), .b(n_44112), .c(n_33613), .o(n_34575) );
na02f80 g753662 ( .a(n_26504), .b(n_26591), .o(n_26592) );
no02f80 g748268 ( .a(n_31835), .b(n_30646), .o(n_31863) );
na02f80 g784111 ( .a(n_6851), .b(n_6895), .o(n_45858) );
no02f80 g771531 ( .a(n_9268), .b(n_9389), .o(n_9445) );
no02f80 g741196 ( .a(FE_OCP_RBN2637_n_38806), .b(FE_OCP_RBN2351_n_38534), .o(n_38986) );
na02f80 g762039 ( .a(n_18847), .b(n_18614), .o(n_18911) );
in01f80 FE_RC_2595_0 ( .a(n_2882), .o(FE_RN_1074_0) );
ao12f80 g747883 ( .a(n_31794), .b(n_31938), .c(n_31862), .o(n_32001) );
no02f80 g771444 ( .a(n_9377), .b(n_9337), .o(n_9567) );
no03m80 g777819 ( .a(n_3229), .b(n_3213), .c(n_2654), .o(n_3454) );
in01f80 FE_OCPC1526_n_26587 ( .a(FE_OCPN1525_n_26587), .o(FE_OCPN1526_n_26587) );
in01f80 newInst_2071 ( .a(newNet_2070), .o(newNet_2071) );
no02f80 g763072 ( .a(n_17452), .b(n_17449), .o(n_17450) );
oa12f80 g780635 ( .a(n_745), .b(n_809), .c(n_808), .o(n_811) );
in01f80 g764251 ( .a(n_16490), .o(n_16491) );
in01f80 g778491 ( .a(n_2428), .o(n_2400) );
in01f80 FE_RC_3546_0 ( .a(FE_RN_1537_0), .o(n_32821) );
no02f80 g767075 ( .a(n_13591), .b(n_13590), .o(n_13637) );
in01f80 newInst_1235 ( .a(newNet_1234), .o(newNet_1235) );
in01f80 FE_OFC825_n_5067 ( .a(FE_OFN842_n_5067), .o(FE_OFN825_n_5067) );
na02f80 g739621 ( .a(n_40607), .b(n_44610), .o(n_40653) );
na02f80 g781021 ( .a(sin_out_22), .b(FE_OFN4_n_43918), .o(n_310) );
in01f80 FE_OCPC1748_n_23354 ( .a(FE_OCPN1747_n_23354), .o(FE_RN_1643_0) );
ao12f80 g761359 ( .a(n_18278), .b(n_18864), .c(n_18313), .o(n_18951) );
in01f80 newInst_1735 ( .a(newNet_1734), .o(newNet_1735) );
in01f80 FE_OCP_RBC2336_n_8269 ( .a(n_8269), .o(FE_OCP_RBN2336_n_8269) );
no02f80 g767526 ( .a(n_13382), .b(n_13354), .o(n_13355) );
oa22f80 g779869 ( .a(n_44652), .b(n_1048), .c(n_44637), .d(n_998), .o(n_1309) );
no02f80 g756993 ( .a(n_23215), .b(n_23250), .o(n_23252) );
in01f80 FE_RC_4183_0 ( .a(n_33855), .o(FE_RN_1829_0) );
in01f80 FE_OCP_RBC2528_n_3421 ( .a(FE_OCP_RBN2527_n_3421), .o(FE_OCP_RBN2528_n_3421) );
in01f80 g758226 ( .a(n_22654), .o(n_22655) );
no02f80 g746910 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_14_), .o(n_33160) );
in01f80 newInst_3629 ( .a(newNet_3628), .o(newNet_3629) );
no02f80 FE_RC_4078_0 ( .a(FE_RN_1777_0), .b(n_16876), .o(n_17001) );
no02f80 g754469 ( .a(n_26514), .b(n_26416), .o(n_26578) );
in01f80 g773285 ( .a(n_7599), .o(n_7617) );
no02f80 g769288 ( .a(n_11439), .b(FE_OCP_RBN2916_n_10644), .o(n_11478) );
in01f80 g748509 ( .a(n_31471), .o(n_31472) );
in01f80 g739569 ( .a(n_41343), .o(n_40658) );
no02f80 g779052 ( .a(n_2086), .b(delay_add_ln22_unr2_stage2_stallmux_q_15_), .o(n_2097) );
in01f80 g755218 ( .a(n_25201), .o(n_25315) );
in01f80 g757474 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n_22936) );
in01f80 g748603 ( .a(n_31401), .o(n_31402) );
in01f80 newInst_534 ( .a(newNet_533), .o(newNet_534) );
na02f80 g771277 ( .a(n_9588), .b(n_9379), .o(n_9657) );
in01f80 FE_RC_190_0 ( .a(n_13829), .o(FE_RN_64_0) );
in01f80 g744697 ( .a(n_36574), .o(n_36596) );
no02f80 g772854 ( .a(n_8001), .b(n_8021), .o(n_8022) );
na02f80 g766228 ( .a(n_14254), .b(FE_OCP_RBN2231_n_13141), .o(n_14415) );
in01f80 FE_OCP_RBC2143_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2140_FE_OCPN861_n_45450), .o(FE_OCP_RBN2143_FE_OCPN861_n_45450) );
no02f80 g756488 ( .a(n_23850), .b(n_23765), .o(n_23879) );
na02f80 g774019 ( .a(n_6974), .b(n_6973), .o(n_6975) );
na03f80 g737728 ( .a(n_42339), .b(n_42414), .c(n_42413), .o(n_42415) );
na02f80 g745376 ( .a(FE_OCP_RBN2987_n_35539), .b(n_35389), .o(n_35847) );
na02f80 g758159 ( .a(n_22149), .b(n_20979), .o(n_22197) );
in01f80 g778080 ( .a(n_4587), .o(n_3012) );
oa22f80 g779871 ( .a(n_44659), .b(n_981), .c(n_44623), .d(n_924), .o(n_1357) );
no02f80 g776832 ( .a(n_3887), .b(n_3864), .o(n_3888) );
in01f80 FE_OCPC3754_n_1451 ( .a(n_1451), .o(FE_OCPN3754_n_1451) );
oa22f80 FE_RC_3095_0 ( .a(n_23353), .b(FE_OCP_RBN3656_n_25997), .c(FE_OCPN1494_n_23398), .d(n_25997), .o(FE_RN_1367_0) );
oa12f80 g736275 ( .a(n_328), .b(n_43864), .c(FE_OFN3_n_43918), .o(n_43896) );
in01f80 g777072 ( .a(n_3941), .o(n_3975) );
in01f80 g758667 ( .a(n_22431), .o(n_22453) );
oa12f80 g761899 ( .a(n_18401), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_18544) );
na02f80 g758857 ( .a(n_21803), .b(n_21762), .o(n_21838) );
no02f80 g747228 ( .a(n_34497), .b(n_33929), .o(n_33972) );
na02f80 g766319 ( .a(n_14359), .b(n_13515), .o(n_14402) );
no02f80 g779418 ( .a(n_1587), .b(n_1603), .o(n_1624) );
in01f80 FE_OCP_RBC2746_n_47011 ( .a(n_47011), .o(FE_OCP_RBN2746_n_47011) );
in01f80 g745593 ( .a(n_34401), .o(n_34402) );
in01f80 g763941 ( .a(n_16611), .o(n_16612) );
na02f80 g779364 ( .a(n_1541), .b(n_1447), .o(n_1560) );
oa22f80 g747890 ( .a(n_32109), .b(n_32161), .c(n_32110), .d(n_32162), .o(n_32235) );
in01f80 g745690 ( .a(n_34261), .o(n_34291) );
in01f80 g757298 ( .a(n_23077), .o(n_23043) );
in01f80 g773205 ( .a(n_7913), .o(n_7763) );
oa12f80 g770964 ( .a(n_9594), .b(n_9764), .c(n_9571), .o(n_9851) );
in01f80 g737660 ( .a(n_42585), .o(n_42586) );
na02f80 g778165 ( .a(n_2860), .b(n_2673), .o(n_2888) );
in01f80 g755546 ( .a(n_24576), .o(n_24577) );
in01f80 g741532 ( .a(n_38729), .o(n_38730) );
in01f80 FE_OCP_RBC3542_n_44575 ( .a(n_44575), .o(FE_OCP_RBN3542_n_44575) );
ao12f80 g740810 ( .a(n_39242), .b(n_39291), .c(n_39303), .o(n_39352) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_19_ ( .ck(newNet_2394), .d(n_36460), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_) );
in01f80 g765313 ( .a(n_15264), .o(n_15265) );
in01f80 newInst_2728 ( .a(newNet_2727), .o(newNet_2728) );
ao12f80 g761367 ( .a(n_19787), .b(n_19607), .c(n_19928), .o(n_19989) );
na02f80 g776495 ( .a(n_4449), .b(n_4128), .o(n_4502) );
in01f80 g759800 ( .a(n_20476), .o(n_20505) );
in01f80 g775641 ( .a(n_5618), .o(n_5567) );
no02f80 g767068 ( .a(n_13624), .b(n_13639), .o(n_13668) );
in01f80 FE_OCP_RBC3571_n_44563 ( .a(n_44563), .o(FE_OCP_RBN3571_n_44563) );
no02f80 g775409 ( .a(n_5684), .b(n_5679), .o(n_5751) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_28_ ( .ck(newNet_2832), .d(n_12143), .o(delay_add_ln22_unr8_stage4_stallmux_q_28_) );
in01f80 newInst_3639 ( .a(newNet_3638), .o(newNet_3639) );
ao12f80 g748699 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32558), .c(n_32462), .o(n_32608) );
in01f80 g779617 ( .a(n_1945), .o(n_1946) );
na02f80 g764780 ( .a(n_15702), .b(n_15701), .o(n_15736) );
in01f80 FE_OCP_DRV_C1568_n_19751 ( .a(FE_OCP_DRV_N1567_n_19751), .o(FE_OCP_DRV_N1568_n_19751) );
oa12f80 g756255 ( .a(n_24669), .b(n_24668), .c(n_24667), .o(n_24767) );
na02f80 g773898 ( .a(n_7037), .b(n_7036), .o(n_7045) );
in01f80 newInst_742 ( .a(newNet_741), .o(newNet_742) );
no02f80 g754068 ( .a(n_26102), .b(n_26123), .o(n_26249) );
in01f80 g756694 ( .a(n_23572), .o(n_23678) );
no02f80 g778251 ( .a(n_2725), .b(n_2563), .o(n_2792) );
na02f80 g759921 ( .a(n_21051), .b(n_21169), .o(n_21252) );
no02f80 g778696 ( .a(n_2256), .b(n_1887), .o(n_2533) );
na02f80 g749779 ( .a(n_31284), .b(n_31571), .o(n_31317) );
in01f80 g737307 ( .a(n_42910), .o(n_42911) );
na02f80 g778280 ( .a(n_2535), .b(n_2527), .o(n_2754) );
in01f80 FE_OCPC3165_n_44267 ( .a(n_44267), .o(FE_OCPN3165_n_44267) );
no02f80 g775034 ( .a(n_5946), .b(n_4875), .o(n_5973) );
na02f80 g737129 ( .a(n_43009), .b(n_43012), .o(n_43015) );
na02f80 g768430 ( .a(n_12428), .b(delay_add_ln22_unr8_stage4_stallmux_q_11_), .o(n_12491) );
in01f80 newInst_2865 ( .a(newNet_41), .o(newNet_2865) );
ao12f80 g751291 ( .a(n_29051), .b(n_29708), .c(n_29072), .o(n_29747) );
na02f80 g765077 ( .a(n_15344), .b(n_15305), .o(n_15383) );
in01f80 FE_OCP_RBC1297_n_30451 ( .a(FE_OCP_RBN1296_n_30451), .o(FE_OCP_RBN1297_n_30451) );
no03m80 g743348 ( .a(n_37814), .b(n_37829), .c(n_36854), .o(n_37922) );
in01f80 g757170 ( .a(n_23616), .o(n_23646) );
no02f80 g771440 ( .a(n_9080), .b(n_8309), .o(n_9163) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_19_ ( .ck(newNet_1625), .d(n_27247), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_19_) );
in01f80 g776411 ( .a(n_4472), .o(n_4473) );
oa22f80 g780053 ( .a(n_1231), .b(n_1054), .c(n_1235), .d(n_1055), .o(n_1244) );
na02f80 g749533 ( .a(n_30387), .b(n_30223), .o(n_30452) );
in01f80 g738890 ( .a(n_41319), .o(n_41330) );
no02f80 g777689 ( .a(n_3331), .b(n_2641), .o(n_3371) );
in01f80 FE_OCP_RBC2802_n_15706 ( .a(FE_OCP_RBN2801_n_15706), .o(FE_OCP_RBN2802_n_15706) );
no02f80 g754943 ( .a(n_25505), .b(n_25553), .o(n_25561) );
in01f80 g777642 ( .a(n_3521), .o(n_3522) );
oa12f80 g763032 ( .a(n_16976), .b(n_17452), .c(n_17454), .o(n_17493) );
na02f80 g762175 ( .a(n_18191), .b(n_18166), .o(n_18266) );
in01f80 g750991 ( .a(n_30399), .o(n_28996) );
in01f80 g741829 ( .a(n_38389), .o(n_38451) );
in01f80 g752471 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_21_), .o(n_28541) );
no02f80 g772494 ( .a(n_8617), .b(n_8642), .o(n_8647) );
in01f80 g754295 ( .a(n_25902), .o(n_25903) );
in01f80 newInst_1741 ( .a(newNet_1451), .o(newNet_1741) );
na02f80 g776116 ( .a(n_4856), .b(n_4741), .o(n_4947) );
in01f80 FE_RC_2317_0 ( .a(n_35958), .o(FE_RN_881_0) );
in01f80 FE_OCP_RBC2880_n_21132 ( .a(n_21132), .o(FE_OCP_RBN2880_n_21132) );
no02f80 g762288 ( .a(n_18834), .b(n_18490), .o(n_19544) );
na02f80 g736468 ( .a(n_43691), .b(n_43227), .o(n_43728) );
oa12f80 g780194 ( .a(n_813), .b(n_837), .c(n_812), .o(n_854) );
in01f80 g775643 ( .a(n_5538), .o(n_5569) );
ao22s80 FE_RC_396_0 ( .a(n_14887), .b(n_14225), .c(n_14265), .d(n_14886), .o(n_14982) );
in01f80 FE_OCP_RBC2323_n_33942 ( .a(n_33942), .o(FE_OCP_RBN2323_n_33942) );
in01f80 newInst_1092 ( .a(newNet_416), .o(newNet_1092) );
in01f80 newInst_937 ( .a(newNet_635), .o(newNet_937) );
na02f80 g771348 ( .a(n_9048), .b(n_9016), .o(n_9271) );
no02f80 g763200 ( .a(n_17287), .b(n_16839), .o(n_17288) );
no02f80 g753895 ( .a(n_26361), .b(FE_OCPN1498_n_26360), .o(n_26392) );
ao12f80 g780247 ( .a(n_1098), .b(n_1046), .c(FE_OFN50_n_1045), .o(n_1089) );
in01f80 fopt783927 ( .a(n_45635), .o(n_45633) );
na02f80 g759005 ( .a(n_21571), .b(n_45080), .o(n_21604) );
na02f80 FE_RC_1712_0 ( .a(FE_RN_471_0), .b(FE_OCP_RBN2879_n_15553), .o(FE_RN_473_0) );
no02f80 g760910 ( .a(n_20118), .b(n_19993), .o(n_20057) );
no02f80 g755701 ( .a(n_24503), .b(n_24502), .o(n_24449) );
na02f80 g748573 ( .a(n_32658), .b(n_32656), .o(n_32657) );
in01f80 g755425 ( .a(n_24910), .o(n_24964) );
oa12f80 g780682 ( .a(n_513), .b(n_657), .c(n_536), .o(n_662) );
in01f80 g758687 ( .a(n_21960), .o(n_22012) );
in01f80 newInst_2767 ( .a(newNet_2766), .o(newNet_2767) );
in01f80 newInst_3213 ( .a(newNet_2845), .o(newNet_3213) );
in01f80 g769671 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_16_), .o(n_12537) );
na02f80 g758150 ( .a(n_22154), .b(FE_OCP_RBN3857_FE_RN_779_0), .o(n_22295) );
na02f80 g777019 ( .a(n_3813), .b(n_3735), .o(n_3875) );
in01f80 newInst_685 ( .a(newNet_684), .o(newNet_685) );
in01f80 g760602 ( .a(n_19857), .o(n_19858) );
in01f80 FE_OCP_RBC2102_n_44962 ( .a(FE_OCP_RBN3334_n_44962), .o(FE_OCP_RBN2102_n_44962) );
na04m80 g747100 ( .a(n_32721), .b(n_32549), .c(n_32790), .d(FE_OCPN1236_n_32791), .o(n_32792) );
in01f80 g771573 ( .a(n_9190), .o(n_9134) );
no02f80 g746168 ( .a(n_33715), .b(n_33714), .o(n_33731) );
ao22s80 FE_RC_1248_0 ( .a(n_37575), .b(FE_OCP_RBN2183_FE_RN_464_0), .c(n_37581), .d(n_37644), .o(n_37657) );
ao22s80 g779141 ( .a(n_1895), .b(n_1790), .c(n_1894), .d(n_1791), .o(n_2270) );
na02f80 g737366 ( .a(n_42861), .b(n_42846), .o(n_43211) );
in01f80 newInst_3219 ( .a(newNet_3218), .o(newNet_3219) );
no02f80 g751570 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_28_), .o(n_28828) );
in01f80 newInst_1149 ( .a(newNet_1148), .o(newNet_1149) );
no02f80 g754699 ( .a(n_26163), .b(n_26162), .o(n_26164) );
no02f80 g748975 ( .a(n_31024), .b(n_27518), .o(n_31136) );
ao22s80 FE_RC_1197_0 ( .a(n_8203), .b(n_8370), .c(n_8439), .d(n_8185), .o(n_8489) );
no02f80 g752912 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_29_), .o(n_28199) );
na02f80 g764897 ( .a(n_15614), .b(n_15645), .o(n_15792) );
no02f80 g779816 ( .a(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .o(n_1517) );
oa12f80 g759908 ( .a(n_20473), .b(n_20370), .c(FE_OCPN1261_n_20242), .o(n_20474) );
na02f80 g762850 ( .a(n_17596), .b(n_17445), .o(n_17689) );
na02f80 g766331 ( .a(n_14199), .b(n_14243), .o(n_14200) );
ao22s80 g736503 ( .a(n_43699), .b(n_43264), .c(n_43700), .d(n_43263), .o(n_43723) );
oa12f80 g764338 ( .a(n_15930), .b(n_16673), .c(n_16059), .o(n_16741) );
na04m80 g762914 ( .a(n_17561), .b(n_17458), .c(n_17593), .d(n_17560), .o(n_17680) );
in01f80 g778116 ( .a(n_3626), .o(n_2994) );
na02f80 g740755 ( .a(n_39352), .b(n_39363), .o(n_39444) );
na02f80 g743941 ( .a(n_36901), .b(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_36902) );
no02f80 g765516 ( .a(n_15565), .b(n_16246), .o(n_15563) );
no02f80 g739072 ( .a(n_41096), .b(n_40811), .o(n_41109) );
na02f80 g746048 ( .a(n_33955), .b(n_33974), .o(n_34224) );
in01f80 g763799 ( .a(n_17467), .o(n_17573) );
in01f80 g780217 ( .a(n_1093), .o(n_1094) );
oa12f80 g771243 ( .a(n_9835), .b(n_9834), .c(n_9833), .o(n_9916) );
in01f80 newInst_2271 ( .a(newNet_2270), .o(newNet_2271) );
in01f80 g775671 ( .a(n_5688), .o(n_5689) );
in01f80 newInst_3037 ( .a(newNet_3036), .o(newNet_3037) );
in01f80 g767091 ( .a(n_13513), .o(n_13532) );
in01f80 g772585 ( .a(n_8439), .o(n_8370) );
na02f80 g772021 ( .a(FE_OCPN996_n_44460), .b(n_9321), .o(n_9475) );
oa12f80 g755745 ( .a(n_25290), .b(n_25192), .c(n_25160), .o(n_25309) );
in01f80 newInst_2851 ( .a(newNet_2850), .o(newNet_2851) );
no02f80 g736777 ( .a(n_43270), .b(n_46938), .o(n_43219) );
na02f80 g765095 ( .a(n_15381), .b(n_15460), .o(n_15533) );
na02f80 g770145 ( .a(n_10599), .b(n_10329), .o(n_10672) );
ao22s80 g781000 ( .a(n_276), .b(n_154), .c(n_277), .d(n_153), .o(n_439) );
na02f80 g747220 ( .a(n_32696), .b(n_32733), .o(n_32755) );
in01f80 g738766 ( .a(n_41370), .o(n_41371) );
no02f80 g740685 ( .a(n_39473), .b(n_39501), .o(n_39554) );
in01f80 g766763 ( .a(n_13753), .o(n_13754) );
in01f80 newInst_1779 ( .a(newNet_1778), .o(newNet_1779) );
in01f80 newInst_1074 ( .a(newNet_1073), .o(newNet_1074) );
na02f80 g777190 ( .a(n_5187), .b(n_5287), .o(n_5342) );
in01f80 newInst_638 ( .a(newNet_637), .o(newNet_638) );
in01f80 FE_OCPC3775_n_14730 ( .a(FE_OCPN3774_n_14730), .o(FE_OCPN3775_n_14730) );
in01f80 g778676 ( .a(n_2331), .o(n_2350) );
oa12f80 g744220 ( .a(n_35429), .b(n_35495), .c(n_35459), .o(n_35537) );
na02f80 g743196 ( .a(n_36876), .b(n_36875), .o(n_36877) );
oa12f80 g764553 ( .a(n_16548), .b(n_16547), .c(n_16546), .o(n_16593) );
ao12f80 g761890 ( .a(n_18674), .b(n_18284), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_27_), .o(n_18707) );
no02f80 g777848 ( .a(n_3272), .b(n_3144), .o(n_3302) );
no02f80 g736492 ( .a(n_43664), .b(n_43692), .o(n_43705) );
no02f80 g738393 ( .a(n_41595), .b(n_41511), .o(n_41512) );
in01f80 g757637 ( .a(n_23746), .o(n_23294) );
in01f80 newInst_1869 ( .a(newNet_802), .o(newNet_1869) );
no02f80 g744275 ( .a(n_44174), .b(n_34967), .o(n_35739) );
na02f80 g742057 ( .a(FE_OCP_RBN2255_n_37844), .b(n_37894), .o(n_37955) );
in01f80 g770009 ( .a(n_11005), .o(n_11006) );
ao12f80 g780724 ( .a(n_615), .b(n_619), .c(n_614), .o(n_757) );
na02f80 g743004 ( .a(n_36983), .b(n_37047), .o(n_37159) );
no02f80 g767580 ( .a(n_12958), .b(n_13137), .o(n_13239) );
in01f80 g747923 ( .a(n_33372), .o(n_33571) );
in01f80 g778337 ( .a(n_2624), .o(n_2625) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_4_ ( .ck(newNet_622), .d(n_46385), .o(delay_xor_ln21_unr9_stage4_stallmux_q_4_) );
no02f80 g752341 ( .a(n_27822), .b(FE_OCP_RBN3306_n_44722), .o(n_27891) );
in01f80 g760524 ( .a(n_19922), .o(n_19923) );
in01f80 newInst_2263 ( .a(newNet_2262), .o(newNet_2263) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_19_ ( .ck(newNet_3424), .d(n_27686), .o(delay_add_ln22_unr17_stage7_stallmux_q_19_) );
in01f80 g758638 ( .a(n_22523), .o(n_22524) );
na02f80 g743975 ( .a(n_35948), .b(n_35980), .o(n_35981) );
no02f80 g754163 ( .a(n_26128), .b(n_25993), .o(n_26083) );
in01f80 g747935 ( .a(n_33315), .o(n_33372) );
in01f80 newInst_1713 ( .a(newNet_1712), .o(newNet_1713) );
in01f80 g739879 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(n_40299) );
in01f80 newInst_380 ( .a(newNet_379), .o(newNet_380) );
ao12f80 g763011 ( .a(n_17486), .b(n_17561), .c(n_17560), .o(n_17562) );
in01f80 newInst_2363 ( .a(newNet_2362), .o(newNet_2363) );
na02f80 g758622 ( .a(n_21983), .b(n_20273), .o(n_22034) );
in01f80 g742831 ( .a(n_37311), .o(n_37296) );
no02f80 g772353 ( .a(n_8613), .b(n_8588), .o(n_8589) );
in01f80 g779023 ( .a(n_2204), .o(n_2205) );
ao12f80 g752767 ( .a(n_27929), .b(n_27875), .c(n_27791), .o(n_27955) );
oa22f80 g758597 ( .a(n_21914), .b(n_21869), .c(n_21913), .d(n_21870), .o(n_21967) );
in01f80 FE_OCP_RBC2859_n_10399 ( .a(FE_OCP_RBN2857_n_10399), .o(FE_OCP_RBN2859_n_10399) );
in01f80 g738793 ( .a(n_41537), .o(n_41716) );
in01f80 g740879 ( .a(n_39220), .o(n_39237) );
no02f80 g752811 ( .a(n_27903), .b(n_27902), .o(n_28351) );
in01f80 g780102 ( .a(n_1217), .o(n_1216) );
in01f80 FE_OCP_RBC3469_n_7886 ( .a(FE_OCP_RBN3462_n_7886), .o(FE_OCP_RBN3469_n_7886) );
ao12f80 g741072 ( .a(n_38835), .b(FE_OCPN957_n_39096), .c(n_38144), .o(n_39337) );
na02f80 g745814 ( .a(n_44102), .b(n_34143), .o(n_34477) );
no02f80 g748575 ( .a(n_31515), .b(n_31361), .o(n_31547) );
na02f80 g763053 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_17556) );
in01f80 FE_OCP_RBC2808_n_35285 ( .a(n_35285), .o(FE_OCP_RBN2808_n_35285) );
oa12f80 g773889 ( .a(n_7059), .b(n_7058), .c(n_7060), .o(n_7991) );
no02f80 g754024 ( .a(n_26176), .b(FE_OCPN1494_n_23398), .o(n_26277) );
no02f80 g764919 ( .a(n_15679), .b(n_15678), .o(n_15790) );
no02f80 g744574 ( .a(n_35331), .b(n_35363), .o(n_35397) );
na02f80 g751831 ( .a(n_28208), .b(n_26972), .o(n_28286) );
na02f80 FE_RC_534_0 ( .a(FE_RN_165_0), .b(FE_RN_166_0), .o(FE_RN_167_0) );
no02f80 g742006 ( .a(n_38087), .b(n_38032), .o(n_38056) );
na02f80 g736852 ( .a(n_43514), .b(n_43458), .o(n_43545) );
na02f80 g758000 ( .a(n_22047), .b(n_22022), .o(n_22081) );
no02f80 g760405 ( .a(n_20031), .b(n_19919), .o(n_20104) );
na02f80 g742112 ( .a(n_37930), .b(n_37969), .o(n_38001) );
in01f80 g749811 ( .a(n_31567), .o(n_31568) );
na02f80 g765876 ( .a(n_14856), .b(n_14859), .o(n_14881) );
no02f80 g778043 ( .a(n_2980), .b(n_2777), .o(n_3063) );
no02f80 g743490 ( .a(n_36582), .b(n_36561), .o(n_36646) );
in01f80 FE_OFC831_n_19807 ( .a(n_19807), .o(FE_OFN831_n_19807) );
na02f80 g739027 ( .a(n_41103), .b(n_41102), .o(n_41104) );
oa12f80 g758977 ( .a(n_22010), .b(n_22009), .c(n_22008), .o(n_22055) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_2_ ( .ck(newNet_795), .d(n_1301), .o(delay_xor_ln21_unr3_stage2_stallmux_q_2_) );
no02f80 g736964 ( .a(n_43120), .b(n_43250), .o(n_43316) );
na02f80 g774503 ( .a(FE_OCPN895_n_6521), .b(n_6142), .o(n_6783) );
oa22f80 FE_RC_1152_0 ( .a(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .b(n_25933), .c(n_23354), .d(n_25934), .o(n_26097) );
na02f80 g778912 ( .a(n_2305), .b(n_1973), .o(n_2354) );
na02f80 g748154 ( .a(n_31847), .b(FE_OCP_RBN1297_n_30451), .o(n_31874) );
na02f80 g745262 ( .a(n_35766), .b(FE_OCP_RBN2993_n_35539), .o(n_35853) );
no02f80 g740361 ( .a(n_39739), .b(n_39738), .o(n_39751) );
oa12f80 g740696 ( .a(n_39335), .b(n_39386), .c(n_39211), .o(n_39477) );
na02f80 g740823 ( .a(n_39382), .b(n_39404), .o(n_39538) );
in01f80 g766005 ( .a(n_14763), .o(n_14762) );
in01f80 newInst_2018 ( .a(newNet_2017), .o(newNet_2018) );
in01f80 FE_RC_3048_0 ( .a(n_26704), .o(FE_RN_1335_0) );
na02f80 g765269 ( .a(n_15047), .b(FE_OCP_RBN2506_n_13896), .o(n_15082) );
in01f80 g767054 ( .a(n_13972), .o(n_14040) );
in01f80 FE_OCPC1733_n_16143 ( .a(n_16143), .o(FE_OCPN1733_n_16143) );
na02f80 g745097 ( .a(n_34790), .b(n_34789), .o(n_34791) );
na02f80 g752145 ( .a(n_28620), .b(n_28619), .o(n_28621) );
na02f80 g776049 ( .a(n_5115), .b(n_4496), .o(n_5176) );
no02f80 g742143 ( .a(FE_OCP_RBN2257_n_37844), .b(n_37519), .o(n_37939) );
no02f80 g756561 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_22_), .o(n_24182) );
in01f80 newInst_3384 ( .a(newNet_3383), .o(newNet_3384) );
in01f80 g760460 ( .a(n_20160), .o(n_20211) );
na02f80 g774924 ( .a(n_6201), .b(n_6189), .o(n_6270) );
na02f80 g761476 ( .a(n_19845), .b(n_19844), .o(n_19903) );
na02f80 g773551 ( .a(n_7472), .b(n_7448), .o(n_7486) );
no02f80 g752486 ( .a(n_27668), .b(n_27384), .o(n_27717) );
oa22f80 FE_RC_4112_0 ( .a(n_12705), .b(FE_OCP_RBN1151_n_13460), .c(n_12684), .d(n_13460), .o(n_13557) );
in01f80 newInst_3303 ( .a(newNet_3302), .o(newNet_3303) );
na02f80 FE_RC_3619_0 ( .a(FE_RN_1582_0), .b(n_20650), .o(FE_RN_1583_0) );
na02f80 g771767 ( .a(n_9034), .b(FE_OCP_RBN3554_n_44575), .o(n_9180) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_8_ ( .ck(newNet_2606), .d(FE_OCP_DRV_N1612_n_21706), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_) );
no02f80 g756899 ( .a(n_23237), .b(n_23108), .o(n_23238) );
no02f80 g760978 ( .a(n_19914), .b(n_19853), .o(n_20118) );
na02f80 g779256 ( .a(n_1767), .b(delay_add_ln22_unr2_stage2_stallmux_q_7_), .o(n_1845) );
oa22f80 g779850 ( .a(n_44652), .b(n_1132), .c(n_44637), .d(n_1106), .o(n_1350) );
in01f80 newInst_3481 ( .a(newNet_3480), .o(newNet_3481) );
no02f80 g742183 ( .a(n_44887), .b(n_38268), .o(n_38301) );
no02f80 g757982 ( .a(n_22164), .b(n_22078), .o(n_22165) );
in01f80 g753597 ( .a(n_26750), .o(n_26751) );
in01f80 g779176 ( .a(n_1903), .o(n_1904) );
na02f80 g756459 ( .a(n_23586), .b(n_23584), .o(n_23612) );
in01f80 g744603 ( .a(n_35317), .o(n_35318) );
in01f80 g755294 ( .a(n_25246), .o(n_25094) );
oa22f80 g743601 ( .a(n_36382), .b(n_35860), .c(n_36383), .d(n_35859), .o(n_36432) );
in01f80 g751966 ( .a(n_28940), .o(n_28922) );
in01f80 g766194 ( .a(n_14571), .o(n_14628) );
no02f80 g753581 ( .a(n_26652), .b(n_26663), .o(n_26699) );
in01f80 g751424 ( .a(n_28649), .o(n_28650) );
na02f80 g753521 ( .a(n_27450), .b(n_26793), .o(n_27537) );
in01f80 FE_OCP_RBC3832_n_19204 ( .a(FE_OCP_RBN3829_n_19204), .o(FE_OCP_RBN3832_n_19204) );
na02f80 g760704 ( .a(n_19720), .b(n_19719), .o(n_19721) );
na02f80 g757447 ( .a(n_23033), .b(FE_OCPN930_n_44083), .o(n_23094) );
no02f80 g752936 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_), .o(n_27881) );
in01f80 g770876 ( .a(n_10134), .o(n_10135) );
ao12f80 g757074 ( .a(n_23570), .b(n_23569), .c(n_23568), .o(n_24088) );
na02f80 g750858 ( .a(n_29157), .b(n_29155), .o(n_29156) );
in01f80 g774305 ( .a(n_6976), .o(n_6977) );
na02f80 g759280 ( .a(n_21757), .b(n_21756), .o(n_21758) );
in01f80 g746686 ( .a(FE_OCP_RBN2598_n_34388), .o(n_34473) );
ao12f80 g747165 ( .a(n_32850), .b(n_32849), .c(n_32848), .o(n_33714) );
in01f80 g757224 ( .a(n_23523), .o(n_23524) );
no02f80 g780485 ( .a(n_887), .b(n_900), .o(n_927) );
in01f80 g736487 ( .a(n_43719), .o(n_43720) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_12_ ( .ck(newNet_2788), .d(n_16575), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_) );
na02f80 g773859 ( .a(n_7028), .b(n_6871), .o(n_7065) );
na02f80 g754885 ( .a(n_25276), .b(n_25302), .o(n_25394) );
no02f80 g746131 ( .a(n_33757), .b(n_33756), .o(n_33829) );
in01f80 newInst_467 ( .a(newNet_466), .o(newNet_467) );
in01f80 g779283 ( .a(n_1827), .o(n_1828) );
na02f80 g756670 ( .a(n_23505), .b(n_23160), .o(n_23581) );
na02f80 g760088 ( .a(n_20340), .b(n_20343), .o(n_20375) );
no02f80 g767774 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_31_), .o(n_13082) );
in01f80 newInst_3447 ( .a(newNet_3446), .o(newNet_3447) );
in01f80 newInst_1502 ( .a(newNet_1501), .o(newNet_1502) );
in01f80 g757786 ( .a(n_22540), .o(n_22514) );
in01f80 g753876 ( .a(n_26329), .o(n_26330) );
in01f80 newInst_2679 ( .a(newNet_2678), .o(newNet_2679) );
na02f80 FE_RC_1791_0 ( .a(n_7017), .b(FE_RN_527_0), .o(n_7258) );
no02f80 g761498 ( .a(n_19613), .b(n_19575), .o(n_19576) );
na02f80 g779093 ( .a(n_2038), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_), .o(n_2081) );
in01f80 g768224 ( .a(FE_OCP_RBN3416_n_12739), .o(n_12914) );
ao22s80 FE_RC_3908_0 ( .a(n_30875), .b(FE_OCP_RBN2913_n_30949), .c(n_30949), .d(n_30876), .o(n_31056) );
na02f80 g749181 ( .a(n_30807), .b(n_30347), .o(n_30856) );
na02f80 g778394 ( .a(n_2512), .b(n_1836), .o(n_2627) );
no02f80 g762826 ( .a(n_17801), .b(n_17800), .o(n_17822) );
na02f80 g766644 ( .a(n_13918), .b(FE_OCP_RBN2243_n_13017), .o(n_13948) );
ao12f80 g753609 ( .a(n_26462), .b(n_26599), .c(n_26518), .o(n_26705) );
in01f80 newInst_2903 ( .a(newNet_2902), .o(newNet_2903) );
oa22f80 g740616 ( .a(n_39625), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .c(n_39617), .d(n_45841), .o(n_39680) );
no02f80 g762690 ( .a(n_17998), .b(n_17967), .o(n_18020) );
in01f80 g765616 ( .a(n_15021), .o(n_15048) );
oa22f80 g743076 ( .a(n_36590), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .d(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .o(n_37086) );
oa12f80 g770477 ( .a(n_10251), .b(n_10481), .c(n_10342), .o(n_10575) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_19_ ( .ck(newNet_730), .d(n_46181), .o(delay_xor_ln21_unr6_stage3_stallmux_q_19_) );
na02f80 FE_RC_3410_0 ( .a(FE_RN_1475_0), .b(FE_RN_1476_0), .o(FE_RN_1477_0) );
oa12f80 g740981 ( .a(n_38983), .b(n_39005), .c(n_38870), .o(n_39108) );
na02f80 g747727 ( .a(n_33373), .b(n_33601), .o(n_33994) );
in01f80 FE_OFC78_n_4117 ( .a(FE_OFN77_n_4117), .o(FE_OFN78_n_4117) );
oa12f80 g739916 ( .a(n_39904), .b(n_40049), .c(n_39820), .o(n_40164) );
na02f80 g773134 ( .a(n_7802), .b(n_8030), .o(n_8059) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_6_ ( .ck(newNet_776), .d(n_1287), .o(delay_xor_ln21_unr3_stage2_stallmux_q_6_) );
na02f80 g767520 ( .a(n_12981), .b(FE_OCP_RBN3415_n_12739), .o(n_13057) );
na02f80 g768645 ( .a(n_12100), .b(delay_add_ln22_unr8_stage4_stallmux_q_6_), .o(n_12191) );
no02f80 g744680 ( .a(n_35229), .b(n_44713), .o(n_35271) );
na02f80 g776914 ( .a(n_3853), .b(n_3760), .o(n_3932) );
ao12f80 g756952 ( .a(n_23644), .b(n_23643), .c(n_23642), .o(n_24028) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_18_ ( .ck(newNet_2959), .d(n_6233), .o(delay_add_ln22_unr5_stage3_stallmux_q_18_) );
in01f80 g763865 ( .a(n_16643), .o(n_16665) );
no02f80 g762780 ( .a(FE_OCP_RBN2140_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_10_), .o(n_17825) );
oa12f80 g780302 ( .a(n_1113), .b(n_941), .c(FE_OFN50_n_1045), .o(n_1007) );
ms00f80 delay_sub_ln23_0_unr23_stage8_stallmux_q_reg ( .ck(newNet_1552), .d(n_31530), .o(delay_sub_ln23_0_unr23_stage8_stallmux_q) );
in01f80 FE_OCP_RBC3843_n_24972 ( .a(n_24972), .o(FE_OCP_RBN3843_n_24972) );
no02f80 g739325 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_26_), .o(n_40843) );
in01f80 newInst_1926 ( .a(newNet_1925), .o(newNet_1926) );
in01f80 g771291 ( .a(n_9659), .o(n_9568) );
ao12f80 g758134 ( .a(n_22692), .b(FE_OCP_RBN2050_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n_23356) );
in01f80 FE_OCP_RBC2567_n_8904 ( .a(n_8904), .o(FE_OCP_RBN2567_n_8904) );
na02f80 g759998 ( .a(n_20660), .b(FE_OCP_RBN3521_n_19663), .o(n_20709) );
no02f80 g772878 ( .a(n_7974), .b(n_7973), .o(n_8006) );
oa12f80 g748613 ( .a(n_31271), .b(n_31308), .c(n_31268), .o(n_31334) );
in01f80 FE_RC_3895_0 ( .a(n_24645), .o(FE_RN_1691_0) );
no02f80 g778530 ( .a(n_2516), .b(n_2108), .o(n_2556) );
na02f80 g769264 ( .a(n_11627), .b(n_11007), .o(n_11651) );
na02f80 g761926 ( .a(n_18268), .b(n_17772), .o(n_18512) );
no02f80 g756902 ( .a(n_23325), .b(n_23371), .o(n_23498) );
na02f80 g745314 ( .a(n_35961), .b(n_35929), .o(n_35992) );
no02f80 g746808 ( .a(n_33253), .b(n_33231), .o(n_33267) );
no02f80 g753644 ( .a(n_26627), .b(n_26626), .o(n_26654) );
oa22f80 g784522 ( .a(n_12217), .b(FE_OFN802_n_46285), .c(n_12190), .d(FE_OFN771_n_46337), .o(n_46344) );
in01f80 g753333 ( .a(n_27086), .o(n_27087) );
na02f80 g761038 ( .a(n_19207), .b(n_19182), .o(n_19249) );
na02f80 g771744 ( .a(n_8790), .b(n_8189), .o(n_8795) );
in01f80 g750354 ( .a(n_29672), .o(n_29673) );
na02f80 g743586 ( .a(n_36458), .b(n_36032), .o(n_36488) );
no02f80 g757180 ( .a(n_23535), .b(n_22850), .o(n_23536) );
ao12f80 g774203 ( .a(n_6964), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_13_), .o(n_7064) );
in01f80 newInst_2394 ( .a(newNet_2393), .o(newNet_2394) );
na02f80 g778654 ( .a(FE_OCP_RBN2318_n_2367), .b(n_2413), .o(n_2450) );
na02f80 g749050 ( .a(n_30994), .b(n_30964), .o(n_31073) );
na02f80 g736827 ( .a(n_43127), .b(n_42906), .o(n_43140) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_6_ ( .ck(newNet_2050), .d(n_5244), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_) );
no02f80 FE_RC_2188_0 ( .a(n_21659), .b(n_21707), .o(FE_RN_783_0) );
no02f80 g750544 ( .a(n_29399), .b(n_47251), .o(n_29428) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_29_ ( .ck(newNet_3606), .d(n_17835), .o(delay_add_ln22_unr11_stage5_stallmux_q_29_) );
no02f80 g747173 ( .a(n_32830), .b(n_32651), .o(n_32869) );
in01f80 g781272 ( .a(n_153), .o(n_154) );
in01f80 newInst_1317 ( .a(newNet_943), .o(newNet_1317) );
na02f80 g778022 ( .a(n_2996), .b(n_2248), .o(n_3019) );
na02f80 FE_RC_2451_0 ( .a(FE_RN_980_0), .b(n_13587), .o(n_13636) );
na02f80 g771004 ( .a(n_10045), .b(n_10002), .o(n_10003) );
no02f80 g751952 ( .a(n_28793), .b(n_28901), .o(n_28924) );
na02f80 g741721 ( .a(n_38457), .b(n_38349), .o(n_38477) );
na02f80 g745245 ( .a(n_36681), .b(FE_OCP_RBN2994_n_35539), .o(n_36086) );
na02f80 g748627 ( .a(n_31443), .b(n_31236), .o(n_31463) );
in01f80 newInst_574 ( .a(newNet_573), .o(newNet_574) );
no02f80 g762334 ( .a(n_18386), .b(n_18385), .o(n_18387) );
no02f80 g752983 ( .a(n_27086), .b(n_27156), .o(n_27236) );
na02f80 g768504 ( .a(n_12360), .b(FE_OCPN1002_n_45660), .o(n_12411) );
na02f80 g776967 ( .a(n_3879), .b(n_3840), .o(n_3880) );
no02f80 g768035 ( .a(FE_OCPN860_n_12880), .b(n_13073), .o(n_13113) );
na02f80 g751836 ( .a(n_28250), .b(n_28211), .o(n_28265) );
na02f80 g762102 ( .a(n_18177), .b(n_18060), .o(n_18195) );
in01f80 newInst_2206 ( .a(newNet_788), .o(newNet_2206) );
na02f80 g743981 ( .a(n_35691), .b(n_35663), .o(n_35746) );
in01f80 g736845 ( .a(n_43039), .o(n_43072) );
na02f80 g744249 ( .a(n_44180), .b(n_35521), .o(n_36184) );
in01f80 g763430 ( .a(n_17268), .o(n_17269) );
na02f80 g778470 ( .a(n_2582), .b(n_2542), .o(n_2640) );
in01f80 FE_OCP_RBC3578_n_8774 ( .a(n_8774), .o(FE_OCP_RBN3578_n_8774) );
na02f80 g738826 ( .a(n_41342), .b(n_41341), .o(n_41357) );
oa12f80 FE_RC_4165_0 ( .a(FE_RN_1814_0), .b(n_12574), .c(n_13059), .o(n_13232) );
oa22f80 g747683 ( .a(n_32260), .b(n_31989), .c(n_32261), .d(n_31988), .o(n_32325) );
no02f80 FE_RC_4177_0 ( .a(FE_RN_1822_0), .b(FE_RN_1823_0), .o(FE_RN_1824_0) );
na02f80 g755161 ( .a(n_25201), .b(n_24316), .o(n_25412) );
ao22s80 FE_RC_4266_0 ( .a(n_13577), .b(n_13630), .c(n_13629), .d(n_13593), .o(n_13722) );
no02f80 g760709 ( .a(n_19640), .b(FE_OCP_RBN1839_n_19528), .o(n_19700) );
in01f80 FE_OCPUNCOC1802_n_29375 ( .a(FE_OCPUNCON1801_n_29375), .o(FE_OCPUNCON1802_n_29375) );
in01f80 g744385 ( .a(n_46208), .o(n_36805) );
in01f80 g753979 ( .a(n_26278), .o(n_26279) );
in01f80 FE_OCP_RBC2602_n_39126 ( .a(n_39126), .o(FE_OCP_RBN2602_n_39126) );
in01f80 g747856 ( .a(n_33334), .o(n_33335) );
na02f80 g768385 ( .a(n_12467), .b(n_12440), .o(n_12441) );
no02f80 g751790 ( .a(n_28271), .b(n_28031), .o(n_28269) );
in01f80 g740164 ( .a(n_39950), .o(n_40041) );
na02f80 g770360 ( .a(n_10567), .b(n_10610), .o(n_10656) );
no02f80 g752060 ( .a(n_28982), .b(n_28669), .o(n_28690) );
no02f80 g749122 ( .a(n_30939), .b(n_27246), .o(n_30995) );
no02f80 g776579 ( .a(n_4360), .b(FE_OCP_RBN2528_n_3421), .o(n_4411) );
in01f80 g774901 ( .a(n_6261), .o(n_6262) );
na02f80 g738563 ( .a(n_41570), .b(n_41569), .o(n_41664) );
na02f80 g780587 ( .a(n_663), .b(n_554), .o(n_675) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_27_ ( .ck(newNet_1975), .d(n_12217), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_27_) );
no02f80 g771964 ( .a(n_44464), .b(n_9544), .o(n_9591) );
no02f80 g741331 ( .a(n_38869), .b(n_38842), .o(n_39033) );
in01f80 FE_RC_3272_0 ( .a(n_11426), .o(FE_RN_1441_0) );
no02f80 g762434 ( .a(FE_OCPN854_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_19_), .o(n_18005) );
no02f80 g770218 ( .a(n_10668), .b(n_10648), .o(n_10742) );
no02f80 g740024 ( .a(n_40008), .b(FE_OCP_RBN3715_n_39913), .o(n_40081) );
na02f80 g777332 ( .a(n_3564), .b(n_4587), .o(n_3566) );
na02f80 g771189 ( .a(n_9143), .b(n_9196), .o(n_9419) );
in01f80 FE_OCP_RBC3400_n_37670 ( .a(n_37670), .o(FE_OCP_RBN3400_n_37670) );
no02f80 g764273 ( .a(n_16290), .b(n_16237), .o(n_16407) );
na02f80 g761767 ( .a(n_18645), .b(n_18676), .o(n_18709) );
in01f80 FE_OCP_RBC1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01f80 newInst_2804 ( .a(newNet_2803), .o(newNet_2804) );
in01f80 g776599 ( .a(n_4391), .o(n_4392) );
in01f80 g743014 ( .a(n_36958), .o(n_36959) );
na02f80 g770485 ( .a(n_10367), .b(n_10325), .o(n_10483) );
na02f80 g749450 ( .a(n_30465), .b(n_30466), .o(n_30502) );
na02f80 g768821 ( .a(n_11822), .b(n_11883), .o(n_11980) );
na02f80 g769765 ( .a(n_11123), .b(n_11065), .o(n_11169) );
no02f80 g749926 ( .a(n_30262), .b(n_30214), .o(n_30243) );
in01f80 g761100 ( .a(n_19152), .o(n_19456) );
na02f80 g780827 ( .a(n_488), .b(n_458), .o(n_641) );
no02f80 g761025 ( .a(n_19315), .b(FE_OCP_DRV_N1554_n_19314), .o(n_19350) );
na02f80 g779642 ( .a(n_1480), .b(n_1479), .o(n_1499) );
no02f80 g780384 ( .a(n_937), .b(n_878), .o(n_879) );
oa22f80 FE_RC_1453_0 ( .a(n_32566), .b(n_32305), .c(n_28336), .d(n_32282), .o(n_32350) );
in01f80 FE_OCPC1451_n_27518 ( .a(n_27518), .o(FE_OCPN1451_n_27518) );
ao12f80 g772503 ( .a(n_8010), .b(n_8369), .c(n_7989), .o(n_8503) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_17_ ( .ck(newNet_2772), .d(n_46975), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_17_) );
na02f80 g740910 ( .a(n_39336), .b(n_39308), .o(n_40202) );
na02f80 g771669 ( .a(n_9097), .b(n_9005), .o(n_9203) );
na02f80 g745558 ( .a(n_34650), .b(n_34621), .o(n_34702) );
oa22f80 g753409 ( .a(n_26809), .b(n_26719), .c(n_26808), .d(n_26718), .o(n_26881) );
na02f80 g753437 ( .a(n_26964), .b(n_26962), .o(n_27041) );
na02f80 g742423 ( .a(FE_OCP_RBN2212_n_37720), .b(FE_OCP_RBN3400_n_37670), .o(n_37736) );
in01f80 newInst_1367 ( .a(newNet_392), .o(newNet_1367) );
oa12f80 g775211 ( .a(n_5951), .b(n_5950), .c(n_5949), .o(n_5992) );
no02f80 g743841 ( .a(n_37138), .b(n_36805), .o(n_37168) );
ao22s80 FE_RC_1352_0 ( .a(n_38778), .b(n_38610), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .d(n_38609), .o(n_38657) );
in01f80 FE_RC_1648_0 ( .a(n_20823), .o(FE_RN_460_0) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_13_ ( .ck(newNet_2213), .d(FE_OFN760_n_45813), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_13_) );
in01f80 FE_RC_3607_0 ( .a(FE_OCPN1483_n_18953), .o(FE_RN_1577_0) );
in01f80 g755282 ( .a(n_25686), .o(n_26417) );
no02f80 g742379 ( .a(n_37763), .b(n_37710), .o(n_37794) );
in01f80 g758698 ( .a(n_21843), .o(n_21844) );
na02f80 g766796 ( .a(n_14429), .b(n_14562), .o(n_14563) );
in01f80 g763585 ( .a(n_16899), .o(n_16973) );
na02f80 g770336 ( .a(FE_OCP_RBN2887_n_10570), .b(FE_OCP_RBN2874_n_10477), .o(n_10623) );
no02f80 g775580 ( .a(FE_OCP_RBN3695_n_5284), .b(n_4556), .o(n_5352) );
in01f80 g749193 ( .a(n_30887), .o(n_30852) );
no02f80 g742749 ( .a(n_37390), .b(n_37254), .o(n_37480) );
in01f80 g774827 ( .a(n_6386), .o(n_6310) );
in01f80 FE_RC_1870_0 ( .a(n_32598), .o(FE_RN_577_0) );
na02f80 g781229 ( .a(n_102), .b(n_61), .o(n_112) );
no02f80 g758057 ( .a(n_22688), .b(n_22843), .o(n_23448) );
no02f80 g760351 ( .a(n_20128), .b(n_19884), .o(n_20172) );
na03f80 FE_RC_2238_0 ( .a(FE_RN_817_0), .b(n_23437), .c(n_23438), .o(n_23494) );
in01f80 newInst_1466 ( .a(newNet_343), .o(newNet_1466) );
ao22s80 g779117 ( .a(n_1967), .b(n_1774), .c(n_1999), .d(n_1773), .o(n_2034) );
no02f80 g765898 ( .a(n_14826), .b(FE_OCPN1046_n_13570), .o(n_14854) );
in01f80 g765089 ( .a(n_15494), .o(n_15495) );
no02f80 g774362 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_11_), .o(n_6873) );
na02f80 g773409 ( .a(n_7518), .b(delay_add_ln22_unr5_stage3_stallmux_q_25_), .o(n_7567) );
in01f80 FE_OCPC3767_n_14439 ( .a(FE_OCPN3766_n_14439), .o(FE_OCPN3767_n_14439) );
na02f80 g750514 ( .a(n_29543), .b(n_29542), .o(n_29544) );
na02f80 g773971 ( .a(n_6931), .b(n_6987), .o(n_7008) );
na02f80 g751893 ( .a(n_29043), .b(n_29042), .o(n_29653) );
no02f80 g745031 ( .a(n_34859), .b(n_34564), .o(n_34901) );
no02f80 g784771 ( .a(n_20249), .b(FE_OCP_RBN1176_n_18981), .o(n_47257) );
no02f80 g742195 ( .a(n_44871), .b(n_37889), .o(n_37890) );
no02f80 g770889 ( .a(n_9992), .b(FE_OFN755_n_44461), .o(n_10050) );
in01f80 FE_OCP_RBC3065_n_22170 ( .a(FE_OCP_RBN3064_n_22170), .o(FE_OCP_RBN3065_n_22170) );
no02f80 g765972 ( .a(n_15090), .b(n_15063), .o(n_15064) );
in01f80 g743082 ( .a(n_36935), .o(n_36990) );
ao12f80 g756449 ( .a(n_24196), .b(n_24195), .c(n_24194), .o(n_25002) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_7_ ( .ck(newNet_396), .d(n_32515), .o(delay_xor_ln22_unr21_stage8_stallmux_q_7_) );
oa22f80 FE_RC_3374_0 ( .a(n_18630), .b(n_19539), .c(FE_RN_1464_0), .d(n_19519), .o(n_19663) );
in01f80 g753157 ( .a(n_27484), .o(n_27485) );
ao12f80 g741817 ( .a(n_38311), .b(n_38368), .c(n_38352), .o(n_38423) );
no02f80 g748064 ( .a(n_32882), .b(n_32881), .o(n_32883) );
in01f80 g777979 ( .a(n_47021), .o(n_3137) );
no02f80 g756637 ( .a(n_24190), .b(n_24189), .o(n_24191) );
in01f80 g742701 ( .a(n_37882), .o(n_38293) );
ao12f80 g765633 ( .a(n_15070), .b(n_15003), .c(n_14916), .o(n_15225) );
in01f80 g762617 ( .a(n_18021), .o(n_18043) );
oa12f80 g764767 ( .a(n_15494), .b(n_45136), .c(n_15492), .o(n_15768) );
na02f80 g778975 ( .a(n_2204), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_18_), .o(n_2263) );
in01f80 newInst_3581 ( .a(newNet_3580), .o(newNet_3581) );
na02f80 g776604 ( .a(n_4355), .b(n_4204), .o(n_4356) );
no02f80 g781255 ( .a(n_135), .b(n_71), .o(n_237) );
in01f80 g777719 ( .a(n_3331), .o(n_3332) );
na02f80 g758749 ( .a(n_21616), .b(n_21506), .o(n_21663) );
no02f80 g743555 ( .a(n_36444), .b(n_36095), .o(n_36462) );
in01f80 newInst_490 ( .a(newNet_489), .o(newNet_490) );
no02f80 g761866 ( .a(n_18786), .b(n_18593), .o(n_18675) );
no02f80 g772768 ( .a(n_7990), .b(n_7972), .o(n_9304) );
no02f80 FE_RC_3956_0 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .b(n_23581), .o(FE_RN_1714_0) );
in01f80 FE_OCP_RBC2699_n_4238 ( .a(FE_OCP_RBN2698_n_4238), .o(FE_OCP_RBN2699_n_4238) );
ao12f80 g737286 ( .a(n_42418), .b(n_42847), .c(n_42746), .o(n_42898) );
in01f80 g752236 ( .a(n_28058), .o(n_28184) );
na02f80 g756558 ( .a(n_23843), .b(delay_add_ln22_unr14_stage6_stallmux_q_28_), .o(n_23876) );
no02f80 g756168 ( .a(n_24101), .b(n_21852), .o(n_24146) );
no02f80 g764188 ( .a(n_16407), .b(n_16335), .o(n_16499) );
in01f80 g745589 ( .a(n_34324), .o(n_34290) );
no02f80 g749068 ( .a(n_30991), .b(n_27366), .o(n_31075) );
no02f80 g764729 ( .a(n_17158), .b(n_16503), .o(n_16540) );
na02f80 g765654 ( .a(n_15008), .b(n_15043), .o(n_15097) );
no04s80 g762135 ( .a(n_18137), .b(n_17977), .c(n_18115), .d(n_18026), .o(n_18177) );
in01f80 newInst_2355 ( .a(newNet_2354), .o(newNet_2355) );
in01f80 g780013 ( .a(n_1267), .o(n_1268) );
na02f80 g769558 ( .a(n_11349), .b(n_11304), .o(n_11354) );
ao12f80 g745566 ( .a(n_34157), .b(n_34250), .c(n_34197), .o(n_34298) );
oa22f80 g753613 ( .a(n_27202), .b(n_26889), .c(n_27201), .d(n_26888), .o(n_27323) );
no02f80 g751869 ( .a(n_28248), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .o(n_28371) );
na02f80 g758045 ( .a(n_22840), .b(n_22656), .o(n_22841) );
no02f80 g761198 ( .a(n_19083), .b(n_19082), .o(n_19084) );
no02f80 g776652 ( .a(n_4340), .b(n_4339), .o(n_4382) );
oa12f80 g766748 ( .a(n_13804), .b(n_13803), .c(n_13827), .o(n_13879) );
na02f80 g745933 ( .a(n_34064), .b(n_33942), .o(n_34065) );
oa12f80 g779193 ( .a(n_1848), .b(n_1847), .c(n_1846), .o(n_1908) );
in01f80 newInst_1529 ( .a(newNet_1012), .o(newNet_1529) );
in01f80 g756366 ( .a(n_23890), .o(n_23891) );
in01f80 newInst_800 ( .a(newNet_799), .o(newNet_800) );
in01f80 FE_RC_3258_0 ( .a(FE_RN_1305_0), .o(FE_RN_1437_0) );
ao12f80 g767909 ( .a(n_12392), .b(n_12615), .c(n_12420), .o(n_12655) );
na02f80 g780558 ( .a(n_662), .b(n_545), .o(n_670) );
na02f80 g752995 ( .a(n_27184), .b(n_27098), .o(n_27272) );
in01f80 g750556 ( .a(n_29425), .o(n_29426) );
ao12f80 g766750 ( .a(n_14012), .b(n_14011), .c(n_14010), .o(n_15788) );
in01f80 g741275 ( .a(n_39041), .o(n_38980) );
na02f80 g775319 ( .a(n_5901), .b(n_5558), .o(n_5974) );
no02f80 g771210 ( .a(n_9299), .b(FE_OCP_RBN2522_n_8951), .o(n_9416) );
no02f80 g739961 ( .a(n_40157), .b(n_40041), .o(n_40197) );
no02f80 g759951 ( .a(n_20753), .b(n_20667), .o(n_20815) );
na02f80 g768798 ( .a(n_12021), .b(delay_add_ln22_unr8_stage4_stallmux_q_3_), .o(n_12130) );
na02f80 g747799 ( .a(n_33372), .b(n_33370), .o(n_33702) );
no02f80 g753563 ( .a(n_26725), .b(n_26332), .o(n_26780) );
in01f80 g749496 ( .a(n_30500), .o(n_30510) );
no02f80 g773580 ( .a(n_45865), .b(n_7428), .o(n_7429) );
no02f80 g744077 ( .a(n_44222), .b(FE_OCP_RBN2615_n_35005), .o(n_36098) );
in01f80 g770679 ( .a(n_10349), .o(n_10350) );
no02f80 FE_RC_2500_0 ( .a(FE_RN_1013_0), .b(n_42038), .o(FE_RN_1014_0) );
no02f80 g753943 ( .a(FE_OCP_RBN2908_n_26173), .b(n_23398), .o(n_26260) );
in01f80 g747844 ( .a(n_32238), .o(n_32264) );
no02f80 g756301 ( .a(n_24609), .b(n_23911), .o(n_24668) );
in01f80 g750657 ( .a(n_29329), .o(n_29345) );
oa22f80 FE_RC_1328_0 ( .a(n_9669), .b(n_9718), .c(n_9668), .d(n_9719), .o(n_9859) );
in01f80 FE_OCP_RBC3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_ ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_) );
in01f80 FE_RC_3557_0 ( .a(FE_OCPN1464_n_29630), .o(FE_RN_1544_0) );
in01f80 g777105 ( .a(n_5384), .o(n_5341) );
no02f80 g773944 ( .a(n_6959), .b(n_6621), .o(n_7013) );
na02f80 g740333 ( .a(n_39995), .b(n_40269), .o(n_40392) );
in01f80 newInst_3318 ( .a(newNet_2895), .o(newNet_3318) );
in01f80 newInst_515 ( .a(newNet_514), .o(newNet_515) );
in01f80 newInst_916 ( .a(newNet_915), .o(newNet_916) );
na02f80 g741503 ( .a(n_38709), .b(n_38681), .o(n_38711) );
in01f80 g769716 ( .a(n_11229), .o(n_11271) );
ao12f80 g746700 ( .a(n_33026), .b(n_33039), .c(n_33025), .o(n_34222) );
na02f80 g750146 ( .a(n_29869), .b(n_29114), .o(n_29954) );
no02f80 g737950 ( .a(n_42201), .b(n_41948), .o(n_42372) );
no02f80 g747465 ( .a(FE_OCP_RBN3333_n_44962), .b(n_32543), .o(n_32593) );
na02f80 g750281 ( .a(n_29807), .b(n_29776), .o(n_29826) );
in01f80 newInst_2785 ( .a(newNet_2784), .o(newNet_2785) );
in01f80 newInst_112 ( .a(newNet_111), .o(newNet_112) );
in01f80 newInst_1218 ( .a(newNet_1217), .o(newNet_1218) );
in01f80 g757199 ( .a(n_23246), .o(n_23263) );
in01f80 newInst_730 ( .a(newNet_729), .o(newNet_730) );
oa22f80 g777224 ( .a(n_3564), .b(n_3195), .c(n_3596), .d(n_4761), .o(n_3733) );
na02f80 g780565 ( .a(n_666), .b(n_695), .o(n_700) );
ao12f80 g739390 ( .a(n_40849), .b(FE_OCPN897_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n_41306) );
no02f80 g758998 ( .a(n_21537), .b(n_45080), .o(n_21572) );
no02f80 g765241 ( .a(n_15126), .b(n_15191), .o(n_15343) );
no02f80 FE_RC_2708_0 ( .a(FE_RN_1137_0), .b(FE_RN_1138_0), .o(FE_RN_1139_0) );
ms00f80 mux_while_ln12_psv_q_reg_6_ ( .ck(newNet_104), .d(n_227), .o(mux_while_ln12_psv_q_6_) );
in01f80 newInst_3110 ( .a(newNet_3109), .o(newNet_3110) );
in01f80 g773239 ( .a(n_7639), .o(n_7640) );
in01f80 g747693 ( .a(n_33443), .o(n_33444) );
no02f80 FE_RC_2365_0 ( .a(n_1749), .b(FE_RN_915_0), .o(FE_RN_916_0) );
no02f80 FE_RC_1959_0 ( .a(n_14466), .b(FE_RN_631_0), .o(n_14503) );
no02f80 g737219 ( .a(n_42928), .b(n_42673), .o(n_42950) );
na02f80 g739153 ( .a(n_40960), .b(n_40882), .o(n_40961) );
in01f80 FE_OCP_RBC3140_n_6477 ( .a(n_6477), .o(FE_OCP_RBN3140_n_6477) );
in01f80 g761878 ( .a(n_18639), .o(n_18640) );
in01f80 g738727 ( .a(n_41502), .o(n_41457) );
na02f80 g770130 ( .a(n_10742), .b(FE_OCP_RBN2621_n_44561), .o(n_10782) );
na02f80 g748075 ( .a(n_32843), .b(n_32781), .o(n_32882) );
na02f80 g754923 ( .a(n_25270), .b(n_24305), .o(n_25421) );
no02f80 g779547 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_15_), .o(n_1770) );
na02f80 g745016 ( .a(n_34930), .b(n_34929), .o(n_34931) );
na03f80 g784143 ( .a(n_37897), .b(n_46252), .c(n_37898), .o(n_45890) );
no02f80 g763069 ( .a(n_17452), .b(n_17454), .o(n_17455) );
no02f80 g768318 ( .a(n_12545), .b(n_12544), .o(n_12546) );
na02f80 FE_RC_2904_0 ( .a(FE_RN_1258_0), .b(FE_RN_1260_0), .o(FE_RN_1261_0) );
no02f80 g740869 ( .a(n_39377), .b(n_39158), .o(n_39434) );
na03f80 FE_RC_1042_0 ( .a(FE_RN_302_0), .b(n_32689), .c(n_32851), .o(n_32889) );
no02f80 g757097 ( .a(n_23566), .b(n_23565), .o(n_23567) );
in01f80 FE_OCP_RBC2424_n_47023 ( .a(n_47023), .o(FE_OCP_RBN2424_n_47023) );
na02f80 g778069 ( .a(n_3024), .b(n_3023), .o(n_3101) );
na02f80 g767378 ( .a(n_13361), .b(n_13301), .o(n_13386) );
no02f80 g747587 ( .a(n_32333), .b(n_47271), .o(n_32366) );
no02f80 g763854 ( .a(n_16639), .b(n_15083), .o(n_16777) );
no02f80 g771676 ( .a(n_9240), .b(FE_OCP_RBN3549_n_44575), .o(n_9269) );
in01f80 g753418 ( .a(n_26882), .o(n_26852) );
na02f80 g764191 ( .a(n_16495), .b(n_16442), .o(n_16533) );
in01f80 FE_OFC785_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN782_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01f80 g761684 ( .a(n_18756), .o(n_18717) );
in01f80 g736282 ( .a(n_43894), .o(n_43895) );
no02f80 g749930 ( .a(n_30279), .b(n_30278), .o(n_30280) );
in01f80 g764654 ( .a(n_15948), .o(n_15993) );
no02f80 g784602 ( .a(n_11049), .b(n_44464), .o(n_44453) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_4_ ( .ck(newNet_299), .d(n_1328), .o(delay_xor_ln22_unr3_stage2_stallmux_q_4_) );
na02f80 g770606 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .o(n_10458) );
in01f80 g756014 ( .a(n_25191), .o(n_25166) );
ao12f80 g761361 ( .a(n_19676), .b(n_20086), .c(n_19650), .o(n_20120) );
na02f80 g777046 ( .a(n_3844), .b(n_3804), .o(n_4023) );
no02f80 g747330 ( .a(FE_OCP_RBN2103_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_6_), .o(n_32818) );
na02f80 g751561 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_20_), .o(n_28533) );
na02f80 g775411 ( .a(n_5444), .b(n_5494), .o(n_5495) );
in01f80 FE_OCP_RBC3475_n_7886 ( .a(FE_OCP_RBN3471_n_7886), .o(FE_OCP_RBN3475_n_7886) );
ao12f80 g745143 ( .a(n_34821), .b(n_34820), .c(n_34819), .o(n_34894) );
in01f80 g777668 ( .a(n_3478), .o(n_3479) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_6_ ( .ck(newNet_1000), .d(n_17144), .o(delay_xor_ln21_unr12_stage5_stallmux_q_6_) );
na02f80 g768584 ( .a(n_12234), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(n_12235) );
in01f80 g745759 ( .a(n_34198), .o(n_34199) );
na02f80 g775773 ( .a(n_5029), .b(FE_OCP_RBN2728_n_4219), .o(n_5204) );
oa12f80 g753732 ( .a(n_26335), .b(n_26377), .c(FE_OCPN1026_n_25481), .o(n_26502) );
in01f80 newInst_2941 ( .a(newNet_2175), .o(newNet_2941) );
in01f80 FE_OCP_RBC1354_n_33584 ( .a(FE_OCP_RBN1353_n_33584), .o(FE_OCP_RBN1354_n_33584) );
no02f80 g765400 ( .a(n_15186), .b(n_15149), .o(n_15338) );
in01f80 newInst_2328 ( .a(newNet_2327), .o(newNet_2328) );
in01f80 g743572 ( .a(n_36545), .o(n_36581) );
in01f80 g747817 ( .a(n_33313), .o(n_33516) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_7_ ( .ck(newNet_1791), .d(n_16414), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_) );
in01f80 newInst_2482 ( .a(newNet_35), .o(newNet_2482) );
in01f80 g771040 ( .a(n_9747), .o(n_9748) );
no02f80 g753137 ( .a(n_27390), .b(n_27345), .o(n_27494) );
na02f80 g743259 ( .a(n_36844), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_), .o(n_36864) );
na02f80 g779770 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_), .o(n_1479) );
oa12f80 g777635 ( .a(n_2954), .b(n_3423), .c(n_2781), .o(n_3466) );
no02f80 g743967 ( .a(n_35909), .b(n_35911), .o(n_35952) );
na02f80 g743426 ( .a(n_36628), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36671) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_29_ ( .ck(newNet_1709), .d(n_22659), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_) );
in01f80 FE_OCPC1481_n_22207 ( .a(n_22207), .o(FE_OCPN1481_n_22207) );
in01f80 g750940 ( .a(n_29054), .o(n_29080) );
in01f80 FE_RC_2630_0 ( .a(FE_RN_1095_0), .o(n_12420) );
no02f80 g742102 ( .a(n_37874), .b(n_37889), .o(n_37909) );
no02f80 g762828 ( .a(n_17889), .b(n_17885), .o(n_17907) );
in01f80 g743617 ( .a(n_37517), .o(n_37586) );
in01f80 newInst_2168 ( .a(newNet_2167), .o(newNet_2168) );
in01f80 g754708 ( .a(n_26345), .o(n_26866) );
no02f80 g758330 ( .a(n_22187), .b(n_21324), .o(n_22292) );
in01f80 g780404 ( .a(n_800), .o(n_801) );
oa22f80 FE_RC_3745_0 ( .a(n_25831), .b(n_25816), .c(FE_OCPN1748_n_23354), .d(FE_OCP_RBN1139_n_25816), .o(n_25912) );
na02f80 g755123 ( .a(n_25315), .b(n_24310), .o(n_25349) );
in01f80 newInst_3105 ( .a(newNet_3104), .o(newNet_3105) );
in01f80 FE_OCPC1799_FE_OFN780_n_17093 ( .a(FE_OFN780_n_17093), .o(FE_OCPN1799_FE_OFN780_n_17093) );
oa22f80 g737654 ( .a(FE_OCPN887_n_42367), .b(n_42459), .c(n_42392), .d(n_42483), .o(n_42797) );
na02f80 g777130 ( .a(n_3671), .b(n_3695), .o(n_3770) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_11_ ( .ck(newNet_3655), .d(n_16425), .o(delay_add_ln22_unr11_stage5_stallmux_q_11_) );
in01f80 newInst_3754 ( .a(newNet_3753), .o(newNet_3754) );
in01f80 g749894 ( .a(n_31276), .o(n_31342) );
na02f80 g749078 ( .a(n_30954), .b(n_31655), .o(n_30989) );
na02f80 g780904 ( .a(n_420), .b(n_465), .o(n_581) );
in01f80 newInst_1487 ( .a(newNet_1486), .o(newNet_1487) );
in01f80 g776071 ( .a(n_5093), .o(n_5094) );
in01f80 g750564 ( .a(n_29481), .o(n_29473) );
in01f80 g776559 ( .a(n_4424), .o(n_4425) );
ao12f80 g762703 ( .a(n_17872), .b(FE_OCP_RBN2148_FE_OCPN861_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_16_), .o(n_17918) );
in01f80 g780799 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_1_), .o(n_607) );
no02f80 g740066 ( .a(n_40116), .b(n_40009), .o(n_40010) );
in01f80 g780282 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n_792) );
in01f80 g740304 ( .a(n_39816), .o(n_39913) );
ao12f80 g782658 ( .a(n_15142), .b(n_15228), .c(n_14239), .o(n_44051) );
in01f80 g737435 ( .a(n_42738), .o(n_42734) );
no02f80 g737711 ( .a(n_42392), .b(n_42421), .o(n_42467) );
in01f80 newInst_3063 ( .a(newNet_2112), .o(newNet_3063) );
no02f80 g769054 ( .a(FE_OCP_RBN3270_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_4_), .o(n_11737) );
in01f80 g769163 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_0_), .o(n_11592) );
no02f80 g754950 ( .a(n_25210), .b(n_24221), .o(n_25272) );
in01f80 newInst_187 ( .a(newNet_137), .o(newNet_187) );
na02f80 g773094 ( .a(n_7641), .b(n_8226), .o(n_7656) );
ao12f80 g750488 ( .a(n_29466), .b(n_29558), .c(n_29516), .o(n_29564) );
oa12f80 g757528 ( .a(n_23321), .b(n_23320), .c(n_23319), .o(n_23801) );
na02f80 g759941 ( .a(n_21374), .b(n_21595), .o(n_21668) );
no02f80 g763809 ( .a(n_17106), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_), .o(n_17107) );
ao12f80 g773112 ( .a(n_7806), .b(n_8232), .c(n_7215), .o(n_8556) );
na02f80 g775123 ( .a(n_5870), .b(n_5766), .o(n_5871) );
na02f80 FE_RC_2858_0 ( .a(FE_OFN755_n_44461), .b(n_10270), .o(FE_RN_1231_0) );
na02f80 g752049 ( .a(n_28714), .b(n_28713), .o(n_28715) );
no02f80 g763766 ( .a(n_16748), .b(n_16777), .o(n_16778) );
na02f80 g777146 ( .a(n_3679), .b(n_3653), .o(n_3695) );
no02f80 g750640 ( .a(n_29271), .b(n_29379), .o(n_29304) );
no02f80 g772521 ( .a(n_8419), .b(n_8455), .o(n_8456) );
in01f80 FE_RC_2495_0 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_2_), .o(FE_RN_1011_0) );
oa12f80 g759527 ( .a(FE_OCP_RBN3612_FE_OCPN1797_n_20333), .b(n_20767), .c(n_20332), .o(n_20799) );
no02f80 g753539 ( .a(n_26757), .b(n_26780), .o(n_26874) );
in01f80 g769016 ( .a(n_11761), .o(n_11842) );
na02f80 g763352 ( .a(FE_OCP_RBN3205_n_44365), .b(n_16881), .o(n_17040) );
in01f80 g779210 ( .a(n_1959), .o(n_1934) );
na02f80 FE_RC_2074_0 ( .a(FE_RN_707_0), .b(n_30558), .o(n_30603) );
in01f80 g773073 ( .a(n_8048), .o(n_8049) );
in01f80 FE_OCP_RBC3604_n_8981 ( .a(n_8981), .o(FE_OCP_RBN3604_n_8981) );
in01f80 g774782 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_22_), .o(n_7467) );
na02f80 g742261 ( .a(n_44875), .b(n_37511), .o(n_38120) );
no02f80 g760398 ( .a(n_20167), .b(FE_OCPN1438_FE_OCP_RBN1330_n_18866), .o(n_20168) );
in01f80 FE_OCPC1241_n_7721 ( .a(FE_OCPN1240_n_7721), .o(FE_OCPN1241_n_7721) );
in01f80 g766560 ( .a(n_13928), .o(n_13929) );
in01f80 g756077 ( .a(n_24208), .o(n_24209) );
in01f80 g766533 ( .a(n_14564), .o(n_14621) );
in01f80 g769052 ( .a(n_11882), .o(n_11692) );
na02f80 g765052 ( .a(n_15533), .b(n_15532), .o(n_15534) );
in01f80 g741005 ( .a(n_39109), .o(n_39083) );
in01f80 fopt783279 ( .a(n_10599), .o(n_44853) );
na02f80 g763690 ( .a(n_16739), .b(FE_OCP_RBN2787_n_15079), .o(n_16809) );
in01f80 FE_OCPC1252_n_8348 ( .a(n_8348), .o(FE_OCPN1252_n_8348) );
oa12f80 g745248 ( .a(n_34119), .b(n_34275), .c(n_34149), .o(n_34520) );
in01f80 g749310 ( .a(n_30676), .o(n_30677) );
na02f80 FE_RC_3927_0 ( .a(n_11774), .b(FE_RN_1698_0), .o(n_11817) );
oa12f80 g773381 ( .a(n_7557), .b(n_7558), .c(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n_7590) );
in01f80 newInst_2724 ( .a(newNet_2723), .o(newNet_2724) );
in01f80 FE_RC_2609_0 ( .a(n_17977), .o(FE_RN_1085_0) );
in01f80 newInst_437 ( .a(newNet_436), .o(newNet_437) );
no02f80 FE_RC_2570_0 ( .a(n_12620), .b(FE_RN_1055_0), .o(n_13413) );
na02f80 g740412 ( .a(FE_OCP_RBN3022_n_39942), .b(n_39582), .o(n_40054) );
in01f80 g737335 ( .a(n_42856), .o(n_43172) );
oa22f80 g739977 ( .a(n_39875), .b(n_39814), .c(n_39874), .d(n_39815), .o(n_39958) );
in01f80 newInst_1605 ( .a(newNet_1009), .o(newNet_1605) );
in01f80 g763386 ( .a(n_16957), .o(n_17037) );
na02f80 g780509 ( .a(n_674), .b(n_670), .o(n_714) );
in01f80 g747467 ( .a(n_32578), .o(n_32595) );
in01f80 g748195 ( .a(n_31742), .o(n_31774) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_11_ ( .ck(newNet_2880), .d(n_10885), .o(delay_add_ln22_unr8_stage4_stallmux_q_11_) );
in01f80 FE_OCP_RBC2867_n_16088 ( .a(n_16088), .o(FE_OCP_RBN2867_n_16088) );
in01f80 g745817 ( .a(n_34203), .o(n_34179) );
no02f80 g748799 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_25_), .o(n_32461) );
no02f80 g755609 ( .a(n_24596), .b(n_24615), .o(n_24748) );
in01f80 newInst_2511 ( .a(newNet_2510), .o(newNet_2511) );
na02f80 g765272 ( .a(FE_OCP_RBN2673_n_14991), .b(n_14758), .o(n_15058) );
ao22s80 g779513 ( .a(n_1372), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln22_unr3_stage2_stallmux_q_5_), .o(n_1453) );
na03f80 FE_RC_161_0 ( .a(n_17560), .b(n_17561), .c(n_17458), .o(n_17683) );
in01f80 g748314 ( .a(n_31842), .o(n_31843) );
ao22s80 g756629 ( .a(n_23474), .b(n_23544), .c(n_23473), .d(n_23579), .o(n_25022) );
in01f80 g761452 ( .a(n_20133), .o(n_20134) );
no02f80 g748183 ( .a(n_31684), .b(n_31704), .o(n_31808) );
no02f80 g776323 ( .a(n_4762), .b(n_4761), .o(n_4919) );
na02f80 FE_RC_1076_0 ( .a(n_12541), .b(n_12542), .o(FE_RN_318_0) );
in01f80 FE_OCP_RBC3601_FE_OCPN1243_n_44460 ( .a(FE_OCP_RBN3598_FE_OCPN1243_n_44460), .o(FE_OCP_RBN3601_FE_OCPN1243_n_44460) );
no02f80 g745398 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35840), .o(n_35958) );
in01f80 g764341 ( .a(n_16424), .o(n_16456) );
na02f80 g738585 ( .a(n_41536), .b(n_41187), .o(n_41566) );
oa12f80 g739065 ( .a(n_40926), .b(n_41031), .c(n_40797), .o(n_41073) );
na02f80 FE_RC_559_0 ( .a(FE_RN_168_0), .b(FE_RN_169_0), .o(FE_RN_170_0) );
in01f80 newInst_2102 ( .a(newNet_2101), .o(newNet_2102) );
in01f80 g745214 ( .a(n_36228), .o(n_36178) );
na02f80 g775246 ( .a(n_6002), .b(n_6001), .o(n_6003) );
oa22f80 g752450 ( .a(n_27639), .b(n_27423), .c(n_45638), .d(n_27424), .o(n_27739) );
in01f80 FE_OCP_RBC3646_n_44490 ( .a(FE_OCP_RBN3641_n_44490), .o(FE_OCP_RBN3646_n_44490) );
in01f80 g758651 ( .a(n_22032), .o(n_22033) );
no02f80 g767011 ( .a(FE_OCP_RBN2503_n_13896), .b(n_13975), .o(n_14137) );
no02f80 g752785 ( .a(n_27881), .b(n_27903), .o(n_27905) );
no02f80 g754141 ( .a(n_26004), .b(n_26003), .o(n_26068) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_6_ ( .ck(newNet_1794), .d(n_16413), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_6_) );
in01f80 newInst_1787 ( .a(newNet_1786), .o(newNet_1787) );
in01f80 g771598 ( .a(n_9268), .o(n_9335) );
in01f80 g743451 ( .a(n_36583), .o(n_36584) );
no02f80 g738502 ( .a(FE_OCPN953_n_41540), .b(n_41406), .o(n_41743) );
in01f80 FE_OCP_RBC3513_n_13960 ( .a(FE_OCP_RBN2411_n_13960), .o(FE_OCP_RBN3513_n_13960) );
in01f80 g751391 ( .a(n_28705), .o(n_28770) );
no03m80 FE_RC_2277_0 ( .a(n_17533), .b(FE_RN_849_0), .c(n_18237), .o(n_45524) );
na02f80 g749361 ( .a(n_30724), .b(FE_RN_1486_0), .o(n_30791) );
no02f80 g784413 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_21_), .o(n_46225) );
oa12f80 g743627 ( .a(n_36105), .b(n_36410), .c(n_47266), .o(n_36457) );
no02f80 g761880 ( .a(n_18994), .b(n_18993), .o(n_18995) );
in01f80 g747258 ( .a(n_33764), .o(n_33765) );
no02f80 g750368 ( .a(n_30663), .b(n_30084), .o(n_30662) );
in01f80 g766163 ( .a(n_14678), .o(n_14679) );
in01f80 FE_OCP_RBC3600_FE_OCPN1243_n_44460 ( .a(FE_OCP_RBN3598_FE_OCPN1243_n_44460), .o(FE_OCP_RBN3600_FE_OCPN1243_n_44460) );
in01f80 newInst_162 ( .a(newNet_161), .o(newNet_162) );
no02f80 g766725 ( .a(n_13732), .b(n_13261), .o(n_13759) );
in01f80 g752152 ( .a(n_28040), .o(n_28041) );
na02f80 g762964 ( .a(n_17509), .b(n_17518), .o(n_17656) );
na02f80 g770320 ( .a(n_10614), .b(n_10665), .o(n_10692) );
na02f80 FE_RC_1748_0 ( .a(FE_RN_489_0), .b(FE_RN_492_0), .o(n_44426) );
in01f80 newInst_2586 ( .a(newNet_2585), .o(newNet_2586) );
in01f80 newInst_2655 ( .a(newNet_2654), .o(newNet_2655) );
na02f80 g771583 ( .a(n_9025), .b(n_9007), .o(n_9079) );
na02f80 g771237 ( .a(n_9148), .b(FE_OCP_RBN2524_n_8951), .o(n_9155) );
oa12f80 g770521 ( .a(n_10398), .b(n_10474), .c(n_10286), .o(n_10525) );
in01f80 g754725 ( .a(n_26636), .o(n_26709) );
no02f80 g745749 ( .a(n_34201), .b(n_34200), .o(n_34202) );
no02f80 g743471 ( .a(n_37712), .b(n_36941), .o(n_37787) );
in01f80 g753090 ( .a(n_27274), .o(n_27229) );
ao12f80 g764755 ( .a(n_15725), .b(n_15889), .c(n_15793), .o(n_16030) );
no02f80 g751165 ( .a(n_29944), .b(n_29767), .o(n_30088) );
in01f80 g741183 ( .a(n_39358), .o(n_39359) );
oa12f80 g754491 ( .a(n_26383), .b(n_26349), .c(n_26160), .o(n_26454) );
oa22f80 g753508 ( .a(n_27451), .b(n_26895), .c(n_27452), .d(n_26894), .o(n_27539) );
in01f80 FE_RC_2526_0 ( .a(n_23003), .o(FE_RN_1030_0) );
in01f80 g743337 ( .a(n_36677), .o(n_36696) );
in01f80 newInst_3040 ( .a(newNet_3039), .o(newNet_3040) );
oa12f80 g746364 ( .a(n_33472), .b(n_33471), .c(n_33470), .o(n_33545) );
in01f80 newInst_2967 ( .a(newNet_228), .o(newNet_2967) );
in01f80 newInst_1046 ( .a(newNet_42), .o(newNet_1046) );
no02f80 g769780 ( .a(n_11113), .b(n_10984), .o(n_11172) );
oa12f80 g746373 ( .a(n_33537), .b(n_33536), .c(n_33535), .o(n_33604) );
in01f80 FE_OCP_RBC2270_n_13489 ( .a(n_13489), .o(FE_OCP_RBN2270_n_13489) );
ao12f80 g768104 ( .a(n_12632), .b(n_12589), .c(n_12631), .o(n_12694) );
in01f80 g761216 ( .a(n_19058), .o(n_19078) );
in01f80 g765558 ( .a(n_15258), .o(n_15178) );
na02f80 g747327 ( .a(n_32624), .b(n_44962), .o(n_32855) );
no02f80 g739004 ( .a(n_41192), .b(n_40775), .o(n_41204) );
oa12f80 g765863 ( .a(n_14967), .b(n_15032), .c(n_14966), .o(n_15093) );
in01f80 FE_RC_3900_0 ( .a(n_29697), .o(FE_RN_1694_0) );
na02f80 FE_RC_2600_0 ( .a(FE_RN_1075_0), .b(FE_RN_1078_0), .o(n_3564) );
na02f80 g737569 ( .a(n_42224), .b(n_42239), .o(n_42290) );
na02f80 g747517 ( .a(n_33398), .b(n_33315), .o(n_33446) );
in01f80 g750030 ( .a(n_31038), .o(n_31039) );
in01f80 g759156 ( .a(n_21127), .o(n_21128) );
in01f80 g767756 ( .a(n_13278), .o(n_13279) );
in01f80 newInst_2443 ( .a(newNet_2442), .o(newNet_2443) );
oa12f80 g747877 ( .a(n_32138), .b(n_32073), .c(n_32110), .o(n_32214) );
in01f80 g751581 ( .a(n_28842), .o(n_28843) );
na02f80 g777940 ( .a(n_3137), .b(FE_OCPN848_n_3597), .o(n_3194) );
ao12f80 g762424 ( .a(n_18328), .b(n_18327), .c(n_18326), .o(n_18414) );
in01f80 newInst_3184 ( .a(newNet_2619), .o(newNet_3184) );
in01f80 newInst_2090 ( .a(newNet_1730), .o(newNet_2090) );
na02f80 g753178 ( .a(n_27207), .b(n_25789), .o(n_27421) );
ao22s80 FE_RC_841_0 ( .a(n_44575), .b(FE_OCP_RBN3603_n_8981), .c(FE_OCP_RBN3572_n_44563), .d(n_8981), .o(n_9102) );
ao22s80 g763454 ( .a(n_17577), .b(n_17527), .c(n_17503), .d(n_17526), .o(n_18419) );
na02f80 FE_RC_2479_0 ( .a(n_40054), .b(n_40100), .o(FE_RN_1000_0) );
na02f80 g745164 ( .a(n_36056), .b(n_36112), .o(n_36252) );
in01f80 g756808 ( .a(n_23439), .o(n_23453) );
no02f80 g754157 ( .a(n_25983), .b(n_24218), .o(n_26293) );
in01f80 FE_OFC84_n_46137 ( .a(FE_OFN773_n_46137), .o(FE_OFN84_n_46137) );
in01f80 newInst_1758 ( .a(newNet_1757), .o(newNet_1758) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_10_ ( .ck(newNet_2221), .d(n_990), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_) );
in01f80 newInst_1943 ( .a(newNet_711), .o(newNet_1943) );
na02f80 g736819 ( .a(n_43048), .b(n_43052), .o(n_43053) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_6_ ( .ck(newNet_2903), .d(n_5273), .o(delay_add_ln22_unr5_stage3_stallmux_q_6_) );
ao12f80 g768377 ( .a(n_11898), .b(n_12413), .c(n_11960), .o(n_12486) );
in01f80 newInst_1456 ( .a(newNet_1455), .o(newNet_1456) );
in01f80 g774195 ( .a(n_7154), .o(n_7155) );
no02f80 g776238 ( .a(n_4508), .b(n_4550), .o(n_4647) );
no02f80 FE_RC_4239_0 ( .a(n_21490), .b(n_21572), .o(FE_RN_1862_0) );
in01f80 g741153 ( .a(n_38836), .o(n_38821) );
na02f80 g763959 ( .a(n_16606), .b(n_16605), .o(n_16686) );
ao12f80 g768861 ( .a(n_11458), .b(n_44355), .c(n_11658), .o(n_11947) );
na02f80 g763592 ( .a(n_16892), .b(n_16972), .o(n_17192) );
na02f80 g769817 ( .a(n_11164), .b(n_44454), .o(n_11181) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_31_ ( .ck(newNet_2526), .d(n_27781), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_31_) );
in01f80 newInst_2054 ( .a(newNet_2053), .o(newNet_2054) );
in01f80 fopt783523 ( .a(n_15510), .o(n_45134) );
in01f80 g759021 ( .a(n_21283), .o(n_21324) );
no02f80 g759581 ( .a(n_20685), .b(n_20474), .o(n_20821) );
in01f80 g740706 ( .a(n_39584), .o(n_39583) );
in01f80 newInst_335 ( .a(newNet_334), .o(newNet_335) );
in01f80 g751528 ( .a(n_29359), .o(n_29335) );
no02f80 g736870 ( .a(n_43470), .b(n_43503), .o(n_43609) );
na02f80 FE_RC_1161_0 ( .a(FE_RN_348_0), .b(FE_RN_349_0), .o(FE_RN_350_0) );
in01f80 g767831 ( .a(n_12727), .o(n_12751) );
in01f80 g779792 ( .a(n_1506), .o(n_1420) );
in01f80 g744108 ( .a(n_35574), .o(n_35593) );
in01f80 g746592 ( .a(n_34756), .o(n_34805) );
na02f80 g771427 ( .a(FE_OCP_RBN2543_n_9082), .b(n_9012), .o(n_9193) );
na02f80 g736762 ( .a(n_43110), .b(n_43106), .o(n_43112) );
in01f80 g743578 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .o(n_36461) );
no02f80 FE_RC_1871_0 ( .a(FE_RN_576_0), .b(FE_RN_577_0), .o(FE_RN_578_0) );
na02f80 g763671 ( .a(n_17372), .b(n_17257), .o(n_17374) );
in01f80 newInst_865 ( .a(newNet_864), .o(newNet_865) );
ao12f80 g775568 ( .a(n_5580), .b(n_5590), .c(n_5579), .o(n_5676) );
no02f80 g769260 ( .a(n_11585), .b(n_10613), .o(n_11584) );
oa22f80 g758662 ( .a(n_22286), .b(n_21821), .c(n_22287), .d(n_21822), .o(n_22398) );
na02f80 g766050 ( .a(n_14949), .b(n_14428), .o(n_15090) );
na02f80 g765493 ( .a(n_15719), .b(n_15957), .o(n_16255) );
in01f80 newInst_56 ( .a(newNet_42), .o(newNet_56) );
na02f80 g739338 ( .a(n_40676), .b(delay_add_ln22_unr27_stage10_stallmux_q_3_), .o(n_40742) );
in01f80 g754829 ( .a(n_26005), .o(n_26006) );
na02f80 g745223 ( .a(n_34520), .b(n_34519), .o(n_34521) );
in01f80 g749713 ( .a(n_31395), .o(n_31457) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_23_ ( .ck(newNet_2743), .d(n_17591), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_) );
in01f80 FE_OCP_RBC1326_n_36489 ( .a(n_36489), .o(FE_OCP_RBN1326_n_36489) );
in01f80 g754371 ( .a(n_26646), .o(n_26613) );
no02f80 g770408 ( .a(n_10330), .b(n_10442), .o(n_10506) );
no02f80 g741084 ( .a(n_39154), .b(n_39180), .o(n_39249) );
na02f80 g767006 ( .a(FE_OCP_RBN2503_n_13896), .b(n_14038), .o(n_14213) );
no02f80 g778463 ( .a(n_2694), .b(n_2109), .o(n_2722) );
in01f80 g741500 ( .a(n_38786), .o(n_38787) );
na02f80 g773530 ( .a(n_7477), .b(n_7476), .o(n_7478) );
oa12f80 g746094 ( .a(FE_OCP_RBN2169_n_32892), .b(n_33677), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_30_), .o(n_33719) );
oa22f80 g766858 ( .a(n_13869), .b(FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__), .c(n_13870), .d(FE_OCP_RBN1923_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_14044) );
na02f80 g767787 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n_12900) );
no02f80 g737934 ( .a(n_42180), .b(n_41516), .o(n_42207) );
no02f80 g780748 ( .a(n_590), .b(n_587), .o(n_588) );
in01f80 g774398 ( .a(n_6643), .o(n_6587) );
in01f80 g765744 ( .a(n_14959), .o(n_14960) );
oa12f80 g741697 ( .a(n_38089), .b(n_38478), .c(n_37949), .o(n_38521) );
na02f80 g773861 ( .a(n_7071), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_10_), .o(n_7134) );
in01f80 g778309 ( .a(n_2895), .o(n_2946) );
no02f80 g746796 ( .a(n_32963), .b(n_32962), .o(n_32974) );
in01f80 newInst_1206 ( .a(newNet_1205), .o(newNet_1206) );
no02f80 FE_RC_3303_0 ( .a(n_17972), .b(FE_RN_1454_0), .o(n_18077) );
in01f80 FE_OCP_RBC3272_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3272_n_45224) );
in01f80 g751540 ( .a(n_28494), .o(n_28495) );
no02f80 FE_RC_973_0 ( .a(n_26302), .b(FE_RN_281_0), .o(n_26327) );
no02f80 FE_RC_1240_0 ( .a(n_8806), .b(n_8815), .o(FE_RN_373_0) );
in01f80 newInst_1692 ( .a(newNet_1691), .o(newNet_1692) );
in01f80 newInst_3727 ( .a(newNet_3726), .o(newNet_3727) );
na02f80 g744282 ( .a(n_44180), .b(n_35684), .o(n_35780) );
in01f80 g745059 ( .a(n_36315), .o(n_36386) );
oa12f80 g738884 ( .a(n_41250), .b(n_41249), .c(n_41248), .o(n_41562) );
no02f80 g778985 ( .a(n_2201), .b(n_1947), .o(n_2214) );
in01f80 g775777 ( .a(n_5563), .o(n_5564) );
in01f80 g768023 ( .a(n_13080), .o(n_12988) );
no02f80 g751205 ( .a(n_29818), .b(n_29360), .o(n_30307) );
na02f80 g783821 ( .a(n_2575), .b(n_2349), .o(n_45506) );
no02f80 g738139 ( .a(n_42018), .b(n_42017), .o(n_42019) );
in01f80 g744136 ( .a(n_35737), .o(n_35738) );
in01f80 g746744 ( .a(n_34227), .o(n_34228) );
no02f80 g765193 ( .a(n_15828), .b(n_15839), .o(n_15880) );
in01f80 newInst_1533 ( .a(newNet_1532), .o(newNet_1533) );
na02f80 g775347 ( .a(n_5876), .b(n_5659), .o(n_5826) );
no02f80 g740783 ( .a(n_39442), .b(n_39407), .o(n_39891) );
in01f80 g741723 ( .a(n_38546), .o(n_38547) );
ao12f80 g755341 ( .a(n_24837), .b(n_24784), .c(n_24760), .o(n_24861) );
oa12f80 g739710 ( .a(n_40337), .b(n_40505), .c(n_40113), .o(n_40517) );
na02f80 g761730 ( .a(n_18679), .b(n_18646), .o(n_18824) );
na02f80 g768859 ( .a(n_11791), .b(n_11664), .o(n_11914) );
in01f80 fopt782735 ( .a(n_28319), .o(n_44143) );
na02f80 g740971 ( .a(n_39191), .b(n_39130), .o(n_39192) );
ao12f80 g761645 ( .a(n_19487), .b(n_19486), .c(n_19485), .o(n_19927) );
in01f80 g739084 ( .a(n_41096), .o(n_41097) );
no02f80 g771955 ( .a(FE_OFN754_n_44461), .b(n_9381), .o(n_9547) );
in01f80 g744874 ( .a(n_35130), .o(n_35165) );
na02f80 g777927 ( .a(n_3096), .b(n_45194), .o(n_3097) );
in01f80 newInst_2633 ( .a(newNet_2632), .o(newNet_2633) );
no02f80 g776337 ( .a(n_4810), .b(n_3715), .o(n_4949) );
in01f80 FE_OCP_DRV_C1549_n_19053 ( .a(n_19053), .o(FE_OCP_DRV_N1549_n_19053) );
no02f80 g776648 ( .a(n_4436), .b(n_4435), .o(n_4589) );
na02f80 g741175 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39230), .o(n_39303) );
ms00f80 sin_out_reg_20_ ( .ck(newNet_59), .d(n_43888), .o(sin_out_20) );
oa12f80 g747752 ( .a(n_32027), .b(n_32188), .c(n_31949), .o(n_32300) );
na02f80 g758936 ( .a(n_21237), .b(n_45070), .o(n_21329) );
in01f80 g771476 ( .a(n_8943), .o(n_8944) );
no02f80 g753808 ( .a(n_26328), .b(n_44443), .o(n_26411) );
in01f80 g759576 ( .a(n_20621), .o(n_20649) );
na02f80 g738190 ( .a(n_41990), .b(n_41729), .o(n_42033) );
in01f80 g763001 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .o(n_18367) );
na02f80 g776060 ( .a(n_4990), .b(n_4787), .o(n_5020) );
oa12f80 g771416 ( .a(n_9444), .b(n_9443), .c(n_9506), .o(n_9655) );
na02f80 g754166 ( .a(n_26076), .b(n_26036), .o(n_26138) );
in01f80 newInst_41 ( .a(newNet_40), .o(newNet_41) );
in01f80 g755765 ( .a(n_24461), .o(n_24486) );
no02f80 g744323 ( .a(FE_OCP_RBN2885_n_35517), .b(n_35516), .o(n_35645) );
na02f80 g755895 ( .a(n_24362), .b(n_24361), .o(n_24393) );
na02f80 g773952 ( .a(n_6914), .b(n_5312), .o(n_7016) );
in01f80 FE_OCPC1253_n_8348 ( .a(FE_OCPN1252_n_8348), .o(FE_OCPN1253_n_8348) );
na02f80 FE_RC_1918_0 ( .a(FE_RN_604_0), .b(n_18354), .o(FE_RN_605_0) );
no02f80 g755044 ( .a(n_25293), .b(FE_OCP_RBN1130_n_24179), .o(n_25294) );
no02f80 g772865 ( .a(n_8064), .b(n_8063), .o(n_8065) );
na02f80 FE_RC_3712_0 ( .a(FE_RN_1631_0), .b(FE_RN_1632_0), .o(FE_RN_1633_0) );
na02f80 g766819 ( .a(n_14306), .b(n_14561), .o(n_14352) );
na02f80 FE_RC_4154_0 ( .a(FE_RN_1806_0), .b(FE_RN_1807_0), .o(FE_RN_161_0) );
in01f80 newInst_1520 ( .a(newNet_1519), .o(newNet_1520) );
na02f80 g776799 ( .a(n_4155), .b(n_4175), .o(n_4156) );
oa12f80 g770348 ( .a(n_10393), .b(n_10659), .c(n_10380), .o(n_10740) );
no02f80 g738712 ( .a(n_41713), .b(n_41198), .o(n_41803) );
na02f80 FE_RC_3631_0 ( .a(FE_RN_1591_0), .b(n_13669), .o(n_13827) );
in01f80 FE_OCPC1769_delay_sub_ln23_0_unr23_stage8_stallmux_q ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(FE_OCPN1769_delay_sub_ln23_0_unr23_stage8_stallmux_q) );
no02f80 g755439 ( .a(n_24704), .b(n_24726), .o(n_24756) );
in01f80 g756136 ( .a(n_25032), .o(n_25026) );
no02f80 g768920 ( .a(n_11881), .b(n_11844), .o(n_11907) );
na02f80 g763800 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_28_), .o(n_17467) );
in01f80 g779351 ( .a(n_2343), .o(n_1687) );
oa22f80 g752708 ( .a(n_27932), .b(n_28021), .c(n_27997), .d(n_28022), .o(n_28993) );
oa22f80 g756533 ( .a(n_23843), .b(delay_add_ln22_unr14_stage6_stallmux_q_31_), .c(n_23572), .d(n_22929), .o(n_24048) );
oa22f80 FE_RC_1461_0 ( .a(n_17336), .b(n_17459), .c(n_17753), .d(n_17441), .o(n_17552) );
in01f80 g776621 ( .a(n_4111), .o(n_4112) );
no02f80 g776180 ( .a(n_4505), .b(n_4564), .o(n_4639) );
na02f80 g757839 ( .a(n_22983), .b(n_22981), .o(n_22982) );
in01f80 g746929 ( .a(n_32915), .o(n_32972) );
ao12f80 g756887 ( .a(n_23743), .b(n_23909), .c(n_23901), .o(n_23910) );
in01f80 g741461 ( .a(n_38794), .o(n_38795) );
ao12f80 g750349 ( .a(n_29670), .b(n_29687), .c(n_29669), .o(n_31164) );
in01f80 FE_OCPC1500_n_26125 ( .a(FE_OCPN1499_n_26125), .o(FE_OCPN1500_n_26125) );
in01f80 g761131 ( .a(n_19219), .o(n_19203) );
no02f80 g772414 ( .a(n_8516), .b(n_8437), .o(n_8626) );
na02f80 g744906 ( .a(n_34883), .b(n_34864), .o(n_34960) );
no02f80 g746625 ( .a(n_34612), .b(n_34667), .o(n_34808) );
in01f80 g751027 ( .a(n_28891), .o(n_28892) );
in01f80 g755676 ( .a(n_24534), .o(n_24601) );
in01f80 newInst_66 ( .a(newNet_65), .o(newNet_66) );
in01f80 FE_RC_2331_0 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_3_), .o(FE_RN_890_0) );
in01f80 FE_RC_2014_0 ( .a(n_13419), .o(FE_RN_665_0) );
in01f80 newInst_3539 ( .a(newNet_3538), .o(newNet_3539) );
na02f80 g742733 ( .a(n_37353), .b(n_37207), .o(n_37397) );
in01f80 g778423 ( .a(n_2731), .o(n_3483) );
in01f80 g763196 ( .a(n_17434), .o(n_17435) );
in01f80 newInst_776 ( .a(newNet_775), .o(newNet_776) );
oa12f80 g773986 ( .a(n_6824), .b(n_6885), .c(n_6945), .o(n_6984) );
na02f80 g741877 ( .a(n_38380), .b(n_38379), .o(n_38381) );
no02f80 g763860 ( .a(n_16682), .b(n_16600), .o(n_16683) );
in01f80 FE_OCP_RBC2577_n_47017 ( .a(n_47017), .o(FE_OCP_RBN2577_n_47017) );
oa12f80 g775524 ( .a(n_5595), .b(n_5594), .c(n_5593), .o(n_5664) );
no02f80 g753477 ( .a(n_26783), .b(n_26748), .o(n_26806) );
in01f80 g763097 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_17508) );
in01f80 g765507 ( .a(n_15837), .o(n_15745) );
in01f80 FE_OCPC3755_n_1451 ( .a(FE_OCPN3754_n_1451), .o(FE_OCPN3755_n_1451) );
na02f80 g745019 ( .a(n_34795), .b(FE_OCP_RBN2451_n_34278), .o(n_34797) );
in01f80 newInst_3611 ( .a(newNet_3610), .o(newNet_3611) );
in01f80 g743691 ( .a(n_36424), .o(n_36425) );
no02f80 g746634 ( .a(n_34473), .b(n_33972), .o(n_34867) );
na02f80 g756082 ( .a(n_24248), .b(n_23762), .o(n_24285) );
no03m80 g743396 ( .a(n_37730), .b(n_37725), .c(n_37632), .o(n_37773) );
no02f80 g781100 ( .a(n_245), .b(n_74), .o(n_252) );
in01f80 g748873 ( .a(n_32420), .o(n_32421) );
in01f80 FE_RC_3894_0 ( .a(n_23995), .o(FE_RN_1690_0) );
oa22f80 g784369 ( .a(FE_OFN774_n_46137), .b(n_6217), .c(FE_OFN805_n_46196), .d(n_6243), .o(n_46175) );
no02f80 g744829 ( .a(n_35035), .b(n_35061), .o(n_35154) );
no02f80 g745607 ( .a(n_34286), .b(n_34314), .o(n_34816) );
in01f80 g765791 ( .a(n_15003), .o(n_15004) );
no02f80 g739088 ( .a(n_41083), .b(n_40826), .o(n_41081) );
in01f80 g757954 ( .a(n_22882), .o(n_22883) );
oa12f80 g773116 ( .a(n_8036), .b(n_8232), .c(n_8062), .o(n_8931) );
na02f80 g744129 ( .a(n_36136), .b(n_36242), .o(n_36260) );
in01f80 g779057 ( .a(n_2118), .o(n_2110) );
ao22s80 g771914 ( .a(n_8875), .b(FE_OCP_RBN3537_n_8597), .c(n_44570), .d(n_8597), .o(n_8980) );
in01f80 g747680 ( .a(n_32223), .o(n_32190) );
in01f80 g766961 ( .a(n_13633), .o(n_13594) );
no02f80 g741009 ( .a(n_39234), .b(n_39278), .o(n_39279) );
na02f80 g770329 ( .a(n_10650), .b(n_10640), .o(n_10641) );
no02f80 g754360 ( .a(n_25777), .b(n_25822), .o(n_25823) );
in01f80 g778203 ( .a(n_2830), .o(n_2831) );
no02f80 g760933 ( .a(n_19417), .b(n_18912), .o(n_19459) );
in01f80 g766609 ( .a(n_14140), .o(n_14141) );
in01f80 newInst_2048 ( .a(newNet_986), .o(newNet_2048) );
in01f80 newInst_2666 ( .a(newNet_2665), .o(newNet_2666) );
in01f80 g775433 ( .a(n_5417), .o(n_5436) );
na02f80 g775133 ( .a(n_5870), .b(n_5868), .o(n_5904) );
no02f80 g763744 ( .a(n_16684), .b(FE_OCP_RBN3061_FE_RN_640_0), .o(n_16733) );
no02f80 g742459 ( .a(n_37609), .b(n_37608), .o(n_37610) );
ao12f80 g763762 ( .a(n_17310), .b(n_17423), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_21_), .o(n_17704) );
na02f80 FE_RC_2803_0 ( .a(FE_RN_1199_0), .b(FE_OCP_RBN2635_n_38806), .o(n_38886) );
in01f80 newInst_1676 ( .a(newNet_11), .o(newNet_1676) );
oa12f80 g755833 ( .a(n_25188), .b(n_25216), .c(n_24813), .o(n_25219) );
no02f80 g772804 ( .a(n_8056), .b(n_8092), .o(n_8199) );
in01f80 newInst_2237 ( .a(newNet_2236), .o(newNet_2237) );
oa12f80 g746569 ( .a(n_34694), .b(n_34666), .c(n_34696), .o(n_35320) );
no02f80 g755778 ( .a(n_24272), .b(n_24295), .o(n_24372) );
in01f80 g775028 ( .a(n_6083), .o(n_6118) );
in01f80 g745432 ( .a(n_35581), .o(n_35582) );
in01f80 FE_OCP_RBC2624_n_3848 ( .a(n_3848), .o(FE_OCP_RBN2624_n_3848) );
in01f80 g752921 ( .a(n_27992), .o(n_27950) );
ao12f80 g737377 ( .a(n_42559), .b(n_42796), .c(n_42581), .o(n_42813) );
ao12f80 g743354 ( .a(n_37803), .b(n_37830), .c(n_46232), .o(n_37857) );
oa12f80 g750972 ( .a(n_30005), .b(FE_OCP_RBN2631_n_29947), .c(n_30003), .o(n_30102) );
no02f80 g780465 ( .a(FE_OFN759_n_45813), .b(FE_OFN50_n_1045), .o(n_821) );
na03f80 FE_RC_724_0 ( .a(n_23246), .b(n_22984), .c(n_23326), .o(n_23327) );
ao12f80 g752771 ( .a(n_27923), .b(n_28132), .c(n_27721), .o(n_28152) );
no02f80 g754227 ( .a(n_25912), .b(FE_OCPN1748_n_23354), .o(n_26002) );
na02f80 g748590 ( .a(n_31584), .b(n_31583), .o(n_31697) );
no02f80 FE_RC_2879_0 ( .a(FE_RN_1243_0), .b(n_14323), .o(FE_RN_1244_0) );
in01f80 g762878 ( .a(n_17866), .o(n_17867) );
na02f80 g765086 ( .a(n_15976), .b(n_15923), .o(n_15977) );
no02f80 g758305 ( .a(FE_OCPN992_n_22249), .b(n_20979), .o(n_22434) );
no02f80 g740549 ( .a(n_39691), .b(n_45738), .o(n_39709) );
in01f80 fopt782911 ( .a(n_27688), .o(n_44360) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_18_ ( .ck(newNet_3427), .d(n_27665), .o(delay_add_ln22_unr17_stage7_stallmux_q_18_) );
na02f80 g750712 ( .a(n_29235), .b(n_29269), .o(n_29376) );
in01f80 g775518 ( .a(n_5711), .o(n_5741) );
na02f80 g751888 ( .a(n_29045), .b(n_28940), .o(n_29650) );
no02f80 g744034 ( .a(n_44223), .b(FE_OCP_DRV_N1598_n_35644), .o(n_35669) );
no02f80 g752612 ( .a(n_28245), .b(n_28244), .o(n_28246) );
no02f80 g768841 ( .a(FE_OCPN867_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_13_), .o(n_12402) );
in01f80 newInst_3619 ( .a(newNet_3618), .o(newNet_3619) );
ao12f80 g784688 ( .a(n_3412), .b(n_3401), .c(n_2695), .o(n_47018) );
no02f80 g774027 ( .a(n_6840), .b(n_6791), .o(n_6918) );
na02f80 g749035 ( .a(n_30945), .b(n_30944), .o(n_30946) );
in01f80 newInst_3452 ( .a(newNet_3451), .o(newNet_3452) );
in01f80 g781216 ( .a(n_160), .o(n_161) );
na02f80 g747110 ( .a(n_33998), .b(n_33624), .o(n_34019) );
na02f80 FE_RC_2025_0 ( .a(FE_RN_672_0), .b(n_14177), .o(FE_RN_673_0) );
no02f80 g775947 ( .a(n_5144), .b(n_4504), .o(n_5193) );
in01f80 g738010 ( .a(n_42175), .o(n_42176) );
na02f80 g747785 ( .a(n_32188), .b(n_31971), .o(n_32260) );
oa12f80 g765230 ( .a(n_15664), .b(n_15928), .c(n_15360), .o(n_15971) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_3_ ( .ck(newNet_2618), .d(n_21124), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_) );
no02f80 g741857 ( .a(n_38262), .b(n_38261), .o(n_38263) );
ao12f80 g748782 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .b(n_32495), .c(n_31887), .o(n_32496) );
in01f80 g773920 ( .a(n_7007), .o(n_6996) );
in01f80 g739783 ( .a(n_40495), .o(n_40513) );
oa22f80 g749476 ( .a(n_31909), .b(n_31319), .c(n_31910), .d(n_31320), .o(n_31976) );
na02f80 g773177 ( .a(n_7802), .b(n_7915), .o(n_7963) );
oa22f80 g779854 ( .a(n_44659), .b(n_1217), .c(n_44637), .d(n_1216), .o(n_1336) );
in01f80 FE_RC_2624_0 ( .a(FE_RN_1093_0), .o(FE_OCPN986_n_28402) );
in01f80 newInst_2153 ( .a(newNet_2152), .o(newNet_2153) );
in01f80 newInst_3506 ( .a(newNet_3505), .o(newNet_3506) );
in01f80 g764975 ( .a(n_16066), .o(n_16026) );
in01f80 FE_OCP_DRV_C1559_n_34288 ( .a(n_34288), .o(FE_OCP_DRV_N1559_n_34288) );
in01f80 g751173 ( .a(n_30126), .o(n_30085) );
in01f80 newInst_1599 ( .a(newNet_1598), .o(newNet_1599) );
na02f80 g745763 ( .a(n_35406), .b(n_34807), .o(n_35417) );
in01f80 g761482 ( .a(n_19792), .o(n_20113) );
no02f80 g753433 ( .a(n_46422), .b(n_26871), .o(n_26988) );
na02f80 g753953 ( .a(n_26195), .b(n_23466), .o(n_26319) );
na02f80 g746505 ( .a(n_33207), .b(n_32918), .o(n_33223) );
na02f80 g767076 ( .a(n_13762), .b(n_13761), .o(n_13763) );
in01f80 newInst_3044 ( .a(newNet_3043), .o(newNet_3044) );
na02f80 g774344 ( .a(n_6507), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6619) );
in01f80 g766072 ( .a(n_14662), .o(n_14687) );
no02f80 g742632 ( .a(n_37413), .b(n_37233), .o(n_37507) );
in01f80 FE_OCP_RBC1712_n_21087 ( .a(n_21087), .o(FE_OCP_RBN1712_n_21087) );
no02f80 g743466 ( .a(n_36607), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36649) );
oa12f80 g738450 ( .a(n_41581), .b(FE_OCPN952_n_41540), .c(n_41629), .o(n_41898) );
in01f80 FE_OCP_RBC2892_n_26152 ( .a(n_26152), .o(FE_OCP_RBN2892_n_26152) );
ao12f80 g745644 ( .a(n_33985), .b(n_34121), .c(n_34041), .o(n_34167) );
in01f80 g772756 ( .a(n_7986), .o(n_8043) );
in01f80 FE_OCP_RBC3557_n_8687 ( .a(n_8687), .o(FE_OCP_RBN3557_n_8687) );
no02f80 g755503 ( .a(n_24539), .b(n_24580), .o(n_24652) );
no02f80 FE_RC_3544_0 ( .a(FE_RN_1535_0), .b(n_18824), .o(n_18858) );
in01f80 g740041 ( .a(n_40018), .o(n_40019) );
in01f80 newInst_1401 ( .a(newNet_1400), .o(newNet_1401) );
no02f80 g738529 ( .a(FE_OCP_RBN2312_n_41420), .b(n_41218), .o(n_41580) );
na02f80 g764379 ( .a(n_16366), .b(n_16365), .o(n_16367) );
no02f80 g737412 ( .a(n_42718), .b(n_42621), .o(n_42740) );
no02f80 g745877 ( .a(n_34052), .b(n_34051), .o(n_34095) );
in01f80 FE_OCP_RBC2921_n_31107 ( .a(n_31107), .o(FE_OCP_RBN2921_n_31107) );
in01f80 FE_OCPC3766_n_14439 ( .a(n_14439), .o(FE_OCPN3766_n_14439) );
na02f80 g744045 ( .a(n_44223), .b(n_35749), .o(n_36295) );
oa12f80 g755235 ( .a(n_24691), .b(n_24970), .c(n_24896), .o(n_25041) );
no02f80 g776701 ( .a(n_4152), .b(n_4025), .o(n_4285) );
no02f80 g754695 ( .a(FE_OCP_RBN3704_n_26231), .b(n_25575), .o(n_26812) );
in01f80 newInst_747 ( .a(newNet_746), .o(newNet_747) );
in01f80 FE_OCP_RBC2777_n_15595 ( .a(n_15595), .o(FE_OCP_RBN2777_n_15595) );
in01f80 FE_RC_3512_0 ( .a(FE_RN_1517_0), .o(FE_OCPN1035_n_28288) );
ao12f80 g745868 ( .a(n_35357), .b(n_35356), .c(n_35355), .o(n_35884) );
no02f80 g752003 ( .a(n_28919), .b(n_28982), .o(n_29000) );
oa12f80 g741903 ( .a(n_38127), .b(n_38126), .c(n_38125), .o(n_38892) );
no02f80 g743997 ( .a(n_35984), .b(n_35950), .o(n_36032) );
na02f80 g743727 ( .a(n_37405), .b(n_46233), .o(n_37359) );
oa12f80 g759609 ( .a(n_20305), .b(FE_OCP_RBN1706_n_20616), .c(FE_OCPN1504_n_47257), .o(n_20686) );
in01f80 g759111 ( .a(n_21491), .o(n_21492) );
in01f80 newInst_2897 ( .a(newNet_2896), .o(newNet_2897) );
no02f80 g770732 ( .a(n_10015), .b(FE_OCP_RBN3601_FE_OCPN1243_n_44460), .o(n_10061) );
in01f80 g753448 ( .a(n_26983), .o(n_26984) );
na02f80 g777742 ( .a(n_3326), .b(n_2839), .o(n_3365) );
oa22f80 FE_RC_3029_0 ( .a(n_40598), .b(n_40577), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_44690), .o(n_40589) );
na02f80 g755757 ( .a(n_24462), .b(n_24339), .o(n_24520) );
na02f80 FE_RC_86_0 ( .a(FE_RN_24_0), .b(FE_RN_25_0), .o(FE_RN_26_0) );
na02f80 g755623 ( .a(n_24521), .b(n_24421), .o(n_24597) );
na03f80 FE_RC_3236_0 ( .a(n_9421), .b(n_9465), .c(n_9504), .o(n_9627) );
na03f80 FE_RC_2391_0 ( .a(n_42395), .b(n_42397), .c(n_42451), .o(FE_RN_938_0) );
oa12f80 g781079 ( .a(n_256), .b(n_255), .c(n_254), .o(n_443) );
na02f80 g761259 ( .a(n_19055), .b(n_17815), .o(n_19057) );
in01f80 fopt782725 ( .a(n_44101), .o(n_44133) );
in01f80 g770988 ( .a(n_9550), .o(n_9551) );
na02f80 g751717 ( .a(n_29132), .b(n_29028), .o(n_29205) );
oa12f80 g768476 ( .a(n_12384), .b(n_12338), .c(FE_OCPN1002_n_45660), .o(n_12674) );
in01f80 g747086 ( .a(n_32985), .o(n_32986) );
no02f80 g774160 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_19_), .o(n_7143) );
no02f80 g749525 ( .a(n_30409), .b(n_30116), .o(n_30411) );
na02f80 g753668 ( .a(n_26504), .b(n_26424), .o(n_26539) );
oa12f80 g738252 ( .a(n_41920), .b(n_41919), .c(n_41918), .o(n_41982) );
ao12f80 g751510 ( .a(n_28723), .b(FE_OCP_RBN3404_n_28597), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n_28764) );
in01f80 g737904 ( .a(n_42193), .o(n_42221) );
oa22f80 g758640 ( .a(n_22396), .b(n_21695), .c(n_22428), .d(n_21696), .o(n_22522) );
no02f80 g748730 ( .a(n_31113), .b(n_31087), .o(n_31207) );
na02f80 g780109 ( .a(n_45818), .b(n_1208), .o(n_1210) );
in01f80 FE_OCP_RBC3526_n_29624 ( .a(n_29624), .o(FE_OCP_RBN3526_n_29624) );
in01f80 newInst_2117 ( .a(newNet_2116), .o(newNet_2117) );
in01f80 g758015 ( .a(n_22385), .o(n_22386) );
in01f80 newInst_2815 ( .a(newNet_232), .o(newNet_2815) );
no02f80 g775127 ( .a(n_5790), .b(n_4875), .o(n_5885) );
in01f80 g770392 ( .a(n_10612), .o(n_10663) );
no02f80 g758755 ( .a(n_21805), .b(n_21490), .o(n_21872) );
no02f80 g775916 ( .a(n_4936), .b(FE_OCP_RBN2722_n_4219), .o(n_5051) );
no02f80 g770625 ( .a(n_10254), .b(n_10311), .o(n_10407) );
in01f80 g751518 ( .a(n_28822), .o(n_28823) );
in01f80 FE_OCPC1246_n_43120 ( .a(FE_OCPN1245_n_43120), .o(FE_OCPN1246_n_43120) );
in01f80 g779414 ( .a(n_1509), .o(n_1510) );
oa12f80 g757065 ( .a(n_23700), .b(n_23800), .c(n_23698), .o(n_24110) );
in01f80 g779498 ( .a(n_1448), .o(n_1449) );
na02f80 g740992 ( .a(n_39141), .b(n_39156), .o(n_39211) );
na02f80 g749027 ( .a(n_31029), .b(n_27246), .o(n_31030) );
oa22f80 g753315 ( .a(n_27626), .b(n_26935), .c(n_27657), .d(n_26936), .o(n_27676) );
in01f80 newInst_1610 ( .a(newNet_1609), .o(newNet_1610) );
na02f80 g738359 ( .a(n_41751), .b(n_41745), .o(n_41752) );
in01f80 g740278 ( .a(n_40363), .o(n_40364) );
in01f80 FE_OFC835_n_4333 ( .a(n_4333), .o(FE_OFN835_n_4333) );
oa12f80 g736320 ( .a(n_332), .b(n_43823), .c(FE_OFN3_n_43918), .o(n_43873) );
oa12f80 g751209 ( .a(n_29770), .b(n_29783), .c(n_29769), .o(n_30165) );
na02f80 FE_RC_4222_0 ( .a(FE_RN_1847_0), .b(FE_RN_1850_0), .o(FE_RN_1851_0) );
in01f80 FE_OCPC1470_n_23818 ( .a(FE_OCPN1469_n_23818), .o(FE_OCPN1470_n_23818) );
na02f80 g752047 ( .a(n_28729), .b(n_28728), .o(n_28730) );
no02f80 g742406 ( .a(n_37743), .b(n_37723), .o(n_37801) );
in01f80 g779809 ( .a(n_2124), .o(n_2125) );
no02f80 g738059 ( .a(n_42091), .b(n_41907), .o(n_42111) );
in01f80 g742645 ( .a(n_37461), .o(n_37462) );
ao22s80 g736302 ( .a(n_43830), .b(n_43617), .c(n_43829), .d(n_43618), .o(n_43864) );
na02f80 g750948 ( .a(n_28971), .b(n_28970), .o(n_28972) );
in01f80 g780570 ( .a(n_818), .o(n_776) );
in01f80 newInst_3593 ( .a(newNet_3592), .o(newNet_3593) );
no02f80 FE_RC_941_0 ( .a(FE_RN_277_0), .b(FE_RN_276_0), .o(FE_RN_278_0) );
oa22f80 g779888 ( .a(n_44652), .b(n_1009), .c(n_44623), .d(FE_OCPN1394_n_962), .o(n_1308) );
in01f80 g770506 ( .a(n_10365), .o(n_10366) );
na02f80 g743789 ( .a(n_37283), .b(n_37259), .o(n_37260) );
no02f80 g781103 ( .a(n_244), .b(n_94), .o(n_245) );
no02f80 g740159 ( .a(n_39812), .b(n_39900), .o(n_40015) );
in01f80 g744669 ( .a(n_35324), .o(n_35325) );
no02f80 g740452 ( .a(n_39769), .b(n_39768), .o(n_39776) );
in01f80 g771527 ( .a(n_9521), .o(n_9522) );
in01f80 g752479 ( .a(n_27772), .o(n_27745) );
oa22f80 g784367 ( .a(FE_OFN86_n_46137), .b(n_6004), .c(FE_OFN805_n_46196), .d(n_46997), .o(n_46173) );
no02f80 g755112 ( .a(n_25201), .b(FE_OCP_RBN1131_n_24179), .o(n_25291) );
na02f80 g754153 ( .a(n_25982), .b(FE_OCPN1514_FE_OFN738_n_22641), .o(n_26100) );
in01f80 g750826 ( .a(n_29258), .o(n_29230) );
in01f80 g776928 ( .a(n_4072), .o(n_4171) );
in01f80 FE_OCP_RBC2407_n_8242 ( .a(FE_OCP_RBN2406_n_8242), .o(FE_OCP_RBN2407_n_8242) );
in01f80 g752460 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_21_), .o(n_28523) );
oa12f80 g771105 ( .a(n_9886), .b(n_9885), .c(n_9921), .o(n_9958) );
in01f80 FE_RC_461_0 ( .a(n_23462), .o(FE_RN_133_0) );
na02f80 g767887 ( .a(n_12843), .b(n_12759), .o(n_12844) );
in01f80 newInst_2559 ( .a(newNet_2558), .o(newNet_2559) );
na02f80 g776361 ( .a(n_4661), .b(n_4172), .o(n_4771) );
in01f80 newInst_1647 ( .a(newNet_1646), .o(newNet_1647) );
in01f80 g752516 ( .a(n_27727), .o(n_27705) );
na02f80 g770370 ( .a(n_10564), .b(n_44490), .o(n_10614) );
oa12f80 g784070 ( .a(n_1002), .b(n_851), .c(n_45808), .o(n_45816) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_18_ ( .ck(newNet_1415), .d(n_36640), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_) );
in01f80 g777655 ( .a(n_3623), .o(n_3624) );
in01f80 newInst_3731 ( .a(newNet_3730), .o(newNet_3731) );
in01f80 g774484 ( .a(n_6667), .o(n_6625) );
no02f80 FE_RC_1283_0 ( .a(FE_RN_378_0), .b(FE_RN_379_0), .o(FE_RN_380_0) );
in01f80 newInst_2703 ( .a(newNet_2702), .o(newNet_2703) );
na02f80 g775187 ( .a(n_5750), .b(n_4675), .o(n_5766) );
na02f80 g771233 ( .a(n_9791), .b(n_9790), .o(n_9838) );
na02f80 g784120 ( .a(n_45873), .b(n_45866), .o(n_45871) );
ao22s80 g737185 ( .a(n_42934), .b(n_42622), .c(n_42933), .d(n_42623), .o(n_42989) );
na02f80 g743321 ( .a(n_36712), .b(n_36695), .o(n_36737) );
in01f80 g780437 ( .a(n_1068), .o(n_1118) );
oa22f80 FE_RC_3898_0 ( .a(n_24461), .b(n_24719), .c(n_24486), .d(n_24681), .o(n_24826) );
na02f80 g742597 ( .a(n_37505), .b(n_37504), .o(n_37716) );
in01f80 g763848 ( .a(n_16751), .o(n_16727) );
na02f80 g741023 ( .a(n_38834), .b(n_38864), .o(n_38865) );
in01f80 FE_OCP_RBC2423_n_24501 ( .a(n_24501), .o(FE_OCP_RBN2423_n_24501) );
na02f80 g738554 ( .a(n_41446), .b(n_41382), .o(n_41541) );
oa12f80 g754500 ( .a(n_25516), .b(n_25515), .c(n_25514), .o(n_25595) );
no02f80 g756538 ( .a(n_23563), .b(n_23562), .o(n_23613) );
oa12f80 g762840 ( .a(n_17672), .b(n_17771), .c(n_17622), .o(n_17846) );
na03f80 g742690 ( .a(n_37375), .b(n_37380), .c(n_36962), .o(n_37376) );
in01f80 newInst_2833 ( .a(newNet_200), .o(newNet_2833) );
in01f80 newInst_677 ( .a(newNet_676), .o(newNet_677) );
in01f80 g766240 ( .a(n_14444), .o(n_14443) );
oa22f80 FE_RC_30_0 ( .a(FE_OFN84_n_46137), .b(n_6477), .c(FE_OFN806_n_46196), .d(FE_OCP_RBN3141_n_6477), .o(n_46182) );
na02f80 FE_RC_754_0 ( .a(FE_RN_234_0), .b(FE_RN_235_0), .o(FE_RN_236_0) );
na02f80 g746896 ( .a(FE_OCP_RBN3384_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_26_), .o(n_33305) );
no02f80 g762140 ( .a(n_18771), .b(n_18818), .o(n_18843) );
ao12f80 g760851 ( .a(n_19382), .b(n_19514), .c(n_19422), .o(n_19602) );
na02f80 FE_RC_2344_0 ( .a(FE_RN_898_0), .b(n_19097), .o(n_19125) );
na02f80 g765103 ( .a(n_15931), .b(n_16023), .o(n_16103) );
in01f80 g751613 ( .a(n_28761), .o(n_28762) );
na02f80 g765209 ( .a(n_15405), .b(n_15403), .o(n_15487) );
oa12f80 g739138 ( .a(n_41013), .b(n_40992), .c(n_40981), .o(n_41044) );
in01f80 newInst_3131 ( .a(newNet_2604), .o(newNet_3131) );
na02f80 FE_RC_1065_0 ( .a(FE_RN_312_0), .b(FE_RN_313_0), .o(FE_RN_314_0) );
na02f80 g780886 ( .a(n_377), .b(n_393), .o(n_400) );
in01f80 FE_OCP_RBC3139_n_40568 ( .a(n_40568), .o(FE_OCP_RBN3139_n_40568) );
in01f80 newInst_586 ( .a(newNet_585), .o(newNet_586) );
ao12f80 g772841 ( .a(n_8068), .b(n_8067), .c(n_8066), .o(n_9640) );
na02f80 g759364 ( .a(n_21207), .b(n_21206), .o(n_21208) );
no02f80 g742374 ( .a(n_37797), .b(n_37796), .o(n_37798) );
na02f80 g760423 ( .a(FE_OCP_RBN1718_n_20090), .b(n_20144), .o(n_20162) );
in01f80 newInst_607 ( .a(newNet_395), .o(newNet_607) );
no02f80 g780315 ( .a(n_995), .b(n_1061), .o(n_991) );
no02f80 g770124 ( .a(n_10804), .b(n_10691), .o(n_10904) );
na02f80 g778171 ( .a(n_2859), .b(n_2858), .o(n_2963) );
no02f80 g773249 ( .a(n_7579), .b(n_7578), .o(n_7580) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_12_ ( .ck(newNet_367), .d(n_1337), .o(delay_xor_ln22_unr3_stage2_stallmux_q_12_) );
no02f80 g777834 ( .a(n_3330), .b(n_3302), .o(n_3391) );
ao22s80 g757629 ( .a(FE_OCP_RBN1195_n_22542), .b(n_22309), .c(n_45497), .d(n_22272), .o(n_22710) );
no02f80 g770772 ( .a(n_10178), .b(n_10216), .o(n_10375) );
in01f80 FE_OCP_RBC2944_FE_RN_1269_0 ( .a(FE_RN_1269_0), .o(FE_OCP_RBN2944_FE_RN_1269_0) );
in01f80 g738487 ( .a(n_41588), .o(n_41589) );
in01f80 g740201 ( .a(n_39824), .o(n_39784) );
oa12f80 g751298 ( .a(n_29639), .b(n_29638), .c(n_29637), .o(n_30083) );
na02f80 g753899 ( .a(n_26227), .b(n_26157), .o(n_26368) );
in01f80 g773925 ( .a(n_7294), .o(n_7295) );
in01f80 g736682 ( .a(n_43094), .o(n_43116) );
na02f80 g738706 ( .a(n_41456), .b(n_41462), .o(n_41488) );
in01f80 newInst_479 ( .a(newNet_478), .o(newNet_479) );
no02f80 g758732 ( .a(n_21872), .b(FE_OCP_RBN2951_n_21489), .o(n_21927) );
in01f80 g771878 ( .a(n_8929), .o(n_8930) );
na02f80 g755053 ( .a(n_25503), .b(n_25502), .o(n_25537) );
na02f80 g772916 ( .a(n_7750), .b(n_7365), .o(n_7804) );
na02f80 g760204 ( .a(FE_OCP_RBN1332_n_20249), .b(n_19641), .o(n_20334) );
in01f80 g762377 ( .a(n_18528), .o(n_18623) );
na02f80 g749663 ( .a(n_30149), .b(n_29968), .o(n_30178) );
no02f80 g746882 ( .a(FE_OCP_RBN3387_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_29_), .o(n_33338) );
in01f80 g749867 ( .a(n_31312), .o(n_31368) );
in01f80 g752735 ( .a(n_27994), .o(n_27995) );
na02f80 g766795 ( .a(n_14526), .b(n_14525), .o(n_14527) );
in01f80 FE_OCP_RBC3210_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3210_n_44365) );
oa22f80 FE_RC_1689_0 ( .a(FE_OFN802_n_46285), .b(n_12196), .c(FE_OFN771_n_46337), .d(n_44766), .o(n_46347) );
in01f80 newInst_1680 ( .a(newNet_150), .o(newNet_1680) );
no02f80 g769028 ( .a(n_11633), .b(n_11738), .o(n_11758) );
ao12f80 g738218 ( .a(n_41958), .b(n_41924), .c(n_41957), .o(n_42065) );
in01f80 g763057 ( .a(n_17641), .o(n_17642) );
oa22f80 g769986 ( .a(n_10972), .b(n_10157), .c(n_11057), .d(n_10156), .o(n_11068) );
in01f80 g758550 ( .a(n_22249), .o(n_22288) );
na02f80 g745631 ( .a(n_34289), .b(FE_OCP_DRV_N1560_n_34288), .o(n_34310) );
na02f80 g748303 ( .a(n_31477), .b(FE_OCPN1418_n_31504), .o(n_31505) );
no02f80 g754856 ( .a(n_25673), .b(n_25672), .o(n_25695) );
in01f80 newInst_235 ( .a(newNet_234), .o(newNet_235) );
na02f80 g774304 ( .a(FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_1_), .o(n_6525) );
in01f80 g746752 ( .a(n_33037), .o(n_33038) );
in01f80 newInst_1800 ( .a(newNet_1629), .o(newNet_1800) );
no02f80 g746319 ( .a(n_33523), .b(n_33544), .o(n_33589) );
in01f80 g754712 ( .a(n_26550), .o(n_26508) );
oa22f80 FE_RC_3024_0 ( .a(n_40277), .b(n_40515), .c(n_40278), .d(n_40516), .o(n_40552) );
na02f80 g763447 ( .a(n_17032), .b(n_17164), .o(n_17321) );
in01f80 newInst_2919 ( .a(newNet_2918), .o(newNet_2919) );
in01f80 g749645 ( .a(n_30250), .o(n_30204) );
in01f80 g780897 ( .a(n_442), .o(n_460) );
no02f80 g760907 ( .a(n_19284), .b(n_18505), .o(n_19365) );
in01f80 g757396 ( .a(n_23122), .o(n_23123) );
no02f80 g769223 ( .a(FE_OCP_RBN3092_n_11475), .b(n_11502), .o(n_11608) );
oa22f80 g778755 ( .a(n_2169), .b(n_1505), .c(n_2200), .d(n_1504), .o(n_2752) );
no02f80 g760871 ( .a(n_19467), .b(n_18010), .o(n_19533) );
in01f80 newInst_1095 ( .a(newNet_982), .o(newNet_1095) );
in01f80 FE_OCP_RBC3006_n_11087 ( .a(n_11087), .o(FE_OCP_RBN3006_n_11087) );
in01f80 g777342 ( .a(n_5005), .o(n_5006) );
na02f80 g766944 ( .a(n_14211), .b(n_14209), .o(n_14299) );
no02f80 g738680 ( .a(n_41564), .b(n_41562), .o(n_41604) );
ao12f80 g748947 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_), .o(n_32502) );
in01f80 g741494 ( .a(n_38772), .o(n_38773) );
in01f80 g740075 ( .a(n_40137), .o(n_40138) );
na02f80 g751386 ( .a(FE_OCP_RBN3396_n_28651), .b(n_28579), .o(n_28745) );
no02f80 g739201 ( .a(n_40679), .b(n_45180), .o(n_40746) );
no02f80 g740601 ( .a(n_39558), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39594) );
na02f80 g753881 ( .a(n_27033), .b(n_26884), .o(n_27054) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_3_ ( .ck(newNet_2522), .d(n_26582), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_) );
no02f80 g769346 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_10_), .o(n_11738) );
na02f80 g750118 ( .a(FE_OCP_RBN2571_n_29922), .b(n_45760), .o(n_30349) );
no02f80 g773549 ( .a(n_45864), .b(n_7481), .o(n_7483) );
na02f80 g759189 ( .a(n_21184), .b(n_21183), .o(n_21185) );
in01f80 g775343 ( .a(n_5982), .o(n_5916) );
in01f80 g747179 ( .a(n_32719), .o(n_32720) );
na02f80 g745187 ( .a(n_34595), .b(n_34762), .o(n_34782) );
in01f80 newInst_1313 ( .a(newNet_1020), .o(newNet_1313) );
oa22f80 FE_RC_104_0 ( .a(n_18632), .b(n_19470), .c(n_18631), .d(n_19471), .o(n_19601) );
na02f80 g739704 ( .a(n_40502), .b(n_40371), .o(n_40531) );
oa22f80 g743813 ( .a(n_35876), .b(n_36262), .c(n_35877), .d(n_36263), .o(n_36337) );
in01f80 FE_OCP_RBC2211_n_37720 ( .a(n_37720), .o(FE_OCP_RBN2211_n_37720) );
in01f80 g744585 ( .a(n_36664), .o(n_36665) );
na02f80 g748908 ( .a(n_32393), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .o(n_32497) );
in01f80 newInst_2268 ( .a(newNet_297), .o(newNet_2268) );
no02f80 g778420 ( .a(n_2672), .b(delay_add_ln22_unr2_stage2_stallmux_q_26_), .o(n_2728) );
in01f80 g776665 ( .a(n_4305), .o(n_4306) );
in01f80 g778924 ( .a(n_2166), .o(n_2167) );
in01f80 g758495 ( .a(FE_OFN735_n_22641), .o(n_22725) );
no02f80 g756452 ( .a(n_23854), .b(n_23853), .o(n_23855) );
in01f80 FE_OCP_DRV_C1564_n_19665 ( .a(FE_OCP_DRV_N1563_n_19665), .o(FE_OCP_DRV_N1564_n_19665) );
no02f80 g740029 ( .a(n_40038), .b(n_40004), .o(n_40080) );
no02f80 g742306 ( .a(n_37837), .b(n_37836), .o(n_37881) );
no02f80 g738915 ( .a(n_41223), .b(n_40983), .o(n_41251) );
in01f80 g778180 ( .a(n_2805), .o(n_2789) );
ao12f80 g778189 ( .a(n_2808), .b(n_2871), .c(n_2870), .o(n_3089) );
na02f80 g743280 ( .a(n_36767), .b(n_36732), .o(n_36789) );
no02f80 g771612 ( .a(n_10340), .b(n_10283), .o(n_10383) );
in01f80 g742045 ( .a(n_38088), .o(n_38051) );
no02f80 g759648 ( .a(n_21629), .b(n_21563), .o(n_21698) );
na02f80 g773786 ( .a(n_7147), .b(n_7146), .o(n_7157) );
no02f80 g757082 ( .a(n_23177), .b(n_21785), .o(n_23250) );
oa12f80 g762004 ( .a(n_18355), .b(n_18593), .c(delay_add_ln22_unr11_stage5_stallmux_q_29_), .o(n_18634) );
na02f80 g769865 ( .a(n_11026), .b(n_11000), .o(n_11062) );
no02f80 g771603 ( .a(n_44056), .b(n_9236), .o(n_9333) );
no02f80 FE_RC_604_0 ( .a(FE_RN_189_0), .b(FE_RN_190_0), .o(FE_RN_191_0) );
in01f80 fopt782892 ( .a(n_17759), .o(n_44334) );
ao22s80 g754800 ( .a(n_25952), .b(n_25709), .c(n_25953), .d(n_25708), .o(n_26643) );
no02f80 g768332 ( .a(n_12490), .b(n_12370), .o(n_12516) );
no02f80 g771206 ( .a(FE_OCP_RBN2589_n_9492), .b(n_9552), .o(n_9476) );
no02f80 g773486 ( .a(n_7526), .b(n_7497), .o(n_7562) );
no02f80 g753926 ( .a(n_26223), .b(n_26191), .o(n_26373) );
oa12f80 g774394 ( .a(n_6854), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_14_), .o(n_7302) );
no02f80 g762737 ( .a(n_17826), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_), .o(n_17849) );
no02f80 g748176 ( .a(n_31929), .b(n_32054), .o(n_32130) );
no02f80 g767067 ( .a(n_13765), .b(n_13764), .o(n_13793) );
in01f80 newInst_2471 ( .a(newNet_2470), .o(newNet_2471) );
na02f80 g743352 ( .a(n_36692), .b(n_36659), .o(n_36706) );
in01f80 g756217 ( .a(n_24175), .o(n_24199) );
in01f80 newInst_619 ( .a(newNet_618), .o(newNet_619) );
na02f80 FE_RC_560_0 ( .a(FE_RN_170_0), .b(n_30675), .o(n_46958) );
ao22s80 FE_RC_1502_0 ( .a(n_25488), .b(n_25732), .c(n_25487), .d(FE_OCP_RBN2764_n_25732), .o(n_25817) );
no02f80 g771220 ( .a(FE_OCP_RBN2703_n_9411), .b(FE_OCP_RBN3550_n_44575), .o(n_9491) );
ao12f80 g742932 ( .a(n_37003), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_11_), .o(n_37354) );
no02f80 g765393 ( .a(n_47261), .b(n_15216), .o(n_15371) );
no02f80 g764501 ( .a(n_16182), .b(n_16271), .o(n_16365) );
no02f80 g765787 ( .a(n_14958), .b(FE_OCP_RBN2756_FE_RN_722_0), .o(n_15005) );
no02f80 g768031 ( .a(n_12790), .b(n_12840), .o(n_12885) );
in01f80 g780372 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_6_), .o(n_912) );
in01f80 g748587 ( .a(n_31585), .o(n_31586) );
in01f80 g763906 ( .a(n_17362), .o(n_17301) );
oa22f80 FE_RC_1496_0 ( .a(n_28948), .b(n_28602), .c(n_28949), .d(n_28601), .o(n_29030) );
in01f80 newInst_2792 ( .a(newNet_2791), .o(newNet_2792) );
oa12f80 g749818 ( .a(n_31282), .b(FE_OCP_RBN3010_n_31117), .c(n_31275), .o(n_31615) );
no02f80 g779750 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_14_), .o(n_1673) );
na02f80 g765284 ( .a(n_15922), .b(n_15784), .o(n_15828) );
in01f80 newInst_1913 ( .a(newNet_11), .o(newNet_1913) );
no02f80 g743828 ( .a(n_36071), .b(n_36204), .o(n_36205) );
in01f80 FE_RC_3991_0 ( .a(n_25016), .o(FE_RN_1731_0) );
ao12f80 g748096 ( .a(n_31698), .b(n_31742), .c(n_31756), .o(n_31853) );
oa22f80 FE_RC_3871_0 ( .a(n_27966), .b(FE_OCP_RBN1149_n_27962), .c(n_27962), .d(FE_OCP_RBN1148_n_27966), .o(n_28116) );
na02f80 g745310 ( .a(n_35724), .b(n_35679), .o(n_35767) );
in01f80 g774080 ( .a(n_6760), .o(n_6823) );
in01f80 g740100 ( .a(n_40324), .o(n_40325) );
in01f80 g764055 ( .a(FE_OFN778_n_17093), .o(n_17661) );
in01f80 newInst_459 ( .a(newNet_458), .o(newNet_459) );
na03f80 FE_RC_445_0 ( .a(n_1455), .b(n_1467), .c(n_1398), .o(n_1533) );
in01f80 FE_OCPC1491_n_22036 ( .a(n_22036), .o(FE_OCPN1491_n_22036) );
na02f80 g773047 ( .a(n_7693), .b(n_7626), .o(n_7713) );
na02f80 g760716 ( .a(n_19568), .b(n_19604), .o(n_19730) );
na02f80 g776090 ( .a(n_4716), .b(n_4602), .o(n_4669) );
no02f80 g776427 ( .a(n_4238), .b(n_3082), .o(n_4328) );
no02f80 g759051 ( .a(n_21421), .b(n_21219), .o(n_21540) );
in01f80 FE_OCP_DRV_C1573_n_28869 ( .a(n_28869), .o(FE_OCP_DRV_N1573_n_28869) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_23_ ( .ck(newNet_232), .d(n_46194), .o(delay_xor_ln22_unr6_stage3_stallmux_q_23_) );
in01f80 newInst_3742 ( .a(newNet_2047), .o(newNet_3742) );
na02f80 g770183 ( .a(n_10813), .b(n_10684), .o(n_10900) );
oa22f80 FE_RC_1298_0 ( .a(n_2913), .b(n_3524), .c(n_4905), .d(n_3029), .o(n_3578) );
in01f80 g777941 ( .a(n_3147), .o(n_3119) );
no02f80 g757567 ( .a(n_23277), .b(n_22700), .o(n_23357) );
in01f80 FE_RC_2663_0 ( .a(n_2261), .o(FE_RN_1112_0) );
in01f80 g745335 ( .a(n_35959), .o(n_35960) );
ao12f80 g784134 ( .a(n_45880), .b(n_7659), .c(n_45884), .o(n_45887) );
na02f80 g765929 ( .a(n_14764), .b(FE_OCP_RBN3536_n_13765), .o(n_14817) );
ao12f80 g759374 ( .a(n_21035), .b(n_20967), .c(n_21036), .o(n_21119) );
in01f80 FE_OCPC1501_n_20723 ( .a(n_20723), .o(FE_OCPN1501_n_20723) );
in01f80 g753427 ( .a(n_27037), .o(n_27038) );
in01f80 g762417 ( .a(n_18568), .o(n_18569) );
oa12f80 g768244 ( .a(n_12572), .b(n_12571), .c(n_12570), .o(n_12612) );
na02f80 g753960 ( .a(n_26216), .b(n_26118), .o(n_26189) );
in01f80 g742987 ( .a(n_37016), .o(n_36969) );
in01f80 newInst_48 ( .a(newNet_47), .o(newNet_48) );
oa22f80 g739850 ( .a(n_40343), .b(n_40318), .c(n_40344), .d(n_40319), .o(n_40420) );
in01f80 g764033 ( .a(n_18032), .o(n_18010) );
in01f80 g768995 ( .a(n_11815), .o(n_11816) );
ao12f80 g739178 ( .a(n_40672), .b(n_40801), .c(n_40735), .o(n_40897) );
no02f80 g758888 ( .a(n_21361), .b(FE_OCPN1524_n_45072), .o(n_21508) );
no02f80 g766134 ( .a(n_14484), .b(n_14479), .o(n_14480) );
na02f80 g773083 ( .a(n_7768), .b(n_7830), .o(n_8160) );
na02f80 g742450 ( .a(n_37693), .b(n_37628), .o(n_37720) );
in01f80 g749156 ( .a(FE_OCP_RBN2912_n_30908), .o(n_30955) );
in01f80 g743159 ( .a(n_36922), .o(n_36914) );
no02f80 g778498 ( .a(n_2340), .b(n_2282), .o(n_2419) );
na02f80 g764882 ( .a(n_15684), .b(n_15683), .o(n_15685) );
oa22f80 FE_RC_1194_0 ( .a(n_7726), .b(n_7693), .c(n_7675), .d(n_7725), .o(n_7747) );
na02f80 g763018 ( .a(n_17715), .b(n_17640), .o(n_17737) );
in01f80 g752725 ( .a(n_27997), .o(n_27932) );
oa12f80 g765945 ( .a(n_14656), .b(n_14750), .c(n_14626), .o(n_14772) );
in01f80 FE_OCP_DRV_C3156_n_15342 ( .a(FE_OCP_DRV_N3155_n_15342), .o(FE_OCP_DRV_N3156_n_15342) );
no02f80 g758295 ( .a(n_22288), .b(n_20555), .o(n_22468) );
in01f80 g740840 ( .a(n_39462), .o(n_39463) );
na02f80 g765578 ( .a(n_15132), .b(n_15091), .o(n_15177) );
oa12f80 g763273 ( .a(n_17228), .b(n_17227), .c(n_17226), .o(n_18559) );
in01f80 g756764 ( .a(n_23537), .o(n_23538) );
no02f80 g750475 ( .a(n_29572), .b(n_29571), .o(n_29622) );
in01f80 g736893 ( .a(n_43587), .o(n_43588) );
in01f80 newInst_1772 ( .a(newNet_863), .o(newNet_1772) );
in01f80 g744212 ( .a(n_35971), .o(n_35972) );
ao12f80 g775857 ( .a(n_5195), .b(n_5240), .c(n_5194), .o(n_5286) );
ao12f80 g757697 ( .a(n_23088), .b(n_23090), .c(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_23221) );
no02f80 g757288 ( .a(n_23223), .b(n_23222), .o(n_23224) );
in01f80 newInst_93 ( .a(newNet_92), .o(newNet_93) );
na02f80 g759345 ( .a(n_20890), .b(n_20829), .o(n_20943) );
ao12f80 g746837 ( .a(n_32940), .b(n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_21_), .o(n_33524) );
in01f80 g768393 ( .a(n_12526), .o(n_12527) );
in01f80 g763511 ( .a(n_16943), .o(n_16982) );
in01f80 FE_OCP_RBC2610_n_3718 ( .a(n_3718), .o(FE_OCP_RBN2610_n_3718) );
na02f80 g775906 ( .a(FE_OCP_RBN3685_n_5217), .b(n_4867), .o(n_5318) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_29_ ( .ck(newNet_2075), .d(n_6719), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_11_ ( .ck(newNet_2593), .d(n_27129), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_11_) );
ao12f80 g757366 ( .a(n_22918), .b(n_23400), .c(n_22808), .o(n_23416) );
no02f80 g760469 ( .a(n_20005), .b(n_19921), .o(n_20006) );
no02f80 g755184 ( .a(n_25042), .b(n_24895), .o(n_25043) );
in01f80 g774218 ( .a(n_6855), .o(n_6856) );
oa22f80 FE_RC_3443_0 ( .a(n_36846), .b(n_36723), .c(n_36722), .d(n_36889), .o(n_36890) );
na02f80 FE_RC_2969_0 ( .a(FE_RN_1297_0), .b(n_26153), .o(FE_RN_1298_0) );
ao22s80 g777868 ( .a(n_4211), .b(n_2913), .c(n_3226), .d(n_2759), .o(n_3250) );
in01f80 g745573 ( .a(n_34348), .o(n_34321) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_23_ ( .ck(newNet_3524), .d(n_22774), .o(delay_add_ln22_unr14_stage6_stallmux_q_23_) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_6_ ( .ck(newNet_1566), .d(n_26796), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_6_) );
in01f80 g743405 ( .a(n_36709), .o(n_36654) );
in01f80 g737053 ( .a(n_43202), .o(n_43203) );
oa22f80 g766610 ( .a(n_46984), .b(n_12868), .c(n_14013), .d(n_12846), .o(n_14140) );
na02f80 FE_RC_1838_0 ( .a(n_23212), .b(FE_RN_554_0), .o(FE_RN_555_0) );
ao12f80 g742164 ( .a(n_38003), .b(n_44887), .c(n_37935), .o(n_38443) );
na02f80 g765668 ( .a(n_15067), .b(n_13479), .o(n_15170) );
oa22f80 g784358 ( .a(FE_OFN775_n_46137), .b(n_5795), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5841), .o(n_46164) );
oa12f80 g776135 ( .a(n_4484), .b(n_4454), .c(n_4394), .o(n_4581) );
na02f80 g755585 ( .a(FE_OCP_RBN2396_n_24451), .b(n_22111), .o(n_24512) );
in01f80 FE_OCP_RBC2978_n_5555 ( .a(FE_OCP_RBN2977_n_5555), .o(FE_OCP_RBN2978_n_5555) );
no02f80 g778182 ( .a(n_2742), .b(n_2479), .o(n_2845) );
in01f80 g742617 ( .a(n_37929), .o(n_37967) );
in01f80 g761874 ( .a(n_18936), .o(n_18937) );
in01f80 g743166 ( .a(n_36919), .o(n_36920) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_27_ ( .ck(newNet_2836), .d(n_12145), .o(delay_add_ln22_unr8_stage4_stallmux_q_27_) );
na02f80 g771136 ( .a(n_47259), .b(n_9593), .o(n_9664) );
no02f80 g740682 ( .a(n_39550), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39588) );
na02f80 g750779 ( .a(n_29167), .b(FE_RN_1513_0), .o(n_29168) );
no02f80 g762131 ( .a(n_18188), .b(delay_add_ln22_unr11_stage5_stallmux_q_18_), .o(n_18265) );
no02f80 g777128 ( .a(n_3547), .b(n_3396), .o(n_3572) );
ao12f80 g750293 ( .a(n_30787), .b(n_30786), .c(n_30785), .o(n_31214) );
ao12f80 g763537 ( .a(n_16751), .b(n_16827), .c(n_16726), .o(n_16938) );
na02f80 FE_RC_3136_0 ( .a(FE_RN_1389_0), .b(FE_RN_1390_0), .o(FE_RN_1391_0) );
no02f80 g764918 ( .a(n_15612), .b(n_15611), .o(n_15615) );
na02f80 g755896 ( .a(n_24305), .b(FE_OCP_RBN2307_n_24288), .o(n_24392) );
ms00f80 cos_out_reg_28_ ( .ck(newNet_3705), .d(n_43904), .o(cos_out_28) );
ao12f80 g738609 ( .a(n_41489), .b(n_41716), .c(n_41140), .o(n_41927) );
na02f80 g760878 ( .a(n_19506), .b(n_19514), .o(n_19507) );
na02f80 g779363 ( .a(n_1588), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_), .o(n_1616) );
oa22f80 g739684 ( .a(n_40491), .b(n_40281), .c(n_40492), .d(n_40282), .o(n_40525) );
in01f80 g779663 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n_1369) );
na02f80 g771380 ( .a(FE_OCP_RBN2678_n_9247), .b(FE_OCP_RBN3550_n_44575), .o(n_9344) );
na02f80 g780450 ( .a(n_764), .b(n_580), .o(n_806) );
in01f80 newInst_2515 ( .a(newNet_2514), .o(newNet_2515) );
in01f80 FE_OCP_RBC2716_n_14982 ( .a(FE_OCP_RBN2714_n_14982), .o(FE_OCP_RBN2716_n_14982) );
ao12f80 g751810 ( .a(n_29131), .b(n_29077), .c(n_28919), .o(n_29823) );
na02f80 g778580 ( .a(n_2476), .b(delay_add_ln22_unr2_stage2_stallmux_q_23_), .o(n_2569) );
no02f80 FE_RC_4179_0 ( .a(FE_RN_1825_0), .b(n_33804), .o(FE_RN_1826_0) );
oa22f80 g739273 ( .a(n_45153), .b(n_40756), .c(n_45155), .d(delay_add_ln22_unr27_stage10_stallmux_q_17_), .o(n_41146) );
no02f80 g743007 ( .a(n_37088), .b(n_37108), .o(n_37279) );
oa22f80 FE_RC_338_0 ( .a(n_12017), .b(n_12330), .c(n_12018), .d(n_12352), .o(n_12428) );
in01f80 newInst_1624 ( .a(newNet_1623), .o(newNet_1624) );
na02f80 g753938 ( .a(n_26220), .b(n_26204), .o(n_26225) );
oa22f80 g758180 ( .a(n_21968), .b(n_21916), .c(n_21990), .d(n_21917), .o(n_22044) );
in01f80 FE_OCP_RBC2128_n_6745 ( .a(n_6745), .o(FE_OCP_RBN2128_n_6745) );
in01f80 newInst_3314 ( .a(newNet_3199), .o(newNet_3314) );
in01f80 g779372 ( .a(n_1608), .o(n_1625) );
na02f80 g764441 ( .a(n_16224), .b(n_16202), .o(n_16274) );
no02f80 g776443 ( .a(n_4486), .b(n_3580), .o(n_4689) );
in01f80 g769918 ( .a(n_11000), .o(n_11027) );
in01f80 fopt783335 ( .a(n_37850), .o(n_44869) );
in01f80 FE_OFC778_n_17093 ( .a(FE_OFN776_n_17093), .o(FE_OFN778_n_17093) );
no02f80 g752245 ( .a(n_28219), .b(n_28032), .o(n_28056) );
ao12f80 g756518 ( .a(n_23993), .b(n_23843), .c(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n_24050) );
in01f80 FE_OCP_RBC3569_n_9188 ( .a(n_9188), .o(FE_OCP_RBN3569_n_9188) );
no02f80 g769382 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_12011) );
in01f80 g755557 ( .a(n_24648), .o(n_24649) );
in01f80 g742464 ( .a(n_37690), .o(n_37691) );
in01f80 g768122 ( .a(n_13412), .o(n_12649) );
no02f80 g774458 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_), .o(n_6940) );
no02f80 g747730 ( .a(n_33840), .b(n_33317), .o(n_33885) );
oa22f80 g774941 ( .a(n_6185), .b(n_5386), .c(n_6184), .d(n_5385), .o(n_6229) );
in01f80 g767195 ( .a(n_14588), .o(n_14730) );
na02f80 g770044 ( .a(n_10932), .b(FE_OCP_RBN3004_n_10930), .o(n_10975) );
na02f80 g737247 ( .a(n_42902), .b(n_42818), .o(n_42945) );
na02f80 g750302 ( .a(n_29766), .b(n_29765), .o(n_29807) );
na02f80 g753571 ( .a(n_26700), .b(n_26726), .o(n_26821) );
in01f80 g738238 ( .a(n_41953), .o(n_42272) );
in01f80 FE_OCP_RBC1357_n_30298 ( .a(n_30298), .o(FE_OCP_RBN1357_n_30298) );
no02f80 g773455 ( .a(n_7510), .b(n_6816), .o(n_7529) );
no02f80 g744895 ( .a(n_34980), .b(n_30504), .o(n_35008) );
na02f80 g763509 ( .a(FE_OCP_RBN3081_n_16977), .b(n_16118), .o(n_17170) );
in01f80 g743031 ( .a(n_37153), .o(n_37154) );
in01f80 g773672 ( .a(n_7306), .o(n_7277) );
in01f80 newInst_511 ( .a(newNet_510), .o(newNet_511) );
ao22s80 FE_RC_3714_0 ( .a(n_38735), .b(n_38784), .c(n_38734), .d(n_38769), .o(n_38818) );
no02f80 g749610 ( .a(n_30483), .b(n_29953), .o(n_30285) );
no02f80 g756476 ( .a(n_23712), .b(n_24182), .o(n_23881) );
in01f80 newInst_1441 ( .a(newNet_830), .o(newNet_1441) );
in01f80 g762906 ( .a(n_18102), .o(n_18103) );
no02f80 g760826 ( .a(n_19462), .b(n_19533), .o(n_19534) );
no02f80 g779503 ( .a(n_1435), .b(n_1405), .o(n_1485) );
oa12f80 g755663 ( .a(n_24443), .b(n_24549), .c(n_24494), .o(n_24556) );
in01f80 g740966 ( .a(n_39215), .o(n_39193) );
in01f80 newInst_3652 ( .a(newNet_3651), .o(newNet_3652) );
na02f80 FE_RC_4174_0 ( .a(FE_RN_1820_0), .b(n_33772), .o(n_33827) );
in01f80 newInst_3084 ( .a(newNet_3083), .o(newNet_3084) );
no02f80 g762610 ( .a(n_45524), .b(n_17734), .o(n_18351) );
in01f80 g781396 ( .a(beta_12), .o(n_27) );
no02f80 FE_RC_2437_0 ( .a(FE_RN_970_0), .b(FE_RN_971_0), .o(FE_RN_972_0) );
in01f80 g746322 ( .a(n_33583), .o(n_34313) );
no02f80 FE_RC_2840_0 ( .a(n_13684), .b(n_13637), .o(FE_RN_1221_0) );
na02f80 g748227 ( .a(FE_OCP_RBN3731_n_31819), .b(n_30522), .o(n_32119) );
na02f80 g769962 ( .a(n_10896), .b(n_10895), .o(n_10998) );
no02f80 g772291 ( .a(n_8587), .b(n_8631), .o(n_8732) );
na02f80 g764703 ( .a(n_16450), .b(n_15838), .o(n_16447) );
oa12f80 g760495 ( .a(n_19910), .b(n_20451), .c(n_19872), .o(n_20559) );
ao12f80 g774268 ( .a(n_6370), .b(n_6513), .c(n_6394), .o(n_6555) );
in01f80 g762365 ( .a(n_18839), .o(n_18693) );
in01f80 newInst_2740 ( .a(newNet_2739), .o(newNet_2740) );
na02f80 g753858 ( .a(n_27053), .b(n_27065), .o(n_27094) );
no02f80 g767327 ( .a(n_13508), .b(n_13482), .o(n_13626) );
na03f80 g761706 ( .a(n_19402), .b(n_19404), .c(n_18808), .o(n_19524) );
na02f80 g754303 ( .a(n_25875), .b(n_25503), .o(n_25925) );
in01f80 g753357 ( .a(n_27070), .o(n_27103) );
ao12f80 g751751 ( .a(n_28302), .b(n_28301), .c(n_28300), .o(n_29504) );
in01f80 g770080 ( .a(n_10984), .o(n_10985) );
na02f80 g766926 ( .a(n_14386), .b(n_14292), .o(n_14387) );
na02f80 g780608 ( .a(n_713), .b(n_712), .o(n_725) );
in01f80 g745347 ( .a(n_36159), .o(n_36160) );
na02f80 g767951 ( .a(n_13078), .b(n_13159), .o(n_13166) );
in01f80 g771395 ( .a(n_9213), .o(n_9214) );
in01f80 newInst_2006 ( .a(newNet_538), .o(newNet_2006) );
in01f80 g772370 ( .a(n_8506), .o(n_8507) );
in01f80 g752192 ( .a(n_28112), .o(n_28113) );
no02f80 g748658 ( .a(n_31439), .b(n_31356), .o(n_31440) );
na02f80 g765321 ( .a(n_15135), .b(FE_OCP_RBN2413_n_13960), .o(n_15263) );
na02f80 g740367 ( .a(n_39787), .b(n_39808), .o(n_39859) );
no02f80 g743875 ( .a(n_35987), .b(n_35867), .o(n_36013) );
in01f80 g741091 ( .a(n_39274), .o(n_39275) );
in01f80 g741219 ( .a(n_39297), .o(n_39298) );
na02f80 g751945 ( .a(n_28221), .b(n_28220), .o(n_28247) );
no02f80 g760156 ( .a(n_20565), .b(n_20605), .o(n_20675) );
in01f80 newInst_3170 ( .a(newNet_3151), .o(newNet_3170) );
in01f80 newInst_2432 ( .a(newNet_2399), .o(newNet_2432) );
no02f80 g759643 ( .a(n_20616), .b(n_20338), .o(n_20617) );
ao12f80 g747594 ( .a(n_31706), .b(n_32190), .c(n_31702), .o(n_32242) );
in01f80 newInst_3713 ( .a(newNet_3712), .o(newNet_3713) );
na02f80 g751984 ( .a(n_28781), .b(n_27995), .o(n_28841) );
in01f80 g774898 ( .a(n_6297), .o(n_6254) );
oa12f80 g741951 ( .a(n_37842), .b(n_44036), .c(n_37881), .o(n_38092) );
no02f80 g771128 ( .a(n_9546), .b(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .o(n_9685) );
in01f80 g736666 ( .a(n_43440), .o(n_43475) );
no02f80 g768467 ( .a(n_12419), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_10_), .o(n_12432) );
oa12f80 g760596 ( .a(n_19879), .b(n_19878), .c(n_19877), .o(n_19961) );
oa12f80 g757724 ( .a(n_23156), .b(n_23155), .c(n_23154), .o(n_23699) );
oa22f80 g773697 ( .a(n_7287), .b(n_7155), .c(n_7261), .d(n_7154), .o(n_7354) );
no02f80 FE_RC_3677_0 ( .a(FE_RN_1615_0), .b(n_46969), .o(n_21125) );
no02f80 g763329 ( .a(n_16882), .b(FE_OCP_RBN1210_n_16814), .o(n_16951) );
in01f80 FE_RC_3857_0 ( .a(FE_RN_1684_0), .o(n_21191) );
in01f80 FE_OCPC1230_n_42201 ( .a(n_42201), .o(FE_OCPN1230_n_42201) );
na02f80 g757004 ( .a(n_23592), .b(n_23591), .o(n_23593) );
no02f80 g760117 ( .a(n_20387), .b(FE_OCP_RBN1697_n_19206), .o(n_20539) );
no02f80 g774151 ( .a(n_6872), .b(delay_xor_ln22_unr6_stage3_stallmux_q_20_), .o(n_7168) );
na02f80 g745806 ( .a(n_44100), .b(n_34123), .o(n_34146) );
na02f80 g773251 ( .a(n_8635), .b(n_7593), .o(n_7631) );
in01f80 FE_OCPC932_n_40736 ( .a(FE_OCPN931_n_40736), .o(FE_OCPN932_n_40736) );
in01f80 FE_OCP_RBC2421_n_24505 ( .a(n_24505), .o(FE_OCP_RBN2421_n_24505) );
no02f80 g750988 ( .a(n_30001), .b(n_29946), .o(n_30002) );
in01f80 g754604 ( .a(n_26884), .o(n_26885) );
ao22s80 g778757 ( .a(n_2167), .b(n_1798), .c(n_2166), .d(n_1799), .o(n_2744) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_25_ ( .ck(newNet_1979), .d(n_12144), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_25_) );
in01f80 newInst_849 ( .a(newNet_369), .o(newNet_849) );
in01f80 FE_OCP_RBC3735_n_31819 ( .a(FE_OCP_RBN3733_n_31819), .o(FE_OCP_RBN3735_n_31819) );
na02f80 g745941 ( .a(n_34086), .b(n_34085), .o(n_34109) );
oa12f80 g776275 ( .a(n_4781), .b(n_4827), .c(n_4780), .o(n_4857) );
oa22f80 FE_RC_3738_0 ( .a(n_17177), .b(n_17487), .c(n_17176), .d(n_17512), .o(n_17688) );
no02f80 g750438 ( .a(n_29588), .b(n_29622), .o(n_29669) );
oa12f80 g778210 ( .a(n_2431), .b(n_2619), .c(n_2274), .o(n_2715) );
oa22f80 g764139 ( .a(n_16823), .b(n_16257), .c(n_16822), .d(n_16256), .o(n_16924) );
na02f80 g737718 ( .a(n_42392), .b(n_41988), .o(n_42747) );
in01f80 g745358 ( .a(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40598) );
in01f80 FE_OCP_RBC3477_n_13756 ( .a(n_13756), .o(FE_OCP_RBN3477_n_13756) );
no02f80 g746156 ( .a(n_33771), .b(n_34037), .o(n_33806) );
oa22f80 g752527 ( .a(n_27582), .b(n_27489), .c(n_45745), .d(n_27488), .o(n_27655) );
oa22f80 FE_RC_1448_0 ( .a(n_32287), .b(FE_OCP_RBN3128_n_32266), .c(n_28336), .d(n_32266), .o(n_32334) );
in01f80 g747413 ( .a(n_32704), .o(n_32709) );
na02f80 g769942 ( .a(n_11107), .b(n_11159), .o(n_11156) );
oa12f80 g770094 ( .a(n_10077), .b(n_10951), .c(n_9951), .o(n_11057) );
no02f80 g777003 ( .a(n_4025), .b(n_4121), .o(n_4096) );
no02f80 g767472 ( .a(n_13303), .b(n_13357), .o(n_13395) );
in01f80 g746999 ( .a(n_32835), .o(n_32836) );
in01f80 newInst_1007 ( .a(newNet_8), .o(newNet_1007) );
na02f80 g744488 ( .a(n_35416), .b(FE_OCPN1860_n_35415), .o(n_35429) );
no02f80 g760732 ( .a(n_19605), .b(n_18099), .o(n_19639) );
oa12f80 g739077 ( .a(n_40958), .b(n_41108), .c(n_41084), .o(n_41131) );
ao12f80 g750630 ( .a(n_30420), .b(n_30419), .c(n_30418), .o(n_31189) );
na02f80 g736991 ( .a(n_43242), .b(n_42771), .o(n_43519) );
ao12f80 g767723 ( .a(n_12748), .b(n_12863), .c(n_12860), .o(n_12938) );
in01f80 g740811 ( .a(n_39535), .o(n_39508) );
no02f80 g741998 ( .a(n_38084), .b(n_38057), .o(n_38399) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_12_ ( .ck(newNet_194), .d(n_46364), .o(delay_xor_ln22_unr9_stage4_stallmux_q_12_) );
in01f80 FE_OCP_RBC2122_n_45224 ( .a(FE_OCP_RBN2119_n_45224), .o(FE_OCP_RBN2122_n_45224) );
in01f80 g766911 ( .a(n_13560), .o(n_13575) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_30_ ( .ck(newNet_1811), .d(n_17102), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_30_) );
in01f80 g745797 ( .a(n_34119), .o(n_34100) );
no02f80 g761438 ( .a(n_18892), .b(FE_OFN779_n_17093), .o(n_18946) );
in01f80 g743086 ( .a(n_37051), .o(n_37052) );
in01f80 FE_RC_533_0 ( .a(FE_RN_167_0), .o(n_22632) );
in01f80 g758257 ( .a(n_22621), .o(n_22694) );
no02f80 g767969 ( .a(n_13079), .b(n_13076), .o(n_13717) );
no02f80 g778770 ( .a(n_2184), .b(n_2183), .o(n_2185) );
na02f80 g770895 ( .a(n_10127), .b(n_10027), .o(n_10170) );
in01f80 g781132 ( .a(n_219), .o(n_220) );
in01f80 g746227 ( .a(n_33697), .o(n_34504) );
no02f80 g761268 ( .a(n_19847), .b(n_20234), .o(n_19932) );
oa12f80 g739942 ( .a(n_40310), .b(n_40122), .c(n_39833), .o(n_40369) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_10_ ( .ck(newNet_2884), .d(n_10739), .o(delay_add_ln22_unr8_stage4_stallmux_q_10_) );
in01f80 g739020 ( .a(n_41462), .o(n_41140) );
ao12f80 g752119 ( .a(n_28618), .b(n_28617), .c(n_28616), .o(n_28939) );
no02f80 g753248 ( .a(n_27287), .b(n_27416), .o(n_27454) );
oa12f80 g749759 ( .a(n_30295), .b(n_30243), .c(n_29846), .o(n_30296) );
no02f80 g777807 ( .a(n_3251), .b(n_2913), .o(n_3308) );
in01f80 g752092 ( .a(n_28897), .o(n_28919) );
na02f80 g753965 ( .a(n_26220), .b(n_26216), .o(n_26251) );
no02f80 g761155 ( .a(n_19237), .b(n_19167), .o(n_19309) );
in01f80 newInst_3476 ( .a(newNet_3475), .o(newNet_3476) );
in01f80 newInst_2285 ( .a(newNet_2284), .o(newNet_2285) );
na02f80 g770901 ( .a(n_9723), .b(n_9674), .o(n_9807) );
na02f80 g764115 ( .a(n_16620), .b(n_16637), .o(n_16656) );
na02f80 g771267 ( .a(n_9313), .b(n_8232), .o(n_9492) );
in01f80 g741684 ( .a(n_38605), .o(n_38606) );
in01f80 newInst_399 ( .a(newNet_398), .o(newNet_399) );
oa12f80 g745117 ( .a(n_34664), .b(n_34663), .c(n_34662), .o(n_35665) );
no02f80 g780836 ( .a(n_395), .b(n_390), .o(n_543) );
ao12f80 g772426 ( .a(n_8640), .b(n_8639), .c(n_8638), .o(n_9598) );
in01f80 g751568 ( .a(n_28784), .o(n_28785) );
in01f80 g740176 ( .a(n_40036), .o(n_40117) );
ao12f80 g738147 ( .a(n_41741), .b(n_42027), .c(n_41762), .o(n_42038) );
in01f80 g770211 ( .a(n_10810), .o(n_10787) );
in01f80 newInst_1191 ( .a(newNet_1190), .o(newNet_1191) );
in01f80 g744598 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_0_), .o(n_35362) );
no02f80 g768396 ( .a(FE_OCP_RBN3394_n_12504), .b(n_12238), .o(n_12525) );
oa12f80 g768695 ( .a(n_11571), .b(n_44451), .c(n_11890), .o(n_12199) );
in01f80 newInst_2638 ( .a(newNet_2637), .o(newNet_2638) );
in01f80 g755287 ( .a(n_24986), .o(n_25011) );
no02f80 g745618 ( .a(n_34369), .b(n_33691), .o(n_34565) );
no02f80 g778035 ( .a(n_3038), .b(n_3058), .o(n_3059) );
oa12f80 g776818 ( .a(n_4085), .b(n_4139), .c(n_4084), .o(n_4192) );
no02f80 g773744 ( .a(n_7194), .b(n_7100), .o(n_7236) );
in01f80 g749044 ( .a(n_30965), .o(n_30966) );
in01f80 g781284 ( .a(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n_151) );
oa22f80 FE_RC_3444_0 ( .a(n_28677), .b(n_28964), .c(n_28676), .d(n_28963), .o(n_29054) );
na02f80 g766259 ( .a(n_14323), .b(n_14376), .o(n_14473) );
in01f80 g780391 ( .a(n_848), .o(n_827) );
in01f80 g772686 ( .a(n_8111), .o(n_8112) );
no02f80 g736953 ( .a(FE_OCPN912_n_43022), .b(n_42925), .o(n_43361) );
in01f80 g743653 ( .a(n_36381), .o(n_36416) );
na02f80 g777054 ( .a(n_3560), .b(n_2847), .o(n_3608) );
no02f80 FE_RC_3065_0 ( .a(FE_OCPN999_n_19311), .b(n_20694), .o(FE_RN_1347_0) );
in01f80 g760914 ( .a(n_19388), .o(n_19428) );
na02f80 FE_RC_2369_0 ( .a(FE_RN_916_0), .b(FE_RN_919_0), .o(n_2148) );
oa12f80 g756892 ( .a(n_23649), .b(n_23648), .c(n_23647), .o(n_24076) );
in01f80 g759722 ( .a(n_20678), .o(n_20679) );
in01f80 g768180 ( .a(n_13418), .o(n_13514) );
no02f80 g766491 ( .a(n_13996), .b(n_13028), .o(n_14067) );
no03m80 g751420 ( .a(n_28877), .b(n_29175), .c(n_28902), .o(n_29287) );
in01f80 g776221 ( .a(n_4741), .o(n_4742) );
ao12f80 g760058 ( .a(n_21100), .b(n_21099), .c(n_21098), .o(n_21593) );
ao22s80 FE_RC_805_0 ( .a(FE_OCP_RBN3464_n_7886), .b(n_8380), .c(n_8379), .d(FE_OCP_RBN2301_n_7817), .o(n_8491) );
in01f80 newInst_80 ( .a(newNet_79), .o(newNet_80) );
na02f80 FE_RC_1721_0 ( .a(FE_RN_474_0), .b(FE_RN_475_0), .o(FE_RN_476_0) );
oa12f80 g741793 ( .a(n_38058), .b(n_38322), .c(n_38084), .o(n_38462) );
no02f80 g776857 ( .a(n_3656), .b(n_3623), .o(n_3722) );
no02f80 g776079 ( .a(n_5048), .b(FE_OCP_RBN2659_n_4101), .o(n_4998) );
ao22s80 FE_RC_3670_0 ( .a(n_21289), .b(FE_OCP_RBN2950_n_21363), .c(n_21363), .d(FE_RN_1612_0), .o(n_21503) );
in01f80 FE_OCP_RBC3208_n_44365 ( .a(FE_OCP_RBN3210_n_44365), .o(FE_OCP_RBN3208_n_44365) );
in01f80 g761776 ( .a(n_19291), .o(n_19825) );
no02f80 g752127 ( .a(FE_OCPN878_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_11_), .o(n_28015) );
in01f80 newInst_3355 ( .a(newNet_3354), .o(newNet_3355) );
no02f80 g759631 ( .a(n_20680), .b(n_20722), .o(n_20789) );
na02f80 g753221 ( .a(n_27120), .b(FE_OCP_RBN2833_n_26081), .o(n_27222) );
no02f80 g763297 ( .a(n_16957), .b(n_17036), .o(n_17191) );
oa12f80 g745778 ( .a(n_34428), .b(n_44112), .c(n_34427), .o(n_34447) );
in01f80 FE_OCP_RBC2755_n_30558 ( .a(n_30558), .o(FE_OCP_RBN2755_n_30558) );
no02f80 g774087 ( .a(n_6832), .b(delay_add_ln22_unr5_stage3_stallmux_q_2_), .o(n_6910) );
in01f80 g772581 ( .a(n_8566), .o(n_8567) );
in01f80 g756206 ( .a(n_24102), .o(n_24125) );
na02f80 g774810 ( .a(n_6228), .b(n_5703), .o(n_6325) );
na02f80 g738065 ( .a(n_42116), .b(n_42115), .o(n_42117) );
no02f80 g764739 ( .a(n_15761), .b(n_14618), .o(n_15905) );
na02f80 g758106 ( .a(FE_OCPN1398_n_21973), .b(FE_OCP_RBN1336_n_20941), .o(n_22022) );
in01f80 FE_OCPC1006_n_13962 ( .a(FE_OCP_RBN2507_n_13896), .o(FE_OCPN1006_n_13962) );
in01f80 g772607 ( .a(n_8294), .o(n_8295) );
ao22s80 g737298 ( .a(n_42867), .b(n_42490), .c(n_42868), .d(n_42489), .o(n_42924) );
no02f80 g762082 ( .a(n_18242), .b(n_17625), .o(n_18337) );
in01f80 newInst_886 ( .a(newNet_885), .o(newNet_886) );
ao12f80 FE_RC_1894_0 ( .a(FE_RN_590_0), .b(FE_RN_591_0), .c(n_12036), .o(n_12173) );
in01f80 g752766 ( .a(n_27955), .o(n_27956) );
in01f80 g757590 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .o(n_22768) );
no02f80 g745752 ( .a(n_47254), .b(n_34256), .o(n_34281) );
no02f80 FE_RC_1912_0 ( .a(n_17732), .b(n_18987), .o(FE_RN_601_0) );
in01f80 g749508 ( .a(n_30598), .o(n_31599) );
no02f80 g749608 ( .a(n_30461), .b(n_30460), .o(n_30462) );
oa12f80 g739260 ( .a(n_40669), .b(n_40699), .c(n_40739), .o(n_40801) );
na02f80 g754892 ( .a(FE_OCP_RBN2596_n_25181), .b(n_24458), .o(n_25452) );
no02f80 g766896 ( .a(n_13740), .b(n_13739), .o(n_13741) );
ao12f80 g752160 ( .a(n_27866), .b(n_28009), .c(n_27867), .o(n_28120) );
in01f80 newInst_665 ( .a(newNet_664), .o(newNet_665) );
in01f80 g746816 ( .a(n_33265), .o(n_33266) );
na02f80 g764569 ( .a(n_15817), .b(n_14588), .o(n_15860) );
na02f80 g772996 ( .a(n_8172), .b(n_8119), .o(n_8173) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_10_ ( .ck(newNet_2424), .d(n_36337), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_) );
ao12f80 g767084 ( .a(n_13735), .b(n_13734), .c(n_13733), .o(n_14253) );
no02f80 g776888 ( .a(n_3893), .b(n_3927), .o(n_4113) );
na02f80 g748146 ( .a(n_31741), .b(n_31773), .o(n_31807) );
ao12f80 g775428 ( .a(n_4871), .b(n_5711), .c(n_4885), .o(n_5814) );
na02f80 g747983 ( .a(n_33040), .b(n_32645), .o(n_33116) );
no02f80 g774320 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_12_), .o(n_6870) );
in01f80 g766172 ( .a(n_14894), .o(n_14895) );
na02f80 g763249 ( .a(FE_OCP_RBN1134_n_16041), .b(n_17140), .o(n_17141) );
in01f80 FE_RC_3069_0 ( .a(n_23353), .o(FE_RN_1349_0) );
in01f80 g773340 ( .a(n_8189), .o(n_8309) );
na02f80 g759784 ( .a(n_21599), .b(n_21374), .o(n_21671) );
in01f80 newInst_176 ( .a(newNet_144), .o(newNet_176) );
na02f80 g767943 ( .a(n_12628), .b(n_12447), .o(n_12669) );
no02f80 g746076 ( .a(n_33873), .b(n_33846), .o(n_33901) );
in01f80 newInst_3706 ( .a(newNet_1044), .o(newNet_3706) );
in01f80 g743527 ( .a(n_36516), .o(n_36517) );
no02f80 g741810 ( .a(n_38469), .b(n_38468), .o(n_38470) );
no02f80 g748801 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_28_), .o(n_32537) );
in01f80 g738158 ( .a(n_42035), .o(n_42036) );
in01f80 fopt782978 ( .a(n_17729), .o(n_44447) );
in01f80 FE_OCPC901_n_44593 ( .a(FE_OCPN899_n_44593), .o(FE_OCPN901_n_44593) );
in01f80 newInst_2197 ( .a(newNet_529), .o(newNet_2197) );
no02f80 g742601 ( .a(n_37547), .b(n_37499), .o(n_37568) );
in01f80 newInst_811 ( .a(newNet_810), .o(newNet_811) );
ao12f80 g780753 ( .a(n_569), .b(n_576), .c(n_568), .o(n_719) );
oa12f80 g739895 ( .a(n_40291), .b(n_40123), .c(n_40214), .o(n_40343) );
in01f80 FE_OCP_RBC3078_FE_OFN807_n_46195 ( .a(FE_OFN807_n_46195), .o(FE_OCP_RBN3078_FE_OFN807_n_46195) );
no02f80 g768415 ( .a(n_12492), .b(n_12147), .o(n_12504) );
na02f80 FE_RC_3125_0 ( .a(FE_OCP_RBN1201_n_25763), .b(FE_RN_1384_0), .o(FE_RN_1385_0) );
no02f80 FE_RC_4182_0 ( .a(FE_RN_1827_0), .b(FE_RN_1828_0), .o(n_33942) );
na02f80 g745734 ( .a(n_34117), .b(n_34130), .o(n_34131) );
ao22s80 g778567 ( .a(n_2251), .b(n_1488), .c(n_2252), .d(n_1487), .o(n_2878) );
in01f80 g773507 ( .a(n_7516), .o(n_7510) );
no02f80 g747121 ( .a(n_32742), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_7_), .o(n_32788) );
in01f80 g765627 ( .a(n_14964), .o(n_14965) );
no02f80 g753576 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_27931) );
no02f80 g758943 ( .a(n_21286), .b(n_19716), .o(n_21432) );
in01f80 g763119 ( .a(n_17200), .o(n_17201) );
in01f80 g769033 ( .a(n_11975), .o(n_11899) );
na02f80 g768014 ( .a(n_12761), .b(n_12461), .o(n_12818) );
no02f80 g759938 ( .a(FE_OCP_RBN3679_n_21051), .b(n_21370), .o(n_21450) );
in01f80 g747563 ( .a(n_32516), .o(n_32465) );
oa12f80 g767651 ( .a(n_12564), .b(n_12727), .c(n_12539), .o(n_12802) );
oa22f80 FE_RC_3803_0 ( .a(n_25355), .b(n_25633), .c(n_25356), .d(n_25602), .o(n_25729) );
in01f80 g748057 ( .a(n_31954), .o(n_31972) );
no02f80 g760367 ( .a(n_20191), .b(n_20170), .o(n_20209) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_1_ ( .ck(newNet_1319), .d(n_1140), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_) );
oa12f80 g739267 ( .a(n_44769), .b(n_40900), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n_40905) );
na02f80 g750484 ( .a(n_29506), .b(n_29484), .o(n_29566) );
no02f80 g762138 ( .a(n_18776), .b(n_18766), .o(n_19402) );
no02f80 g772742 ( .a(n_8133), .b(n_47240), .o(n_8195) );
in01f80 g781351 ( .a(beta_28), .o(n_88) );
in01f80 g746498 ( .a(n_33330), .o(n_33453) );
no02f80 g749301 ( .a(n_46959), .b(n_27130), .o(n_30682) );
no02f80 g759652 ( .a(n_20615), .b(n_20547), .o(n_20641) );
in01f80 g743059 ( .a(n_37173), .o(n_37174) );
in01f80 newInst_2987 ( .a(newNet_2986), .o(newNet_2987) );
in01f80 g746522 ( .a(n_34668), .o(n_34669) );
oa22f80 FE_RC_1704_0 ( .a(n_32287), .b(FE_OCP_RBN3112_n_32254), .c(n_28336), .d(n_32254), .o(n_32304) );
na02f80 g776045 ( .a(n_47004), .b(n_5178), .o(n_5226) );
in01f80 g768441 ( .a(n_12436), .o(n_12437) );
in01f80 g750625 ( .a(n_29417), .o(n_29442) );
no02f80 g781231 ( .a(n_82), .b(n_81), .o(n_83) );
in01f80 newInst_257 ( .a(newNet_256), .o(newNet_257) );
na02f80 g756594 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_), .o(n_23966) );
ao12f80 g746937 ( .a(n_32719), .b(n_32834), .c(n_32722), .o(n_32924) );
na02f80 g750078 ( .a(n_29896), .b(n_29472), .o(n_30245) );
ao12f80 g738971 ( .a(n_41148), .b(n_41147), .c(n_41146), .o(n_41190) );
in01f80 g744397 ( .a(n_35516), .o(n_35529) );
in01f80 FE_OCP_RBC3064_n_22170 ( .a(n_22170), .o(FE_OCP_RBN3064_n_22170) );
na02f80 g742769 ( .a(n_37316), .b(n_37150), .o(n_37350) );
in01f80 g768833 ( .a(n_11956), .o(n_11917) );
in01f80 g749955 ( .a(n_30014), .o(n_30015) );
no02f80 g742681 ( .a(n_37483), .b(n_37482), .o(n_37484) );
na02f80 g755387 ( .a(n_25494), .b(n_25493), .o(n_25495) );
in01f80 g739578 ( .a(n_40647), .o(n_40637) );
na02f80 FE_RC_2292_0 ( .a(FE_RN_858_0), .b(FE_RN_861_0), .o(n_18421) );
no02f80 g760053 ( .a(n_20574), .b(n_20556), .o(n_20672) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_30_ ( .ck(newNet_2257), .d(n_40578), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_) );
in01f80 g756363 ( .a(n_24645), .o(n_24066) );
no02f80 g748122 ( .a(n_31835), .b(n_31850), .o(n_31907) );
in01f80 g776826 ( .a(n_3786), .o(n_3731) );
na02f80 g772517 ( .a(n_8645), .b(n_8644), .o(n_8646) );
in01f80 newInst_3243 ( .a(newNet_3242), .o(newNet_3243) );
ao22s80 FE_RC_1375_0 ( .a(FE_RN_470_0), .b(n_25692), .c(n_25691), .d(FE_OCP_RBN3671_FE_RN_470_0), .o(n_26171) );
in01f80 g757746 ( .a(n_22769), .o(n_22575) );
na02f80 g770497 ( .a(FE_OCP_RBN2904_n_10474), .b(n_10434), .o(n_10501) );
in01f80 g761443 ( .a(n_20176), .o(n_20177) );
na02f80 g755444 ( .a(n_24661), .b(n_24761), .o(n_24662) );
no02f80 g773591 ( .a(n_7425), .b(n_7424), .o(n_7447) );
na02f80 g750085 ( .a(FE_OCP_RBN3561_n_29857), .b(n_29032), .o(n_30021) );
in01f80 newInst_106 ( .a(newNet_105), .o(newNet_106) );
in01f80 g769047 ( .a(n_11762), .o(n_11730) );
in01f80 g767026 ( .a(n_14427), .o(n_14293) );
ao12f80 g777389 ( .a(n_3548), .b(n_3522), .c(n_3615), .o(n_3631) );
in01f80 g740008 ( .a(n_40255), .o(n_40225) );
in01f80 FE_OCP_RBC2371_n_8221 ( .a(n_8221), .o(FE_OCP_RBN2371_n_8221) );
na02f80 g744471 ( .a(n_35458), .b(n_35447), .o(n_35501) );
oa12f80 g760248 ( .a(n_20196), .b(n_20834), .c(n_20234), .o(n_21023) );
in01f80 g740557 ( .a(n_39668), .o(n_39645) );
no02f80 g777114 ( .a(n_3989), .b(n_3912), .o(n_4058) );
in01f80 FE_RC_2683_0 ( .a(FE_OCPN1392_n_7925), .o(FE_RN_1122_0) );
in01f80 FE_OCP_RBC2273_n_2457 ( .a(n_2457), .o(FE_OCP_RBN2273_n_2457) );
in01f80 g768613 ( .a(n_12256), .o(n_12257) );
no02f80 g763089 ( .a(n_17147), .b(n_17046), .o(n_17292) );
no02f80 g752288 ( .a(FE_OCP_RBN2179_FE_RN_526_0), .b(n_28109), .o(n_28538) );
na02f80 g776344 ( .a(n_4580), .b(n_4565), .o(n_4792) );
in01f80 FE_OCPC3791_n_36069 ( .a(FE_OCPN3790_n_36069), .o(FE_OCPN3791_n_36069) );
in01f80 FE_OCP_RBC3205_n_44365 ( .a(FE_OCP_RBN3206_n_44365), .o(FE_OCP_RBN3205_n_44365) );
in01f80 g752218 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_13_), .o(n_27921) );
no02f80 g784081 ( .a(n_8199), .b(n_45820), .o(n_45827) );
no02f80 g748367 ( .a(n_32748), .b(n_32747), .o(n_32749) );
na02f80 g766290 ( .a(n_14438), .b(n_14402), .o(n_14535) );
no02f80 g768078 ( .a(n_12790), .b(n_12789), .o(n_12854) );
ao12f80 g769982 ( .a(n_11041), .b(n_11057), .c(n_10036), .o(n_11069) );
in01f80 g737873 ( .a(n_42614), .o(n_42615) );
oa12f80 g745697 ( .a(n_34190), .b(n_34189), .c(n_34191), .o(n_35415) );
na02f80 g745832 ( .a(FE_OCP_RBN3438_n_33750), .b(n_44104), .o(n_34242) );
in01f80 g765215 ( .a(n_15305), .o(n_15306) );
in01f80 g749766 ( .a(n_31319), .o(n_31320) );
in01f80 g777199 ( .a(n_3593), .o(n_3635) );
na02f80 g760815 ( .a(n_19435), .b(n_19201), .o(n_19518) );
na02f80 g779065 ( .a(n_2000), .b(n_1845), .o(n_2063) );
no02f80 g746517 ( .a(n_34803), .b(n_34840), .o(n_34888) );
na02f80 g743804 ( .a(n_36308), .b(n_36305), .o(n_36369) );
oa12f80 g762662 ( .a(n_17353), .b(n_18237), .c(n_17572), .o(n_18253) );
ao12f80 g778012 ( .a(n_2749), .b(n_3013), .c(n_2816), .o(n_3030) );
oa12f80 g739480 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_16_), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_), .o(n_40713) );
no02f80 g778633 ( .a(n_2913), .b(n_2807), .o(n_2937) );
no02f80 g758069 ( .a(n_22694), .b(n_22693), .o(n_22981) );
no02f80 g777991 ( .a(FE_OCP_RBN2425_n_47023), .b(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(n_3079) );
na02f80 g769694 ( .a(n_11247), .b(n_11168), .o(n_11245) );
oa12f80 g763224 ( .a(n_17712), .b(n_17736), .c(n_17711), .o(n_17785) );
ao12f80 g779656 ( .a(n_1620), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n_1778) );
in01f80 FE_RC_2585_0 ( .a(n_17825), .o(FE_RN_1068_0) );
oa12f80 g751748 ( .a(n_28919), .b(n_29104), .c(n_29172), .o(n_29174) );
in01f80 newInst_2295 ( .a(newNet_2294), .o(newNet_2295) );
in01f80 g740714 ( .a(n_39495), .o(n_39496) );
oa12f80 g751808 ( .a(n_28181), .b(n_28255), .c(n_28139), .o(n_28268) );
no02f80 g761287 ( .a(n_19035), .b(n_18985), .o(n_19083) );
na02f80 g760095 ( .a(FE_OCP_RBN1343_n_19077), .b(n_20372), .o(n_20469) );
no02f80 g748678 ( .a(n_32796), .b(n_32494), .o(n_32781) );
na02f80 g763043 ( .a(n_17252), .b(n_17293), .o(n_17460) );
no02f80 g758193 ( .a(n_22438), .b(n_22366), .o(n_22457) );
no02f80 g744836 ( .a(n_35029), .b(FE_OCPN1796_n_30546), .o(n_35118) );
no02f80 g744806 ( .a(n_35143), .b(FE_OCPN1434_n_30614), .o(n_35169) );
no02f80 g747723 ( .a(n_33680), .b(n_33599), .o(n_34171) );
in01f80 g771369 ( .a(n_9611), .o(n_9612) );
in01f80 FE_OCP_RBC2991_n_35539 ( .a(FE_OCP_RBN2989_n_35539), .o(FE_OCP_RBN2991_n_35539) );
in01f80 g739862 ( .a(n_40263), .o(n_40264) );
na02f80 g771621 ( .a(n_9275), .b(FE_OFN361_n_9391), .o(n_9687) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_11_ ( .ck(newNet_3453), .d(n_27160), .o(delay_add_ln22_unr17_stage7_stallmux_q_11_) );
na02f80 g739053 ( .a(n_41092), .b(n_41041), .o(n_41117) );
no02f80 g760082 ( .a(n_20245), .b(FE_OFN751_n_45003), .o(n_20294) );
na02f80 g767978 ( .a(n_12717), .b(n_12860), .o(n_12821) );
in01f80 g777930 ( .a(n_3183), .o(n_3184) );
no02f80 FE_RC_2287_0 ( .a(n_17093), .b(FE_RN_856_0), .o(FE_RN_857_0) );
no02f80 g756784 ( .a(n_23409), .b(n_23408), .o(n_23410) );
na02f80 g749908 ( .a(n_29968), .b(n_29901), .o(n_30247) );
na02f80 g768874 ( .a(n_12124), .b(n_11871), .o(n_11875) );
ao22s80 g775484 ( .a(n_5398), .b(n_4875), .c(n_5397), .d(n_4759), .o(n_5543) );
in01f80 g779649 ( .a(n_1489), .o(n_1490) );
na02f80 g758191 ( .a(n_22399), .b(n_22368), .o(n_22498) );
oa22f80 g763624 ( .a(n_46977), .b(FE_OFN767_n_15670), .c(n_16705), .d(n_17753), .o(n_16789) );
ao12f80 g749901 ( .a(n_30184), .b(n_30969), .c(n_30186), .o(n_31091) );
na02f80 g779571 ( .a(n_1792), .b(n_1514), .o(n_1809) );
na02f80 g775530 ( .a(n_5506), .b(n_5559), .o(n_5592) );
na02f80 g764477 ( .a(n_16056), .b(n_16092), .o(n_16231) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_31_ ( .ck(newNet_2447), .d(n_32516), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_) );
in01f80 g765533 ( .a(n_15709), .o(n_15830) );
in01f80 g746611 ( .a(n_34417), .o(n_34418) );
no02f80 g743545 ( .a(n_37611), .b(n_37631), .o(n_37713) );
in01f80 newInst_2830 ( .a(newNet_2829), .o(newNet_2830) );
na02f80 g773433 ( .a(n_7530), .b(n_7512), .o(n_7540) );
oa22f80 FE_RC_3437_0 ( .a(n_22498), .b(n_22740), .c(n_22499), .d(FE_OCP_RBN1704_n_22740), .o(n_22897) );
oa12f80 g747192 ( .a(n_32786), .b(n_32817), .c(n_32848), .o(n_32885) );
in01f80 FE_RC_681_0 ( .a(n_32702), .o(FE_RN_220_0) );
ao12f80 g763129 ( .a(n_17368), .b(n_17787), .c(n_17298), .o(n_17863) );
in01f80 g768701 ( .a(n_12238), .o(n_12239) );
in01f80 newInst_3232 ( .a(newNet_3231), .o(newNet_3232) );
no02f80 FE_RC_2142_0 ( .a(n_46419), .b(n_15144), .o(FE_RN_752_0) );
in01f80 FE_OCP_RBC2678_n_9247 ( .a(n_9247), .o(FE_OCP_RBN2678_n_9247) );
oa12f80 g739019 ( .a(n_41118), .b(n_41117), .c(n_41116), .o(n_41490) );
no02f80 g765306 ( .a(FE_OFN764_n_15670), .b(n_15748), .o(n_15840) );
no02f80 g744770 ( .a(n_35173), .b(n_35197), .o(n_35287) );
in01f80 g754075 ( .a(n_26194), .o(n_26195) );
na02f80 g759343 ( .a(n_21888), .b(n_21887), .o(n_21889) );
no02f80 g760313 ( .a(n_20081), .b(n_19921), .o(n_20154) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_30_ ( .ck(newNet_2919), .d(n_6648), .o(delay_add_ln22_unr5_stage3_stallmux_q_30_) );
na02f80 g770138 ( .a(n_10828), .b(FE_OCP_RBN2654_n_9198), .o(n_10940) );
na02f80 g762235 ( .a(n_18163), .b(delay_add_ln22_unr11_stage5_stallmux_q_16_), .o(n_18187) );
in01f80 g746108 ( .a(n_33780), .o(n_33781) );
in01f80 g773442 ( .a(n_8846), .o(n_7691) );
in01f80 g774999 ( .a(n_6102), .o(n_6000) );
in01f80 g739815 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .o(n_40460) );
in01f80 newInst_2218 ( .a(newNet_777), .o(newNet_2218) );
in01f80 FE_OFC49_n_1045 ( .a(n_1045), .o(FE_OFN49_n_1045) );
na02f80 g746593 ( .a(n_34666), .b(n_34735), .o(n_34756) );
no02f80 g743418 ( .a(n_36626), .b(n_36750), .o(n_36689) );
no02f80 g771273 ( .a(n_9261), .b(n_9089), .o(n_9262) );
in01f80 g758909 ( .a(n_21705), .o(n_21648) );
oa22f80 FE_RC_3214_0 ( .a(n_1142), .b(n_44652), .c(n_1130), .d(n_44661), .o(n_1299) );
in01f80 g739968 ( .a(n_40086), .o(n_40122) );
na02f80 g754518 ( .a(n_26739), .b(n_26685), .o(n_26792) );
na02f80 g780916 ( .a(n_403), .b(n_402), .o(n_411) );
ao22s80 g746285 ( .a(n_33616), .b(n_33544), .c(n_33523), .d(n_32728), .o(n_33640) );
na02f80 g743696 ( .a(n_37362), .b(n_46212), .o(n_37436) );
no02f80 FE_RC_2926_0 ( .a(FE_RN_1273_0), .b(FE_RN_1274_0), .o(n_27554) );
no02f80 FE_RC_1640_0 ( .a(FE_RN_456_0), .b(FE_RN_457_0), .o(FE_RN_458_0) );
na02f80 g767673 ( .a(n_13238), .b(n_13777), .o(n_13260) );
na02f80 g738543 ( .a(n_41618), .b(n_41572), .o(n_41666) );
oa12f80 g738303 ( .a(n_41424), .b(n_41648), .c(n_41455), .o(n_41799) );
in01f80 g778263 ( .a(n_2997), .o(n_2998) );
no02f80 g767549 ( .a(n_12944), .b(n_12639), .o(n_13007) );
oa22f80 FE_RC_217_0 ( .a(n_11763), .b(FE_OCP_RBN2137_n_11907), .c(n_11907), .d(FE_OCP_RBN2150_n_11763), .o(n_12062) );
in01f80 FE_OCP_RBC2779_n_15595 ( .a(FE_OCP_RBN2778_n_15595), .o(FE_OCP_RBN2779_n_15595) );
oa12f80 g770160 ( .a(n_10653), .b(n_10813), .c(n_10864), .o(n_10892) );
in01f80 g744130 ( .a(n_35638), .o(n_35639) );
oa12f80 g757769 ( .a(FE_OCP_RBN1709_n_22150), .b(n_22468), .c(n_22531), .o(n_22574) );
na02f80 g744553 ( .a(n_35394), .b(n_35418), .o(n_35456) );
in01f80 g751305 ( .a(n_28748), .o(n_28708) );
in01f80 FE_OCP_RBC2665_n_35207 ( .a(n_35207), .o(FE_OCP_RBN2665_n_35207) );
in01f80 g780254 ( .a(n_1025), .o(n_989) );
in01f80 g777514 ( .a(n_4675), .o(n_5494) );
no02f80 g784590 ( .a(n_32643), .b(FE_OCP_RBN3370_n_32436), .o(n_46413) );
no02f80 g759275 ( .a(n_20865), .b(n_20830), .o(n_20951) );
in01f80 g775762 ( .a(n_5532), .o(n_5533) );
oa22f80 g747757 ( .a(n_32032), .b(n_31737), .c(n_32033), .d(n_31736), .o(n_32113) );
na02f80 g745256 ( .a(n_36083), .b(n_36121), .o(n_36084) );
in01f80 g739164 ( .a(n_40990), .o(n_40975) );
in01f80 g745026 ( .a(n_34878), .o(n_34879) );
na02f80 g753991 ( .a(n_26975), .b(n_26864), .o(n_27031) );
na02f80 g754864 ( .a(n_25242), .b(n_25241), .o(n_25243) );
na02f80 g765139 ( .a(n_15884), .b(n_15874), .o(n_15976) );
in01f80 newInst_1344 ( .a(newNet_723), .o(newNet_1344) );
in01f80 FE_OCP_RBC2976_n_5555 ( .a(n_5555), .o(FE_OCP_RBN2976_n_5555) );
in01f80 newInst_3334 ( .a(newNet_30), .o(newNet_3334) );
in01f80 g744537 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_24_), .o(n_36713) );
oa22f80 FE_RC_829_0 ( .a(n_9493), .b(n_9574), .c(n_9476), .d(n_9573), .o(n_9724) );
ao22s80 FE_RC_1299_0 ( .a(n_39447), .b(n_39188), .c(n_39187), .d(n_39446), .o(n_39542) );
in01f80 g767602 ( .a(n_13005), .o(n_14153) );
na02f80 g756935 ( .a(n_23808), .b(n_23807), .o(n_23809) );
no02f80 g754314 ( .a(n_25830), .b(n_25793), .o(n_25898) );
in01f80 FE_OCP_RBC3685_n_5217 ( .a(n_5217), .o(FE_OCP_RBN3685_n_5217) );
oa22f80 g753542 ( .a(n_27368), .b(n_26924), .c(n_27367), .d(n_26925), .o(n_27479) );
na02f80 g775305 ( .a(n_6007), .b(n_5916), .o(n_5980) );
na02f80 g767933 ( .a(n_12664), .b(n_12683), .o(n_12684) );
in01f80 g747792 ( .a(n_33418), .o(n_33373) );
no02f80 g748607 ( .a(n_31492), .b(n_31237), .o(n_31515) );
in01f80 g766341 ( .a(n_15250), .o(n_14364) );
in01f80 newInst_1326 ( .a(newNet_1325), .o(newNet_1326) );
na02f80 g778198 ( .a(n_3006), .b(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(n_2743) );
in01f80 FE_OCP_RBC3369_n_32436 ( .a(FE_OCP_RBN3368_n_32436), .o(FE_OCP_RBN3369_n_32436) );
oa12f80 g778115 ( .a(n_2846), .b(n_2845), .c(n_2844), .o(n_4207) );
no02f80 g737611 ( .a(n_42240), .b(n_42220), .o(n_42266) );
no02f80 g747433 ( .a(n_32731), .b(n_32620), .o(n_32659) );
no03m80 g743598 ( .a(n_37541), .b(n_37474), .c(n_37540), .o(n_37542) );
na02f80 g754981 ( .a(n_25381), .b(n_25315), .o(n_25451) );
no02f80 g736466 ( .a(n_43716), .b(n_43330), .o(n_43742) );
in01f80 g752575 ( .a(n_28810), .o(n_28327) );
na02f80 g760197 ( .a(FE_OCP_RBN3616_n_20249), .b(n_20266), .o(n_20603) );
na02f80 g776020 ( .a(n_5080), .b(n_5079), .o(n_5081) );
na02f80 g772811 ( .a(n_8103), .b(n_8158), .o(n_8192) );
in01f80 FE_RC_1890_0 ( .a(n_23000), .o(FE_RN_589_0) );
na02f80 g738347 ( .a(n_41812), .b(n_41815), .o(n_41858) );
in01f80 newInst_2962 ( .a(newNet_2961), .o(newNet_2962) );
in01f80 fopt782970 ( .a(n_32339), .o(n_44434) );
in01f80 FE_OCP_RBC3523_n_8242 ( .a(FE_OCP_RBN2407_n_8242), .o(FE_OCP_RBN3523_n_8242) );
in01f80 g746679 ( .a(n_34473), .o(n_34612) );
in01f80 newInst_3152 ( .a(newNet_3151), .o(newNet_3152) );
in01f80 FE_RC_3273_0 ( .a(FE_RN_1441_0), .o(FE_RN_1440_0) );
in01f80 FE_RC_3200_0 ( .a(n_7578), .o(FE_RN_1421_0) );
no02f80 g767982 ( .a(n_12749), .b(n_12719), .o(n_12937) );
in01f80 newInst_858 ( .a(newNet_857), .o(newNet_858) );
na02f80 g779294 ( .a(n_1724), .b(n_1679), .o(n_1760) );
na02f80 g759045 ( .a(n_21127), .b(n_45091), .o(n_21288) );
na02f80 g780289 ( .a(n_908), .b(n_1148), .o(n_909) );
na02f80 g765833 ( .a(n_15290), .b(n_15247), .o(n_15248) );
in01f80 g774515 ( .a(n_6540), .o(n_6541) );
no02f80 g745160 ( .a(n_36056), .b(n_36055), .o(n_36127) );
na02f80 g752780 ( .a(n_27312), .b(n_27357), .o(n_27434) );
in01f80 g778173 ( .a(n_2902), .o(n_2903) );
no02f80 g764613 ( .a(n_15987), .b(n_15845), .o(n_16035) );
in01f80 g765511 ( .a(n_15749), .o(n_15717) );
in01f80 FE_OCP_RBC1163_n_13726 ( .a(n_13726), .o(FE_OCP_RBN1163_n_13726) );
na02f80 g767585 ( .a(n_13055), .b(n_13054), .o(n_13056) );
in01f80 drc784076 ( .a(n_45820), .o(n_45821) );
no02f80 FE_RC_2343_0 ( .a(FE_RN_897_0), .b(n_18696), .o(FE_RN_898_0) );
no02f80 g741066 ( .a(n_38893), .b(FE_OCP_RBN2547_n_44944), .o(n_38963) );
in01f80 g744402 ( .a(n_35532), .o(n_35499) );
no02f80 g739336 ( .a(n_40676), .b(delay_add_ln22_unr27_stage10_stallmux_q_3_), .o(n_40693) );
in01f80 newInst_2435 ( .a(newNet_2434), .o(newNet_2435) );
in01f80 g772639 ( .a(n_8348), .o(n_8366) );
no02f80 g746768 ( .a(n_32922), .b(n_32860), .o(n_32965) );
no02f80 g750921 ( .a(n_29015), .b(n_29014), .o(n_29016) );
in01f80 g760688 ( .a(n_19744), .o(n_19772) );
in01f80 g775362 ( .a(n_5840), .o(n_5789) );
na03f80 g742783 ( .a(n_37288), .b(n_37291), .c(n_36970), .o(n_37289) );
na02f80 g749588 ( .a(n_30286), .b(n_30016), .o(n_30377) );
na02f80 g760727 ( .a(n_19589), .b(n_18119), .o(n_19661) );
no02f80 g778941 ( .a(n_2260), .b(n_2253), .o(n_2254) );
na02f80 g754716 ( .a(FE_OCPN928_n_26231), .b(n_26507), .o(n_26547) );
in01f80 g740725 ( .a(n_39566), .o(n_39567) );
no02f80 g742205 ( .a(n_44867), .b(n_37884), .o(n_37886) );
no02f80 g747583 ( .a(n_33361), .b(n_33257), .o(n_33397) );
na02f80 g740244 ( .a(n_39852), .b(n_39891), .o(n_39892) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_17_ ( .ck(newNet_1242), .d(n_5853), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_17_) );
na02f80 g741657 ( .a(n_38539), .b(n_38239), .o(n_38556) );
na02f80 g737887 ( .a(n_42202), .b(n_42130), .o(n_42307) );
in01f80 newInst_3095 ( .a(newNet_659), .o(newNet_3095) );
in01f80 newInst_313 ( .a(newNet_312), .o(newNet_313) );
no02f80 g750965 ( .a(n_30811), .b(n_30163), .o(n_30229) );
in01f80 newInst_1253 ( .a(newNet_1252), .o(newNet_1253) );
ao12f80 g779650 ( .a(n_1445), .b(n_1452), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_26_), .o(n_1489) );
na02f80 g779296 ( .a(n_1702), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .o(n_1784) );
na02f80 g774185 ( .a(n_6942), .b(n_6939), .o(n_6943) );
na02f80 g757334 ( .a(n_23123), .b(n_23186), .o(n_23223) );
na02f80 g760147 ( .a(n_20456), .b(n_19663), .o(n_20705) );
no02f80 g743011 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_36960) );
in01f80 FE_RC_4255_0 ( .a(FE_OCP_DRV_N3168_FE_RN_1789_0), .o(FE_RN_1873_0) );
na02f80 g741628 ( .a(FE_OCP_RBN3502_n_38592), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38625) );
in01f80 g750645 ( .a(n_29396), .o(n_29397) );
in01f80 g736983 ( .a(n_43389), .o(n_43422) );
na02f80 g757255 ( .a(n_44068), .b(delay_xor_ln22_unr15_stage6_stallmux_q_16_), .o(n_23112) );
oa22f80 g776530 ( .a(n_4101), .b(n_3029), .c(FE_OCP_RBN2658_n_4101), .d(n_3862), .o(n_4343) );
in01f80 FE_OCP_RBC2368_n_38545 ( .a(n_38545), .o(FE_OCP_RBN2368_n_38545) );
in01f80 newInst_1084 ( .a(newNet_1063), .o(newNet_1084) );
ao12f80 g752842 ( .a(n_27991), .b(n_27762), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n_28023) );
no02f80 g780998 ( .a(n_284), .b(n_108), .o(n_283) );
in01f80 g753788 ( .a(n_27095), .o(n_27096) );
no02f80 g779085 ( .a(n_2023), .b(n_2013), .o(n_2014) );
na02f80 g744687 ( .a(n_35235), .b(FE_OCP_RBN2683_n_35213), .o(n_35236) );
oa12f80 g751328 ( .a(n_28403), .b(n_28612), .c(n_28357), .o(n_28685) );
in01f80 g770155 ( .a(n_10920), .o(n_10921) );
na02f80 g775922 ( .a(n_5177), .b(n_5152), .o(n_5315) );
na02f80 g753729 ( .a(n_26529), .b(FE_OCPN1496_n_26528), .o(n_26616) );
no02f80 g772435 ( .a(n_8580), .b(n_7900), .o(n_8594) );
in01f80 g775811 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_7_), .o(n_5362) );
no02f80 g747260 ( .a(n_33724), .b(n_33481), .o(n_33798) );
na02f80 g780598 ( .a(n_779), .b(n_867), .o(n_977) );
in01f80 g780267 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_5_), .o(n_1032) );
na02f80 g741979 ( .a(n_37956), .b(n_37955), .o(n_37957) );
no02f80 g760480 ( .a(n_19972), .b(n_19816), .o(n_20049) );
na02f80 g771858 ( .a(n_10154), .b(n_10038), .o(n_10206) );
in01f80 g746483 ( .a(n_34844), .o(n_34813) );
na02f80 g755040 ( .a(n_25206), .b(n_25205), .o(n_25232) );
na02f80 g748362 ( .a(n_31729), .b(n_31760), .o(n_31825) );
na02f80 g754465 ( .a(n_26938), .b(n_26419), .o(n_26420) );
in01f80 g774794 ( .a(n_6265), .o(n_6295) );
no02f80 g780475 ( .a(n_767), .b(n_724), .o(n_1159) );
na02f80 g779233 ( .a(n_1889), .b(n_1600), .o(n_1924) );
no02f80 g764754 ( .a(n_15732), .b(n_15731), .o(n_15845) );
in01f80 g779745 ( .a(n_1580), .o(n_1553) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_21_ ( .ck(newNet_2096), .d(n_6301), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_) );
no02f80 g746142 ( .a(n_33869), .b(n_33406), .o(n_33937) );
no02f80 g773155 ( .a(n_7712), .b(n_7714), .o(n_7767) );
in01f80 g761202 ( .a(n_19107), .o(n_19108) );
na02f80 g768543 ( .a(n_12230), .b(delay_add_ln22_unr8_stage4_stallmux_q_8_), .o(n_12299) );
in01f80 g737667 ( .a(n_42726), .o(n_42727) );
na02f80 g752671 ( .a(n_28261), .b(n_28153), .o(n_28263) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_1_ ( .ck(newNet_2196), .d(n_1007), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_1_) );
in01f80 FE_OCP_RBC3650_n_35169 ( .a(n_35169), .o(FE_OCP_RBN3650_n_35169) );
in01f80 g740360 ( .a(n_39751), .o(n_39752) );
in01f80 g740574 ( .a(n_39695), .o(n_39765) );
in01f80 g756008 ( .a(n_25679), .o(n_25680) );
na02f80 g766114 ( .a(n_14605), .b(n_14550), .o(n_14632) );
in01f80 FE_OCPC1515_n_35367 ( .a(n_35367), .o(FE_OCPN1515_n_35367) );
oa12f80 g764183 ( .a(n_16313), .b(n_16848), .c(n_16262), .o(n_16887) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_28_ ( .ck(newNet_3295), .d(n_32305), .o(delay_add_ln22_unr20_stage8_stallmux_q_28_) );
ao12f80 g777866 ( .a(n_3158), .b(n_3157), .c(n_3156), .o(n_4597) );
na02f80 g774920 ( .a(n_6138), .b(n_5899), .o(n_6168) );
in01f80 g764044 ( .a(FE_OFN780_n_17093), .o(n_17881) );
no02f80 g767665 ( .a(n_46414), .b(n_13173), .o(n_13174) );
na02f80 g772498 ( .a(n_8509), .b(n_8535), .o(n_8536) );
na02f80 g738960 ( .a(n_41209), .b(n_41046), .o(n_41233) );
in01f80 g754470 ( .a(n_25789), .o(n_25822) );
oa22f80 FE_RC_3439_0 ( .a(n_22961), .b(n_22635), .c(n_22580), .d(n_22614), .o(n_22712) );
in01f80 FE_OCP_RBC2835_n_39586 ( .a(n_39586), .o(FE_OCP_RBN2835_n_39586) );
na02f80 FE_RC_2308_0 ( .a(n_25307), .b(n_25741), .o(FE_RN_875_0) );
in01f80 g763925 ( .a(n_17156), .o(n_17157) );
in01f80 g774784 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_19_), .o(n_7344) );
in01f80 FE_RC_218_0 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_3_), .o(FE_RN_72_0) );
no02f80 g738479 ( .a(FE_OCP_RBN2316_n_41420), .b(n_41543), .o(n_41642) );
in01f80 g744107 ( .a(n_35593), .o(n_35646) );
no02f80 g736811 ( .a(n_43067), .b(n_43066), .o(n_43089) );
in01f80 newInst_1938 ( .a(newNet_1373), .o(newNet_1938) );
ao12f80 g774220 ( .a(n_7006), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_15_), .o(n_7187) );
in01f80 newInst_3425 ( .a(newNet_2273), .o(newNet_3425) );
na02f80 g781032 ( .a(cos_out_31), .b(FE_OFN2_n_43918), .o(n_305) );
ao12f80 g751280 ( .a(n_29713), .b(n_29712), .c(n_29711), .o(n_29993) );
no02f80 g758865 ( .a(n_21500), .b(n_21432), .o(n_21679) );
oa12f80 g778938 ( .a(n_2157), .b(n_2158), .c(n_2156), .o(n_2898) );
na02f80 g748682 ( .a(n_31358), .b(n_31077), .o(n_31381) );
no02f80 g761792 ( .a(n_18378), .b(n_18200), .o(n_18438) );
oa12f80 g766777 ( .a(n_13749), .b(n_13748), .c(n_13747), .o(n_15678) );
na02f80 g747252 ( .a(n_32785), .b(n_31181), .o(n_32845) );
in01f80 newInst_3697 ( .a(newNet_3696), .o(newNet_3697) );
in01f80 FE_RC_2378_0 ( .a(n_45659), .o(FE_RN_926_0) );
no02f80 g739342 ( .a(n_45147), .b(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n_40692) );
no02f80 g764522 ( .a(n_16046), .b(n_16004), .o(n_16197) );
ao22s80 FE_RC_3885_0 ( .a(n_45024), .b(n_21194), .c(n_45026), .d(n_21226), .o(n_21361) );
no02f80 g756611 ( .a(FE_OFN745_n_23604), .b(n_23603), .o(n_23629) );
na02f80 g740072 ( .a(n_40069), .b(n_40073), .o(n_40070) );
na02f80 g757651 ( .a(n_22820), .b(n_22708), .o(n_22748) );
no02f80 g765537 ( .a(n_14982), .b(n_13833), .o(n_15112) );
no02f80 g750457 ( .a(FE_OCP_RBN2376_n_29480), .b(FE_OCPN1464_n_29630), .o(n_29531) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_15_ ( .ck(newNet_2487), .d(n_32259), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_) );
oa22f80 FE_RC_253_0 ( .a(FE_OCP_RBN2505_n_13896), .b(n_14763), .c(n_14762), .d(FE_OCP_RBN2503_n_13896), .o(n_14872) );
in01f80 g767267 ( .a(n_13559), .o(n_13570) );
no02f80 g770227 ( .a(n_10709), .b(FE_OCP_RBN3643_n_44490), .o(n_10755) );
in01f80 g767795 ( .a(n_12968), .o(n_12969) );
in01f80 g744351 ( .a(n_46227), .o(n_36855) );
na02f80 g757936 ( .a(n_22852), .b(n_22736), .o(n_22926) );
in01f80 FE_OCP_RBC2635_n_38806 ( .a(n_38806), .o(FE_OCP_RBN2635_n_38806) );
in01f80 g744912 ( .a(n_35092), .o(n_35113) );
in01f80 g774851 ( .a(n_46994), .o(n_6318) );
in01f80 g741925 ( .a(n_38145), .o(n_38170) );
in01f80 g754890 ( .a(n_25721), .o(n_25722) );
in01f80 g769359 ( .a(n_11896), .o(n_11862) );
ao12f80 g775993 ( .a(n_4918), .b(n_5107), .c(n_4821), .o(n_5208) );
in01f80 g775689 ( .a(n_5527), .o(n_5489) );
no02f80 g780621 ( .a(n_679), .b(FE_OFN50_n_1045), .o(n_692) );
no02f80 g740148 ( .a(FE_OCP_RBN3721_n_39913), .b(n_39864), .o(n_40254) );
ao12f80 g764722 ( .a(n_15843), .b(n_16029), .c(n_15934), .o(n_16142) );
na02f80 FE_RC_3500_0 ( .a(n_27355), .b(n_27433), .o(FE_RN_1510_0) );
in01f80 FE_OCP_RBC2794_n_10106 ( .a(n_10106), .o(FE_OCP_RBN2794_n_10106) );
na02f80 g773981 ( .a(n_6809), .b(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_7276) );
na02f80 g749188 ( .a(n_30800), .b(FE_OCPN1862_n_30319), .o(n_30882) );
na02f80 g743330 ( .a(n_37840), .b(n_37839), .o(n_37841) );
no02f80 g750171 ( .a(n_30836), .b(n_30127), .o(n_30952) );
in01f80 g760164 ( .a(n_20435), .o(n_20461) );
oa22f80 FE_RC_935_0 ( .a(n_26290), .b(FE_OCPN1488_n_23447), .c(FE_RN_1667_0), .d(n_26291), .o(n_26442) );
in01f80 newInst_692 ( .a(newNet_482), .o(newNet_692) );
in01f80 g741052 ( .a(n_39504), .o(n_39505) );
na02f80 g746466 ( .a(n_34942), .b(n_44262), .o(n_34964) );
no02f80 g746914 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_18_), .o(n_33181) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_5_ ( .ck(newNet_2054), .d(n_4992), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_) );
na02f80 g739558 ( .a(n_45511), .b(n_40617), .o(n_40639) );
no02f80 g767578 ( .a(n_13470), .b(n_13377), .o(n_13424) );
oa22f80 FE_RC_4107_0 ( .a(n_22459), .b(n_22612), .c(n_22500), .d(n_22598), .o(n_22774) );
na02f80 g746248 ( .a(n_33707), .b(n_33329), .o(n_33729) );
oa12f80 g768514 ( .a(n_12248), .b(n_12334), .c(n_12182), .o(n_12378) );
na02f80 g744744 ( .a(n_35219), .b(FE_OCPN1434_n_30614), .o(n_35264) );
in01f80 g766106 ( .a(n_14582), .o(n_14607) );
na02f80 g743422 ( .a(n_36611), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36653) );
no02f80 g741860 ( .a(n_38383), .b(n_38382), .o(n_38384) );
oa12f80 g765045 ( .a(n_16102), .b(n_15975), .c(n_15874), .o(n_16312) );
no02f80 g758248 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .o(n_23058) );
in01f80 g759822 ( .a(n_21750), .o(n_21721) );
ao22s80 FE_RC_3820_0 ( .a(n_24830), .b(n_24922), .c(n_24831), .d(n_24921), .o(n_25045) );
in01f80 g760603 ( .a(n_19841), .o(n_19857) );
in01f80 g740139 ( .a(n_39845), .o(n_39904) );
na02f80 g761822 ( .a(n_19126), .b(n_18619), .o(n_19194) );
in01f80 g766475 ( .a(n_14149), .o(n_14148) );
no02f80 g779279 ( .a(n_1736), .b(n_1735), .o(n_1737) );
no02f80 g748970 ( .a(n_31098), .b(n_30987), .o(n_31155) );
na02f80 g773195 ( .a(n_7721), .b(n_7923), .o(n_7917) );
ao12f80 g757305 ( .a(n_23462), .b(n_44068), .c(delay_xor_ln21_unr15_stage6_stallmux_q_14_), .o(n_23167) );
in01f80 FE_RC_3305_0 ( .a(FE_RN_1455_0), .o(FE_RN_1452_0) );
oa12f80 g754125 ( .a(FE_OCPN1522_n_26054), .b(n_26055), .c(FE_OCP_RBN2827_FE_RN_1573_0), .o(n_26089) );
no02f80 g738719 ( .a(n_41382), .b(n_41402), .o(n_41460) );
no02f80 g747337 ( .a(n_33842), .b(n_33841), .o(n_33843) );
na02f80 g746476 ( .a(n_34552), .b(n_34587), .o(n_35809) );
ao12f80 g742882 ( .a(n_37082), .b(n_36954), .c(n_36563), .o(n_37083) );
na02f80 g761457 ( .a(n_19647), .b(n_19796), .o(n_19850) );
in01f80 newInst_2401 ( .a(newNet_2400), .o(newNet_2401) );
in01f80 FE_RC_2706_0 ( .a(n_8326), .o(FE_RN_1138_0) );
oa12f80 g765821 ( .a(n_15248), .b(n_15290), .c(n_15247), .o(n_15665) );
no02f80 g768372 ( .a(n_12471), .b(n_12470), .o(n_12472) );
in01f80 g768971 ( .a(n_12193), .o(n_11867) );
in01f80 g751006 ( .a(n_28871), .o(n_28967) );
oa12f80 g757793 ( .a(n_22436), .b(FE_OCP_RBN1920_n_22476), .c(n_22554), .o(n_22573) );
no02f80 g742999 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n_36999) );
in01f80 FE_OCP_RBC3511_n_19599 ( .a(FE_OCP_RBN3510_n_19599), .o(FE_OCP_RBN3511_n_19599) );
oa12f80 g765908 ( .a(n_14348), .b(n_15088), .c(n_14389), .o(n_15290) );
in01f80 g770663 ( .a(n_10225), .o(n_10202) );
oa12f80 g736518 ( .a(n_319), .b(n_43652), .c(FE_OFN2_n_43918), .o(n_43688) );
no02f80 g738571 ( .a(n_41912), .b(n_41828), .o(n_41570) );
no02f80 g776727 ( .a(n_3786), .b(n_3727), .o(n_3787) );
in01f80 newInst_502 ( .a(newNet_501), .o(newNet_502) );
na02f80 g746589 ( .a(n_34666), .b(n_34738), .o(n_34757) );
no02f80 g753299 ( .a(n_27086), .b(n_25823), .o(n_27168) );
in01f80 FE_OCP_RBC1845_n_20910 ( .a(FE_OCP_RBN1843_n_20910), .o(FE_OCP_RBN1845_n_20910) );
in01f80 FE_OCP_RBC2642_n_34921 ( .a(FE_OCP_RBN2641_n_34921), .o(FE_OCP_RBN2642_n_34921) );
na02f80 g779032 ( .a(n_2127), .b(delay_add_ln22_unr2_stage2_stallmux_q_16_), .o(n_2180) );
na02f80 g737026 ( .a(n_43030), .b(n_43132), .o(n_43553) );
na02f80 g778133 ( .a(FE_OCP_RBN2400_n_2885), .b(n_2823), .o(n_2957) );
in01f80 g752792 ( .a(n_28214), .o(n_28215) );
in01f80 FE_OCP_RBC1993_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_ ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .o(FE_OCP_RBN1993_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
no02f80 g737701 ( .a(n_42203), .b(n_41796), .o(n_42287) );
in01f80 g770814 ( .a(n_10025), .o(n_10026) );
oa12f80 g745250 ( .a(n_35657), .b(n_35656), .c(FE_OFN221_n_35655), .o(n_35726) );
oa22f80 g749011 ( .a(n_32249), .b(n_31574), .c(n_32250), .d(n_31573), .o(n_32294) );
oa22f80 FE_RC_2626_0 ( .a(FE_OCP_RBN3382_n_12365), .b(n_12110), .c(n_12111), .d(n_12365), .o(n_12453) );
in01f80 g752056 ( .a(n_28186), .o(n_28141) );
na02f80 g759505 ( .a(FE_OCP_RBN1217_n_20595), .b(n_20470), .o(n_20619) );
no02f80 FE_RC_2667_0 ( .a(FE_RN_1114_0), .b(n_4111), .o(n_4233) );
oa12f80 g738325 ( .a(n_41445), .b(n_41818), .c(n_41760), .o(n_41833) );
in01f80 g773372 ( .a(FE_OCP_RBN2229_n_7598), .o(n_7721) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_11_ ( .ck(newNet_272), .d(n_46150), .o(delay_xor_ln22_unr6_stage3_stallmux_q_11_) );
in01f80 g762053 ( .a(n_18629), .o(n_18630) );
no02f80 g769959 ( .a(n_10994), .b(n_11047), .o(n_11072) );
ao12f80 g741482 ( .a(n_38776), .b(n_38775), .c(n_38774), .o(n_39740) );
in01f80 g765968 ( .a(n_15088), .o(n_15089) );
ao22s80 g736427 ( .a(n_43754), .b(n_43584), .c(n_43755), .d(n_43583), .o(n_43795) );
in01f80 g750950 ( .a(n_30105), .o(n_30068) );
in01f80 FE_OCP_RBC3120_n_27655 ( .a(n_27655), .o(FE_OCP_RBN3120_n_27655) );
na02f80 g759522 ( .a(n_20426), .b(n_20850), .o(n_20913) );
in01f80 g765362 ( .a(n_15569), .o(n_16341) );
oa22f80 g749566 ( .a(n_31692), .b(n_31532), .c(n_31693), .d(n_31533), .o(n_31779) );
no02f80 g737965 ( .a(n_42182), .b(n_41369), .o(n_42234) );
no02f80 g777321 ( .a(n_3951), .b(n_4207), .o(n_4371) );
no02f80 g769821 ( .a(n_11052), .b(n_44463), .o(n_11053) );
in01f80 FE_RC_3717_0 ( .a(n_5911), .o(FE_RN_1635_0) );
oa22f80 g756957 ( .a(n_23743), .b(n_22811), .c(n_23803), .d(n_22885), .o(n_24075) );
in01f80 newInst_322 ( .a(newNet_280), .o(newNet_322) );
in01f80 g762462 ( .a(n_18130), .o(n_18087) );
in01f80 g778629 ( .a(n_2900), .o(n_2954) );
na02f80 g749357 ( .a(n_30543), .b(n_30584), .o(n_30585) );
no02f80 g769206 ( .a(n_11796), .b(n_11795), .o(n_12264) );
in01f80 newInst_3332 ( .a(newNet_3331), .o(newNet_3332) );
in01f80 g737837 ( .a(n_42285), .o(n_42394) );
na02f80 g779788 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_), .o(n_1462) );
in01f80 g768815 ( .a(n_11952), .o(n_11953) );
in01f80 newInst_837 ( .a(newNet_836), .o(newNet_837) );
no02f80 g765051 ( .a(n_15525), .b(n_44051), .o(n_15604) );
na02f80 g760669 ( .a(n_19746), .b(n_19745), .o(n_19856) );
oa22f80 g740344 ( .a(n_39790), .b(n_39778), .c(n_39791), .d(n_39755), .o(n_39855) );
ao12f80 g780777 ( .a(n_535), .b(n_534), .c(n_533), .o(n_665) );
in01f80 newInst_2690 ( .a(newNet_298), .o(newNet_2690) );
in01f80 g754211 ( .a(n_25972), .o(n_25994) );
in01f80 g746540 ( .a(n_34841), .o(n_34842) );
in01f80 g749702 ( .a(n_31635), .o(n_31636) );
no02f80 g772899 ( .a(n_7887), .b(n_7722), .o(n_7959) );
na02f80 g764584 ( .a(n_16144), .b(FE_OCPN1734_n_16143), .o(n_16181) );
no02f80 g756737 ( .a(n_23441), .b(n_23143), .o(n_23464) );
no02f80 g746706 ( .a(n_33039), .b(n_33025), .o(n_33026) );
na02f80 g743305 ( .a(n_36712), .b(n_36677), .o(n_36725) );
no02f80 g768069 ( .a(n_12753), .b(n_12671), .o(n_12700) );
na02f80 g779268 ( .a(n_1813), .b(n_1520), .o(n_1853) );
no02f80 g773101 ( .a(n_7783), .b(n_7782), .o(n_7975) );
na02f80 g738406 ( .a(n_41731), .b(n_41701), .o(n_42054) );
in01f80 g740442 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_), .o(n_39737) );
na02f80 g771287 ( .a(n_9786), .b(n_9722), .o(n_9885) );
in01f80 FE_OCP_RBC3730_n_31819 ( .a(FE_OCP_RBN3085_n_31819), .o(FE_OCP_RBN3730_n_31819) );
no02f80 g752802 ( .a(n_28106), .b(n_28105), .o(n_28666) );
na02f80 g761723 ( .a(n_19339), .b(n_18910), .o(n_19405) );
na03f80 FE_RC_1291_0 ( .a(n_33833), .b(n_33733), .c(n_33785), .o(n_33906) );
in01f80 g756045 ( .a(n_25163), .o(n_25164) );
in01f80 newInst_3554 ( .a(newNet_568), .o(newNet_3554) );
na02f80 g765964 ( .a(n_14692), .b(n_14678), .o(n_14752) );
in01f80 newInst_3121 ( .a(newNet_3120), .o(newNet_3121) );
in01f80 newInst_3646 ( .a(newNet_3645), .o(newNet_3646) );
in01f80 newInst_38 ( .a(newNet_34), .o(newNet_38) );
no02f80 g779349 ( .a(FE_OCP_RBN2158_n_1614), .b(n_1425), .o(n_1672) );
oa22f80 FE_RC_3371_0 ( .a(n_22961), .b(n_22789), .c(n_22580), .d(n_22739), .o(n_22815) );
in01f80 g759401 ( .a(n_20857), .o(n_20858) );
in01f80 FE_OCP_RBC2612_n_9075 ( .a(n_9075), .o(FE_OCP_RBN2612_n_9075) );
na02f80 g745629 ( .a(n_35462), .b(n_34938), .o(n_35509) );
no02f80 g770615 ( .a(n_10198), .b(FE_OCP_RBN3599_FE_OCPN1243_n_44460), .o(n_10201) );
in01f80 g738071 ( .a(n_42122), .o(n_42139) );
in01f80 g741883 ( .a(n_38468), .o(n_38405) );
ao12f80 g737494 ( .a(n_42377), .b(n_42541), .c(n_42540), .o(n_42552) );
na02f80 g737330 ( .a(n_42831), .b(n_42329), .o(n_42869) );
no04s80 g752055 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_10_), .b(delay_xor_ln21_unr18_stage7_stallmux_q_9_), .c(n_28032), .d(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .o(n_28070) );
ao12f80 g737524 ( .a(n_42203), .b(n_42337), .c(n_42242), .o(n_42381) );
no02f80 g759905 ( .a(n_21374), .b(n_21720), .o(n_21751) );
ao12f80 g775067 ( .a(n_6080), .b(n_6012), .c(n_6039), .o(n_6081) );
in01f80 g746737 ( .a(n_33234), .o(n_33219) );
in01f80 g756293 ( .a(n_24098), .o(n_24093) );
no02f80 g744154 ( .a(n_35575), .b(n_35533), .o(n_35834) );
in01f80 g748865 ( .a(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37709) );
in01f80 FE_RC_635_0 ( .a(n_6876), .o(FE_RN_198_0) );
na02f80 g753165 ( .a(n_27340), .b(n_27383), .o(n_27480) );
oa22f80 g779890 ( .a(n_44652), .b(n_1134), .c(n_44623), .d(n_1120), .o(n_1324) );
ao22s80 FE_RC_1011_0 ( .a(n_12688), .b(n_12527), .c(n_12689), .d(n_12526), .o(n_12800) );
in01f80 g759432 ( .a(n_20997), .o(n_21069) );
no02f80 g756874 ( .a(n_24150), .b(n_24059), .o(n_24354) );
in01f80 FE_OCP_RBC3052_n_39913 ( .a(n_39913), .o(FE_OCP_RBN3052_n_39913) );
in01f80 FE_OCPC969_n_19342 ( .a(FE_OCPN967_n_19342), .o(FE_OCPN969_n_19342) );
in01f80 g776010 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_8_), .o(n_5104) );
na02f80 g751273 ( .a(n_29744), .b(n_29249), .o(n_29783) );
na02f80 g761533 ( .a(n_18719), .b(n_18554), .o(n_18829) );
no02f80 g750276 ( .a(n_29773), .b(FE_OCP_DRV_N1566_n_28654), .o(n_29787) );
in01f80 FE_RC_3984_0 ( .a(n_14503), .o(FE_RN_1727_0) );
na02f80 g741180 ( .a(FE_OCP_RBN2638_n_38806), .b(n_38884), .o(n_38921) );
in01f80 g748022 ( .a(n_31881), .o(n_31882) );
in01f80 g751254 ( .a(n_29837), .o(n_29909) );
in01f80 g753153 ( .a(n_27525), .o(n_27526) );
in01f80 g777249 ( .a(n_3616), .o(n_3610) );
no02f80 FE_RC_3487_0 ( .a(FE_RN_1503_0), .b(FE_RN_1501_0), .o(FE_RN_1502_0) );
na02f80 g767270 ( .a(n_13430), .b(FE_OCP_RBN3428_n_12890), .o(n_13458) );
no02f80 g762922 ( .a(n_17679), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_6_), .o(n_17718) );
na02f80 g761672 ( .a(n_18889), .b(n_18916), .o(n_20345) );
oa22f80 g771099 ( .a(FE_OCP_RBN2721_n_9494), .b(FE_OCPN903_n_44581), .c(n_9494), .d(FE_OCP_RBN2619_n_44561), .o(n_9666) );
oa12f80 g784068 ( .a(n_1111), .b(n_45808), .c(n_936), .o(n_45814) );
ao12f80 g746334 ( .a(n_33562), .b(n_33561), .c(n_33560), .o(n_34160) );
na02f80 g743438 ( .a(n_37750), .b(n_37749), .o(n_37751) );
oa22f80 FE_RC_1231_0 ( .a(n_17336), .b(n_44447), .c(n_16339), .d(n_17729), .o(n_17808) );
in01f80 g764162 ( .a(n_16565), .o(n_16557) );
in01f80 g773813 ( .a(n_7166), .o(n_7167) );
in01f80 newInst_2185 ( .a(newNet_1693), .o(newNet_2185) );
in01f80 FE_RC_3682_0 ( .a(n_23107), .o(FE_RN_1617_0) );
in01f80 g746840 ( .a(n_33287), .o(n_33288) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_2_ ( .ck(newNet_3291), .d(n_31051), .o(delay_add_ln22_unr20_stage8_stallmux_q_2_) );
in01f80 g758831 ( .a(n_21786), .o(n_21804) );
in01f80 g748933 ( .a(n_31156), .o(n_31157) );
in01f80 g749876 ( .a(n_31409), .o(n_31338) );
no02f80 g759076 ( .a(n_21131), .b(n_20667), .o(n_21196) );
oa12f80 g755309 ( .a(n_24822), .b(n_24897), .c(n_24776), .o(n_24974) );
ao12f80 g759478 ( .a(n_20654), .b(n_20442), .c(FE_OCP_RBN1216_n_20595), .o(n_20693) );
in01f80 FE_OCP_RBC1713_FE_RN_664_0 ( .a(FE_RN_664_0), .o(FE_OCP_RBN1713_FE_RN_664_0) );
in01f80 g764536 ( .a(n_16011), .o(n_16050) );
in01f80 FE_OCPC965_n_47020 ( .a(n_47020), .o(FE_OCPN965_n_47020) );
in01f80 g755720 ( .a(n_24518), .o(n_24546) );
no02f80 g773951 ( .a(n_6970), .b(n_6984), .o(n_6971) );
no02f80 g757977 ( .a(n_22028), .b(FE_OCPN1502_n_20723), .o(n_22029) );
in01f80 g772901 ( .a(n_7948), .o(n_7967) );
no02f80 g756170 ( .a(n_24175), .b(n_21852), .o(n_24202) );
ao12f80 g779090 ( .a(n_2052), .b(n_2051), .c(n_2050), .o(n_2104) );
no02f80 g742647 ( .a(n_37852), .b(n_37849), .o(n_37901) );
in01f80 g763566 ( .a(n_16836), .o(n_16923) );
na02f80 g740435 ( .a(n_39726), .b(n_39724), .o(n_39750) );
no02f80 g741031 ( .a(n_39155), .b(n_39154), .o(n_39156) );
in01f80 g774407 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_4_), .o(n_6504) );
na02f80 g778596 ( .a(n_2825), .b(n_2758), .o(n_3314) );
ao12f80 g764808 ( .a(n_46419), .b(n_15588), .c(n_15182), .o(n_15655) );
no02f80 g778281 ( .a(n_3857), .b(n_2988), .o(n_2989) );
no03m80 g747323 ( .a(n_32595), .b(n_32522), .c(n_32599), .o(n_32596) );
oa22f80 FE_RC_3131_0 ( .a(n_31234), .b(n_31463), .c(FE_RN_786_0), .d(FE_RN_787_0), .o(n_31677) );
in01f80 newInst_1630 ( .a(newNet_1629), .o(newNet_1630) );
oa12f80 g736444 ( .a(n_43527), .b(n_43716), .c(n_43331), .o(n_43777) );
in01f80 g764784 ( .a(n_15795), .o(n_15796) );
no02f80 g738138 ( .a(n_42029), .b(n_41708), .o(n_42059) );
in01f80 g780631 ( .a(n_887), .o(n_891) );
in01f80 g757448 ( .a(n_23461), .o(n_23032) );
in01f80 newInst_2180 ( .a(newNet_2179), .o(newNet_2180) );
in01f80 newInst_2130 ( .a(newNet_1793), .o(newNet_2130) );
no02f80 g756942 ( .a(n_24149), .b(n_24037), .o(n_24189) );
in01f80 g761665 ( .a(n_18858), .o(n_18890) );
na02f80 g756780 ( .a(n_24153), .b(n_24105), .o(n_24154) );
na02f80 g775191 ( .a(n_5958), .b(n_5689), .o(n_6023) );
ao22s80 FE_RC_18_0 ( .a(n_5178), .b(n_3734), .c(n_3380), .d(n_3637), .o(n_3805) );
na02f80 FE_RC_2276_0 ( .a(FE_RN_846_0), .b(FE_RN_848_0), .o(FE_RN_849_0) );
na02f80 FE_RC_2893_0 ( .a(n_39869), .b(n_39843), .o(FE_RN_1253_0) );
oa12f80 g760847 ( .a(n_19510), .b(FE_OCP_RBN3841_n_19419), .c(n_19508), .o(n_19626) );
in01f80 g773200 ( .a(n_7916), .o(n_7980) );
oa22f80 FE_RC_1678_0 ( .a(n_8819), .b(n_7606), .c(n_7605), .d(n_8863), .o(n_8923) );
in01f80 g773137 ( .a(n_8018), .o(n_8085) );
na02f80 g765575 ( .a(n_15142), .b(n_14464), .o(n_15448) );
no02f80 g777316 ( .a(n_3604), .b(n_2360), .o(n_3756) );
in01f80 g771611 ( .a(n_10383), .o(n_10384) );
in01f80 newInst_7 ( .a(newNet_6), .o(newNet_7) );
in01f80 FE_OCPC1859_n_35415 ( .a(n_35415), .o(FE_OCPN1859_n_35415) );
in01f80 g777684 ( .a(n_3372), .o(n_3393) );
in01f80 g779438 ( .a(n_1563), .o(n_1564) );
ao12f80 g754581 ( .a(n_25370), .b(n_26163), .c(n_25372), .o(n_26233) );
in01f80 g764281 ( .a(n_16405), .o(n_16406) );
in01f80 newInst_509 ( .a(newNet_508), .o(newNet_509) );
na03f80 FE_RC_3765_0 ( .a(FE_OCP_RBN3401_n_37670), .b(FE_OCP_RBN2211_n_37720), .c(n_37698), .o(n_37763) );
no02f80 g773090 ( .a(n_7962), .b(n_8085), .o(n_8772) );
in01f80 FE_OCP_RBC2591_n_14460 ( .a(n_14460), .o(FE_OCP_RBN2591_n_14460) );
na02f80 g771868 ( .a(n_9480), .b(n_9505), .o(n_10086) );
in01f80 g758905 ( .a(n_21759), .o(n_21760) );
ao12f80 g775639 ( .a(n_4956), .b(n_5031), .c(n_4966), .o(n_5138) );
in01f80 g740127 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_2_), .o(n_40667) );
no02f80 g750742 ( .a(n_29318), .b(n_29317), .o(n_29340) );
in01f80 g741286 ( .a(n_38909), .o(n_39044) );
in01f80 g764816 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_7_), .o(n_17800) );
na02f80 g773414 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_31_), .o(n_7535) );
oa12f80 g739385 ( .a(n_45181), .b(delay_add_ln22_unr27_stage10_stallmux_q_17_), .c(delay_add_ln22_unr27_stage10_stallmux_q_16_), .o(n_40869) );
no02f80 g747818 ( .a(n_33238), .b(n_33370), .o(n_33313) );
in01f80 g757293 ( .a(n_23023), .o(n_23003) );
in01f80 g743364 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_), .o(n_36636) );
na02f80 g773902 ( .a(n_7060), .b(n_6968), .o(n_7061) );
no02f80 g755815 ( .a(n_24442), .b(n_24394), .o(n_24492) );
ao12f80 g755938 ( .a(n_24909), .b(n_24908), .c(n_24907), .o(n_25259) );
in01f80 g762693 ( .a(n_18016), .o(n_18017) );
oa12f80 g737456 ( .a(n_42663), .b(n_42637), .c(n_42583), .o(n_42687) );
na02f80 FE_RC_1860_0 ( .a(n_13634), .b(n_13858), .o(FE_RN_570_0) );
ao22s80 g777677 ( .a(n_3385), .b(n_2913), .c(n_4228), .d(n_2759), .o(n_3481) );
no02f80 g736656 ( .a(n_43332), .b(n_43369), .o(n_43411) );
in01f80 FE_OCP_RBC3537_n_8597 ( .a(n_8597), .o(FE_OCP_RBN3537_n_8597) );
na02f80 g779735 ( .a(n_1379), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_0_), .o(n_1407) );
in01f80 g762220 ( .a(n_18731), .o(n_18814) );
in01f80 g764051 ( .a(n_17093), .o(n_17732) );
no02f80 g750915 ( .a(n_30333), .b(n_30305), .o(n_31294) );
na02f80 g766110 ( .a(n_14634), .b(n_14605), .o(n_14635) );
no02f80 g759788 ( .a(n_21749), .b(n_21748), .o(n_21776) );
na02f80 g765182 ( .a(n_16344), .b(FE_OCP_RBN1924_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_16345) );
no02f80 g774506 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n_6756) );
in01f80 FE_OCP_RBC3489_n_3390 ( .a(FE_OCP_RBN3488_n_3390), .o(FE_OCP_RBN3489_n_3390) );
in01f80 g780213 ( .a(n_1125), .o(n_1144) );
in01f80 g752989 ( .a(n_27353), .o(n_27354) );
in01f80 newInst_2508 ( .a(newNet_2507), .o(newNet_2508) );
ao12f80 g741938 ( .a(n_37990), .b(n_37991), .c(n_37989), .o(n_38067) );
na02f80 g736748 ( .a(n_43430), .b(n_43429), .o(n_43465) );
na02f80 g778587 ( .a(n_2325), .b(n_2306), .o(n_2307) );
in01f80 g771389 ( .a(n_9698), .o(n_9699) );
oa22f80 g758628 ( .a(n_21767), .b(n_21843), .c(n_21766), .d(n_21844), .o(n_21920) );
no02f80 g777634 ( .a(n_3393), .b(n_3154), .o(n_3394) );
in01f80 FE_OCP_RBC3635_n_47260 ( .a(FE_OCP_RBN3634_n_47260), .o(FE_OCP_RBN3635_n_47260) );
na02f80 g766269 ( .a(n_14326), .b(FE_OCP_RBN2459_n_13765), .o(n_14374) );
na02f80 g754007 ( .a(n_26129), .b(n_26083), .o(n_26131) );
na02f80 g754916 ( .a(n_25270), .b(n_24438), .o(n_25485) );
no02f80 g766741 ( .a(n_13725), .b(n_13724), .o(n_13813) );
in01f80 newInst_1197 ( .a(newNet_1196), .o(newNet_1197) );
no02f80 g740790 ( .a(n_39510), .b(n_39509), .o(n_39511) );
in01f80 g780604 ( .a(n_710), .o(n_711) );
in01f80 g742398 ( .a(n_37763), .o(n_37775) );
no02f80 g750931 ( .a(n_28976), .b(n_28653), .o(n_28997) );
no02f80 g764906 ( .a(n_15503), .b(n_15474), .o(n_15623) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_26_ ( .ck(newNet_1978), .d(n_12117), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_26_) );
na02f80 g750851 ( .a(n_29055), .b(FE_RN_1513_0), .o(n_29094) );
in01f80 g780495 ( .a(n_982), .o(n_983) );
na02f80 g754946 ( .a(n_25187), .b(n_25157), .o(n_25158) );
ao12f80 g742696 ( .a(n_37324), .b(n_37323), .c(n_37322), .o(n_37871) );
in01f80 g746296 ( .a(n_33567), .o(n_33584) );
in01f80 g742154 ( .a(n_38197), .o(n_38198) );
in01f80 newInst_1336 ( .a(newNet_263), .o(newNet_1336) );
ao22s80 FE_RC_1351_0 ( .a(n_43609), .b(n_43893), .c(n_43610), .d(n_43892), .o(n_43911) );
na02f80 g750478 ( .a(n_29546), .b(n_29527), .o(n_29547) );
in01f80 g765260 ( .a(n_15376), .o(n_15377) );
in01f80 g765845 ( .a(n_15287), .o(n_15288) );
in01f80 g736508 ( .a(n_43714), .o(n_43715) );
oa12f80 g752020 ( .a(n_28730), .b(n_28729), .c(n_28728), .o(n_29076) );
no02f80 g754412 ( .a(n_25677), .b(n_25378), .o(n_25734) );
ao22s80 FE_RC_1380_0 ( .a(n_20784), .b(n_21165), .c(n_20785), .d(n_21196), .o(n_21358) );
no02f80 g774036 ( .a(n_6848), .b(n_6910), .o(n_6974) );
na02f80 g750955 ( .a(n_28935), .b(n_28652), .o(n_28950) );
oa22f80 FE_RC_4265_0 ( .a(n_17783), .b(FE_OCP_RBN1340_n_19077), .c(n_17900), .d(n_19077), .o(n_19278) );
ao12f80 g741892 ( .a(n_37907), .b(n_38358), .c(n_38267), .o(n_38410) );
in01f80 FE_OCP_DRV_C1597_n_35644 ( .a(n_35644), .o(FE_OCP_DRV_N1597_n_35644) );
no02f80 FE_RC_1519_0 ( .a(FE_RN_426_0), .b(FE_RN_427_0), .o(FE_RN_428_0) );
no02f80 g742491 ( .a(n_37577), .b(n_37709), .o(n_37646) );
na02f80 g768305 ( .a(n_12607), .b(n_12606), .o(n_12608) );
no03m80 FE_RC_480_0 ( .a(n_23462), .b(FE_RN_143_0), .c(n_23460), .o(n_23465) );
in01f80 g780276 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_10_), .o(n_1011) );
oa12f80 g743935 ( .a(n_35529), .b(n_35593), .c(FE_OCP_RBN2885_n_35517), .o(n_35710) );
na02f80 g757778 ( .a(n_23089), .b(n_22657), .o(n_23090) );
na02f80 g744240 ( .a(n_46219), .b(n_36820), .o(n_37259) );
in01f80 g761894 ( .a(n_19650), .o(n_19051) );
in01f80 FE_OCP_RBC2801_n_15706 ( .a(FE_OCP_RBN2800_n_15706), .o(FE_OCP_RBN2801_n_15706) );
no02f80 g740984 ( .a(n_39209), .b(n_39095), .o(n_39235) );
in01f80 newInst_295 ( .a(newNet_294), .o(newNet_295) );
no02f80 g775035 ( .a(n_5977), .b(n_4675), .o(n_6089) );
in01f80 g737866 ( .a(n_42480), .o(n_42481) );
no02f80 g751765 ( .a(n_28268), .b(n_28166), .o(n_28303) );
no02f80 g754538 ( .a(n_26602), .b(n_26636), .o(n_26685) );
in01f80 FE_OCPC3786_n_22156 ( .a(n_22156), .o(FE_OCPN3786_n_22156) );
na02f80 g760706 ( .a(n_19666), .b(FE_OCP_DRV_N1564_n_19665), .o(n_19701) );
in01f80 g751078 ( .a(n_28933), .o(n_28890) );
no02f80 g741982 ( .a(n_38121), .b(n_38057), .o(n_38058) );
na02f80 g784761 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .o(n_47247) );
na02f80 g759531 ( .a(n_20817), .b(n_20796), .o(n_20910) );
no02f80 g773131 ( .a(FE_OCP_RBN3461_n_7886), .b(n_7915), .o(n_8058) );
no02f80 g746786 ( .a(n_33259), .b(n_33323), .o(n_33324) );
in01f80 g768039 ( .a(n_13162), .o(n_13249) );
in01f80 newInst_3066 ( .a(newNet_3065), .o(newNet_3066) );
na02f80 g738578 ( .a(n_41877), .b(n_41901), .o(n_41986) );
na02f80 g741132 ( .a(n_39045), .b(n_39044), .o(n_39074) );
no02f80 g737381 ( .a(n_42811), .b(n_42415), .o(n_42833) );
no02f80 g774586 ( .a(FE_OCP_RBN1990_delay_xor_ln23_unr6_stage3_stallmux_q), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6517) );
in01f80 g763332 ( .a(n_17233), .o(n_17225) );
in01f80 g762771 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_14_), .o(n_17875) );
in01f80 FE_OCP_RBC3310_n_44722 ( .a(n_44722), .o(FE_OCP_RBN3310_n_44722) );
no02f80 g766941 ( .a(n_13823), .b(n_13939), .o(n_13941) );
no02f80 g755524 ( .a(n_25172), .b(n_24995), .o(n_25224) );
in01f80 FE_OCP_RBC3618_n_14841 ( .a(n_14841), .o(FE_OCP_RBN3618_n_14841) );
ao12f80 g748779 ( .a(n_32376), .b(n_32423), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_32539) );
na02f80 g777769 ( .a(n_3291), .b(n_2840), .o(n_3326) );
ao12f80 g742806 ( .a(n_37105), .b(n_37297), .c(n_37045), .o(n_37346) );
no02f80 g775446 ( .a(n_5651), .b(n_4556), .o(n_5679) );
in01f80 g771131 ( .a(n_9624), .o(n_9636) );
no02f80 g742098 ( .a(n_37937), .b(n_38003), .o(n_38004) );
na02f80 g759415 ( .a(n_20967), .b(n_20995), .o(n_21116) );
in01f80 g770959 ( .a(n_10127), .o(n_10128) );
oa12f80 g765029 ( .a(n_15534), .b(n_15533), .c(n_15532), .o(n_15605) );
no02f80 FE_RC_1880_0 ( .a(FE_RN_582_0), .b(FE_OCP_RBN1091_n_45224), .o(FE_RN_584_0) );
na02f80 g744884 ( .a(n_34955), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35059) );
na02f80 g749961 ( .a(n_29833), .b(n_29872), .o(n_30023) );
in01f80 g762097 ( .a(n_18276), .o(n_18277) );
in01f80 newInst_512 ( .a(newNet_511), .o(newNet_512) );
in01f80 newInst_2551 ( .a(newNet_1345), .o(newNet_2551) );
in01f80 g757245 ( .a(n_23210), .o(n_23211) );
na02f80 g777922 ( .a(n_3097), .b(n_3107), .o(n_4211) );
no02f80 g743023 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_29_), .o(n_36938) );
ao12f80 g777820 ( .a(n_3229), .b(n_3228), .c(n_2712), .o(n_3281) );
in01f80 g746304 ( .a(n_33508), .o(n_33529) );
no02f80 g747807 ( .a(n_33372), .b(n_33626), .o(n_33950) );
na02f80 g751972 ( .a(n_28897), .b(n_28665), .o(n_29045) );
na02f80 g756230 ( .a(n_24056), .b(n_23662), .o(n_24071) );
na02f80 g781344 ( .a(n_110), .b(beta_31), .o(n_107) );
in01f80 g773731 ( .a(n_7227), .o(n_7228) );
na02f80 g774485 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_), .o(n_6667) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_15_ ( .ck(newNet_3162), .d(n_40469), .o(delay_add_ln22_unr27_stage10_stallmux_q_15_) );
in01f80 g741075 ( .a(n_39366), .o(n_39367) );
in01f80 FE_RC_4014_0 ( .a(FE_RN_1743_0), .o(n_15392) );
no02f80 g740337 ( .a(n_40057), .b(n_40303), .o(n_40407) );
na02f80 g740868 ( .a(n_39460), .b(n_40177), .o(n_39461) );
in01f80 newInst_1923 ( .a(newNet_1922), .o(newNet_1923) );
in01f80 g755170 ( .a(n_25046), .o(n_25047) );
in01f80 g750930 ( .a(n_28997), .o(n_28998) );
in01f80 g766479 ( .a(n_14069), .o(n_14098) );
in01f80 FE_OCP_RBC1696_n_19206 ( .a(FE_OCP_RBN1695_n_19206), .o(FE_OCP_RBN1696_n_19206) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_11_ ( .ck(newNet_2420), .d(n_36389), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_) );
na02f80 g738559 ( .a(n_41661), .b(n_41525), .o(n_41740) );
oa12f80 g747861 ( .a(n_33129), .b(n_33128), .c(n_33127), .o(n_33743) );
in01f80 FE_OCPC929_n_44083 ( .a(n_44083), .o(FE_OCPN929_n_44083) );
no02f80 g774248 ( .a(n_6715), .b(n_6544), .o(n_6710) );
oa12f80 g759378 ( .a(n_21001), .b(n_21000), .c(n_20999), .o(n_21066) );
in01f80 newInst_1123 ( .a(newNet_496), .o(newNet_1123) );
in01f80 newInst_688 ( .a(newNet_531), .o(newNet_688) );
na02f80 g773856 ( .a(n_7088), .b(n_6992), .o(n_7089) );
no02f80 g765385 ( .a(FE_OCP_RBN3622_n_15135), .b(n_14276), .o(n_15810) );
oa12f80 g781003 ( .a(n_269), .b(n_263), .c(n_88), .o(n_281) );
in01f80 g770607 ( .a(n_10286), .o(n_10287) );
no02f80 g743062 ( .a(n_37094), .b(n_36949), .o(n_37142) );
in01f80 g742473 ( .a(n_37732), .o(n_37733) );
ao22s80 FE_RC_1359_0 ( .a(n_43635), .b(n_43842), .c(n_43634), .d(n_43843), .o(n_43866) );
na02f80 g746622 ( .a(n_34473), .b(n_34582), .o(n_34606) );
no02f80 g748088 ( .a(n_32023), .b(n_32022), .o(n_32078) );
in01f80 FE_OCPC3764_FE_OCP_RBN2222_n_13010 ( .a(FE_OCP_RBN2222_n_13010), .o(FE_OCPN3764_FE_OCP_RBN2222_n_13010) );
in01f80 FE_OCP_RBC2971_n_31239 ( .a(n_31239), .o(FE_OCP_RBN2971_n_31239) );
na02f80 g771437 ( .a(n_9082), .b(n_8309), .o(n_9140) );
in01f80 g742779 ( .a(n_37353), .o(n_37409) );
in01f80 g745017 ( .a(n_34971), .o(n_34994) );
na02f80 g766262 ( .a(n_14362), .b(n_13515), .o(n_14411) );
no02f80 g779152 ( .a(n_1915), .b(delay_add_ln22_unr2_stage2_stallmux_q_11_), .o(n_1936) );
na02f80 g762919 ( .a(n_17994), .b(n_17992), .o(n_17993) );
in01f80 g770466 ( .a(n_10579), .o(n_10864) );
no02f80 FE_RC_1504_0 ( .a(n_20821), .b(n_20396), .o(FE_RN_421_0) );
in01f80 FE_RC_1834_0 ( .a(FE_OCP_RBN1170_n_13756), .o(FE_RN_552_0) );
no02f80 g749246 ( .a(n_30765), .b(n_30318), .o(n_30806) );
ao12f80 g775850 ( .a(n_5229), .b(n_5283), .c(n_5228), .o(n_5350) );
na02f80 g773709 ( .a(n_7284), .b(n_7107), .o(n_7275) );
in01f80 FE_RC_3687_0 ( .a(n_12394), .o(FE_RN_1620_0) );
in01f80 newInst_2453 ( .a(newNet_2452), .o(newNet_2453) );
oa12f80 g756392 ( .a(n_23695), .b(n_23694), .c(n_23693), .o(n_25064) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_5_ ( .ck(newNet_3587), .d(n_15605), .o(delay_add_ln22_unr11_stage5_stallmux_q_5_) );
no02f80 g742711 ( .a(n_37444), .b(n_37445), .o(n_37483) );
in01f80 g764894 ( .a(n_15588), .o(n_15589) );
no02f80 g746820 ( .a(n_32963), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n_32960) );
na02f80 g745858 ( .a(n_35354), .b(n_34844), .o(n_35390) );
na02f80 g767606 ( .a(n_13326), .b(n_13381), .o(n_13470) );
na02f80 g756462 ( .a(n_23711), .b(n_23734), .o(n_23769) );
no02f80 g759237 ( .a(n_20947), .b(n_20607), .o(n_21018) );
ao22s80 FE_RC_4201_0 ( .a(n_34005), .b(n_34084), .c(n_34004), .d(n_34083), .o(n_34183) );
na02f80 g751739 ( .a(n_28322), .b(n_28311), .o(n_28312) );
no02f80 g762001 ( .a(n_18911), .b(n_18587), .o(n_18966) );
oa12f80 g776392 ( .a(n_4615), .b(n_4614), .c(n_4619), .o(n_4679) );
in01f80 newInst_153 ( .a(newNet_152), .o(newNet_153) );
no02f80 g737487 ( .a(n_42685), .b(n_42665), .o(n_43061) );
oa12f80 g751206 ( .a(n_29837), .b(n_29935), .c(n_29408), .o(n_29936) );
ao22s80 FE_RC_611_0 ( .a(n_40139), .b(n_40521), .c(n_40140), .d(n_40531), .o(n_40568) );
na02f80 g767898 ( .a(n_13116), .b(n_13017), .o(n_13168) );
na02f80 g779280 ( .a(n_1736), .b(n_1557), .o(n_1806) );
in01f80 newInst_2449 ( .a(newNet_2222), .o(newNet_2449) );
na02f80 g776026 ( .a(n_4726), .b(FE_OCP_RBN2723_n_4219), .o(n_4807) );
na02f80 g755993 ( .a(n_24204), .b(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24228) );
no02f80 g742146 ( .a(n_37900), .b(n_37391), .o(n_38062) );
na02f80 g776730 ( .a(n_4332), .b(n_4404), .o(n_4518) );
oa22f80 FE_RC_1455_0 ( .a(n_17336), .b(n_17782), .c(n_16339), .d(n_17756), .o(n_17829) );
no02f80 g784398 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n_46210) );
in01f80 g757042 ( .a(n_23932), .o(n_23933) );
in01f80 g763203 ( .a(n_17481), .o(n_17397) );
in01f80 g777179 ( .a(n_5380), .o(n_5381) );
no02f80 g740387 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39878), .o(n_40273) );
na02f80 g756385 ( .a(n_24012), .b(n_24052), .o(n_24053) );
na02f80 FE_RC_4240_0 ( .a(n_21489), .b(n_21786), .o(FE_RN_1863_0) );
oa12f80 g739899 ( .a(n_40309), .b(FE_OCP_RBN3046_n_40231), .c(n_40238), .o(n_40377) );
in01f80 g740106 ( .a(n_40281), .o(n_40282) );
oa22f80 g756252 ( .a(FE_OCPN3164_n_24117), .b(n_22767), .c(n_24116), .d(n_24119), .o(n_26090) );
na02f80 g769379 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_11935) );
in01f80 newInst_1696 ( .a(newNet_711), .o(newNet_1696) );
no02f80 g769681 ( .a(FE_OCP_RBN3706_n_11146), .b(n_44498), .o(n_11183) );
no02f80 g738386 ( .a(n_41642), .b(n_41588), .o(n_41643) );
no02f80 g744606 ( .a(n_35316), .b(n_35315), .o(n_35363) );
in01f80 g749999 ( .a(FE_OCP_RBN3012_n_31117), .o(n_31311) );
in01f80 g747598 ( .a(n_32305), .o(n_32282) );
ao12f80 g771151 ( .a(n_9089), .b(n_9271), .c(n_8309), .o(n_9421) );
in01f80 g758207 ( .a(n_22490), .o(n_22491) );
na02f80 g744675 ( .a(n_35178), .b(n_35123), .o(n_35215) );
in01f80 g768139 ( .a(n_12790), .o(n_12910) );
ao12f80 g768376 ( .a(n_12228), .b(n_12481), .c(n_12294), .o(n_12509) );
in01f80 newInst_3250 ( .a(newNet_3249), .o(newNet_3250) );
no02f80 g737593 ( .a(n_42505), .b(n_42549), .o(n_42524) );
na02f80 g740888 ( .a(n_39290), .b(n_39191), .o(n_39347) );
no02f80 g741972 ( .a(n_38013), .b(n_38007), .o(n_38059) );
no02f80 g762976 ( .a(n_17490), .b(n_16942), .o(n_17566) );
na02f80 g775342 ( .a(n_5909), .b(FE_OCPN1050_n_4459), .o(n_6007) );
in01f80 g745702 ( .a(n_35453), .o(n_35454) );
na02f80 g766937 ( .a(n_13966), .b(n_14006), .o(n_14493) );
ms00f80 delay_sub_ln23_0_unr26_stage9_stallmux_q_reg_0_ ( .ck(newNet_1453), .d(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_) );
na02f80 FE_RC_1105_0 ( .a(n_3361), .b(FE_OCP_RBN2290_n_2438), .o(FE_RN_330_0) );
in01f80 g750519 ( .a(n_30475), .o(n_30552) );
no02f80 g773905 ( .a(n_7094), .b(n_7056), .o(n_7057) );
no02f80 g771631 ( .a(n_8746), .b(n_8701), .o(n_8817) );
in01f80 newInst_183 ( .a(newNet_182), .o(newNet_183) );
na02f80 g769285 ( .a(n_11585), .b(n_11112), .o(n_11579) );
in01f80 g770926 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_10167) );
no02f80 FE_RC_2866_0 ( .a(FE_RN_1234_0), .b(FE_RN_1235_0), .o(FE_RN_1236_0) );
oa22f80 FE_RC_3350_0 ( .a(FE_OCP_RBN3633_n_20568), .b(n_21037), .c(FE_OCP_RBN3632_n_20568), .d(n_21002), .o(n_21203) );
in01f80 FE_RC_3207_0 ( .a(FE_RN_1425_0), .o(FE_RN_1424_0) );
in01f80 g744058 ( .a(n_35784), .o(n_35909) );
na02f80 g770237 ( .a(n_10817), .b(n_10816), .o(n_10818) );
in01f80 g737545 ( .a(n_42510), .o(n_42511) );
no02f80 g752762 ( .a(n_27402), .b(n_27307), .o(n_27512) );
in01f80 g780356 ( .a(n_949), .o(n_1005) );
in01f80 FE_OFC837_n_4298 ( .a(n_4298), .o(FE_OFN837_n_4298) );
in01f80 newInst_1507 ( .a(newNet_1506), .o(newNet_1507) );
na02f80 g769676 ( .a(n_11272), .b(n_11264), .o(n_11314) );
in01f80 g754589 ( .a(n_26890), .o(n_26891) );
na02f80 g769661 ( .a(n_11299), .b(n_11231), .o(n_11315) );
no02f80 g777335 ( .a(n_4759), .b(n_5197), .o(n_5241) );
in01f80 FE_OCP_RBC1927_cordic_combinational_sub_ln23_0_unr12_z_0__ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN1927_cordic_combinational_sub_ln23_0_unr12_z_0__) );
in01f80 newInst_308 ( .a(newNet_307), .o(newNet_308) );
oa12f80 g774618 ( .a(n_6205), .b(n_6485), .c(n_6213), .o(n_6489) );
na02f80 FE_RC_1745_0 ( .a(n_12252), .b(n_12375), .o(FE_RN_490_0) );
in01f80 g749639 ( .a(n_30322), .o(n_30323) );
ao12f80 g757872 ( .a(n_22855), .b(n_22738), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .o(n_22983) );
in01f80 fopt782888 ( .a(n_22874), .o(n_44327) );
in01f80 g743970 ( .a(n_36009), .o(n_36010) );
ao12f80 g762670 ( .a(n_17927), .b(n_17928), .c(n_17926), .o(n_19384) );
oa12f80 g747484 ( .a(n_33721), .b(n_33682), .c(n_33571), .o(n_33815) );
in01f80 g774849 ( .a(n_6319), .o(n_6341) );
in01f80 FE_OCP_RBC3436_n_29163 ( .a(n_29163), .o(FE_OCP_RBN3436_n_29163) );
oa12f80 g739874 ( .a(n_40153), .b(n_40379), .c(n_40274), .o(n_40414) );
na02f80 g751708 ( .a(n_28356), .b(n_28404), .o(n_28417) );
in01f80 g766329 ( .a(n_14436), .o(n_14437) );
ao22s80 FE_RC_118_0 ( .a(n_19052), .b(n_19135), .c(FE_OCP_RBN1691_n_19052), .d(n_19136), .o(n_19315) );
oa12f80 g743821 ( .a(n_35836), .b(n_35835), .c(n_35834), .o(n_35922) );
no02f80 g768052 ( .a(FE_OCPN860_n_12880), .b(n_13074), .o(n_13111) );
in01f80 FE_OCP_RBC2614_n_35005 ( .a(n_35005), .o(FE_OCP_RBN2614_n_35005) );
in01f80 g756469 ( .a(n_23687), .o(n_23688) );
na02f80 g764513 ( .a(n_15918), .b(n_15860), .o(n_16095) );
in01f80 g747841 ( .a(n_33391), .o(n_33353) );
in01f80 newInst_3486 ( .a(newNet_3485), .o(newNet_3486) );
in01f80 newInst_2640 ( .a(newNet_1553), .o(newNet_2640) );
oa12f80 g736346 ( .a(n_43525), .b(n_43814), .c(n_43360), .o(n_43827) );
in01f80 g779548 ( .a(n_1426), .o(n_1427) );
oa12f80 g745888 ( .a(n_34063), .b(n_34048), .c(n_34030), .o(n_34094) );
in01f80 FE_OFC841_n_15791 ( .a(n_15791), .o(FE_OFN841_n_15791) );
na02f80 g741246 ( .a(FE_OCP_RBN2636_n_38806), .b(n_38511), .o(n_39012) );
in01f80 g766517 ( .a(n_16143), .o(n_14355) );
in01f80 newInst_1811 ( .a(newNet_1810), .o(newNet_1811) );
in01f80 newInst_2203 ( .a(newNet_2202), .o(newNet_2203) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_0_ ( .ck(newNet_1152), .d(n_9324), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_0_) );
no02f80 g778320 ( .a(n_2524), .b(n_2523), .o(n_2525) );
in01f80 newInst_621 ( .a(newNet_620), .o(newNet_621) );
no03m80 g743291 ( .a(n_37857), .b(n_37856), .c(n_37827), .o(n_37878) );
oa12f80 g738454 ( .a(n_41679), .b(FE_OCPN952_n_41540), .c(n_41698), .o(n_41853) );
in01f80 newInst_2932 ( .a(newNet_2931), .o(newNet_2932) );
in01f80 g738438 ( .a(n_41904), .o(n_41905) );
in01f80 newInst_564 ( .a(newNet_563), .o(newNet_564) );
oa12f80 g758182 ( .a(n_21899), .b(n_21968), .c(n_21845), .o(n_22020) );
in01f80 newInst_3635 ( .a(newNet_3634), .o(newNet_3635) );
in01f80 newInst_92 ( .a(newNet_50), .o(newNet_92) );
na02f80 g775364 ( .a(n_5668), .b(n_5634), .o(n_5810) );
oa12f80 g748504 ( .a(FE_OCP_RBN3712_n_31466), .b(FE_OCP_RBN2829_n_30731), .c(FE_OCP_RBN2807_n_30643), .o(n_31652) );
in01f80 FE_OFC800_n_46285 ( .a(FE_OFN797_n_46285), .o(FE_OFN800_n_46285) );
oa12f80 g772334 ( .a(n_8718), .b(n_8717), .c(n_8716), .o(n_9647) );
na02f80 FE_RC_2449_0 ( .a(FE_RN_978_0), .b(n_13164), .o(FE_RN_979_0) );
in01f80 newInst_799 ( .a(newNet_798), .o(newNet_799) );
in01f80 g755925 ( .a(n_24293), .o(n_24310) );
in01f80 newInst_3034 ( .a(newNet_3033), .o(newNet_3034) );
no02f80 g762199 ( .a(n_18626), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_18627) );
oa12f80 g752522 ( .a(n_27426), .b(n_27645), .c(n_27343), .o(n_27684) );
na02f80 g750447 ( .a(n_29547), .b(n_25859), .o(n_29604) );
in01f80 g744722 ( .a(n_35184), .o(n_35157) );
in01f80 g775153 ( .a(n_6105), .o(n_6071) );
oa22f80 g784557 ( .a(FE_OFN801_n_46285), .b(n_11297), .c(FE_OCP_RBN3044_n_46337), .d(n_11265), .o(n_46378) );
oa12f80 g760296 ( .a(n_20928), .b(n_20834), .c(n_20927), .o(n_21625) );
no02f80 g746433 ( .a(n_33424), .b(n_33423), .o(n_33425) );
in01f80 g757498 ( .a(n_22867), .o(n_22868) );
na03f80 FE_RC_2230_0 ( .a(FE_RN_808_0), .b(FE_RN_811_0), .c(n_37033), .o(n_37193) );
na02f80 g744984 ( .a(n_34923), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34953) );
in01f80 FE_OCPC910_n_43022 ( .a(FE_OCP_RBN3700_n_43015), .o(FE_OCPN910_n_43022) );
in01f80 FE_OCP_RBC3588_n_9408 ( .a(n_9408), .o(FE_OCP_RBN3588_n_9408) );
no02f80 g750417 ( .a(n_29566), .b(n_29561), .o(n_29643) );
na02f80 g736846 ( .a(n_43026), .b(n_43025), .o(n_43039) );
oa12f80 g738958 ( .a(n_41061), .b(n_41186), .c(n_40935), .o(n_41223) );
in01f80 g770339 ( .a(n_10660), .o(n_10661) );
oa22f80 g770433 ( .a(n_10633), .b(n_9813), .c(n_10551), .d(n_9814), .o(n_10652) );
in01f80 FE_RC_4192_0 ( .a(FE_RN_1836_0), .o(FE_RN_1834_0) );
no02f80 FE_RC_3845_0 ( .a(n_23407), .b(FE_RN_1676_0), .o(FE_RN_1677_0) );
in01f80 FE_RC_2694_0 ( .a(FE_RN_1129_0), .o(n_8855) );
in01f80 g750027 ( .a(n_30367), .o(n_30368) );
no02f80 g736592 ( .a(n_43636), .b(n_43391), .o(n_43649) );
no02f80 g772819 ( .a(n_8019), .b(n_8055), .o(n_8056) );
na02f80 g739460 ( .a(n_40668), .b(n_40667), .o(n_40735) );
ao12f80 g768351 ( .a(n_12444), .b(n_12443), .c(n_12442), .o(n_12838) );
na02f80 g755098 ( .a(n_25180), .b(n_25179), .o(n_25207) );
in01f80 newInst_989 ( .a(newNet_988), .o(newNet_989) );
in01f80 g753505 ( .a(n_26844), .o(n_26845) );
in01f80 g776498 ( .a(n_4441), .o(n_4442) );
na02f80 g770949 ( .a(n_10049), .b(n_10004), .o(n_10005) );
na02f80 g775320 ( .a(n_5830), .b(n_5835), .o(n_5952) );
in01f80 g770810 ( .a(n_10141), .o(n_10142) );
oa22f80 FE_RC_950_0 ( .a(n_20231), .b(n_22914), .c(n_22793), .d(FE_OCP_RBN1223_n_22914), .o(n_22973) );
no02f80 g746610 ( .a(n_34390), .b(n_34389), .o(n_34475) );
no02f80 g776121 ( .a(n_4848), .b(n_4620), .o(n_4837) );
oa12f80 g772253 ( .a(n_8045), .b(n_8760), .c(n_8038), .o(n_8821) );
oa12f80 g770715 ( .a(n_10303), .b(n_10334), .c(n_10302), .o(n_10389) );
na02f80 FE_RC_2850_0 ( .a(n_19739), .b(n_19877), .o(FE_RN_1227_0) );
in01f80 g762061 ( .a(n_18963), .o(n_19406) );
in01f80 newInst_1824 ( .a(newNet_1823), .o(newNet_1824) );
in01f80 FE_OCP_RBC2458_n_13765 ( .a(FE_OCP_RBN2456_n_13765), .o(FE_OCP_RBN2458_n_13765) );
oa22f80 g754192 ( .a(n_25900), .b(n_25616), .c(n_25901), .d(n_25615), .o(n_25997) );
in01f80 newInst_2973 ( .a(newNet_2972), .o(newNet_2973) );
in01f80 g780874 ( .a(n_414), .o(n_415) );
in01f80 g780156 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_3_), .o(n_1178) );
in01f80 g763305 ( .a(n_17085), .o(n_17086) );
na02f80 FE_RC_3486_0 ( .a(n_37375), .b(FE_RN_1499_0), .o(FE_RN_1501_0) );
no02f80 FE_RC_4020_0 ( .a(FE_RN_1745_0), .b(n_20549), .o(FE_RN_1746_0) );
no02f80 g781169 ( .a(n_182), .b(n_58), .o(n_180) );
in01f80 g762855 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_30_), .o(n_17749) );
in01f80 FE_RC_4243_0 ( .a(n_26473), .o(FE_RN_1865_0) );
ao12f80 g766974 ( .a(n_13614), .b(n_13613), .c(n_13612), .o(n_15458) );
no02f80 g768405 ( .a(n_12449), .b(n_11961), .o(n_12459) );
na02f80 g738207 ( .a(n_41977), .b(n_41749), .o(n_41985) );
ao12f80 g751084 ( .a(n_29803), .b(n_29802), .c(n_29801), .o(n_29852) );
in01f80 g756511 ( .a(n_23759), .o(n_23760) );
na02f80 g769824 ( .a(n_11084), .b(n_11122), .o(n_11141) );
in01f80 g771372 ( .a(n_9425), .o(n_9426) );
oa12f80 g757630 ( .a(n_22271), .b(n_45497), .c(n_22130), .o(n_22636) );
in01f80 FE_RC_3541_0 ( .a(FE_RN_1534_0), .o(n_19272) );
in01f80 FE_OCP_RBC1717_n_20734 ( .a(FE_OCP_RBN1716_n_20734), .o(FE_OCP_RBN1717_n_20734) );
in01f80 newInst_196 ( .a(newNet_95), .o(newNet_196) );
no02f80 g745198 ( .a(n_34597), .b(n_34596), .o(n_34598) );
no02f80 g744276 ( .a(n_44180), .b(n_34989), .o(n_36130) );
in01f80 newInst_3710 ( .a(newNet_3709), .o(newNet_3710) );
no02f80 g778906 ( .a(n_2160), .b(n_1956), .o(n_2179) );
no02f80 g744233 ( .a(n_36859), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n_36861) );
no02f80 g746756 ( .a(n_34132), .b(n_33705), .o(n_34172) );
na02f80 g753171 ( .a(n_27410), .b(n_27376), .o(n_27519) );
in01f80 g736822 ( .a(n_43261), .o(n_43262) );
in01f80 g753400 ( .a(n_27081), .o(n_27082) );
oa12f80 g761745 ( .a(n_18480), .b(n_18789), .c(n_18482), .o(n_18822) );
na02f80 g765041 ( .a(FE_OCP_RBN3648_n_15281), .b(n_14210), .o(n_15502) );
in01f80 g737076 ( .a(n_43325), .o(n_43291) );
na02f80 g751949 ( .a(n_28754), .b(n_28753), .o(n_28755) );
in01f80 g765899 ( .a(n_14906), .o(n_14853) );
in01f80 g748103 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_9_), .o(n_32989) );
in01f80 g776986 ( .a(n_3979), .o(n_3980) );
oa12f80 g780346 ( .a(n_45815), .b(n_832), .c(n_831), .o(n_833) );
na02f80 g739030 ( .a(n_41178), .b(n_41177), .o(n_41179) );
no02f80 g747281 ( .a(n_45753), .b(n_33497), .o(n_33748) );
no02f80 g760932 ( .a(n_19255), .b(n_18507), .o(n_19283) );
in01f80 g779325 ( .a(n_1678), .o(n_1679) );
na02f80 g743986 ( .a(n_35646), .b(n_35645), .o(n_35647) );
ao12f80 g780425 ( .a(n_878), .b(n_1203), .c(n_1099), .o(n_902) );
no02f80 g741184 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39324), .o(n_39358) );
na02f80 g741410 ( .a(n_38801), .b(n_38797), .o(n_38798) );
in01f80 fopt782675 ( .a(n_44071), .o(n_44068) );
no02f80 g745319 ( .a(n_35937), .b(n_35763), .o(n_35803) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_21_ ( .ck(newNet_169), .d(n_46350), .o(delay_xor_ln22_unr9_stage4_stallmux_q_21_) );
no02f80 g753920 ( .a(n_26286), .b(n_26262), .o(n_26429) );
na02f80 FE_RC_3755_0 ( .a(FE_OCP_RBN3378_n_40716), .b(FE_RN_1649_0), .o(FE_RN_1650_0) );
na02f80 FE_RC_3047_0 ( .a(n_26727), .b(n_26729), .o(FE_RN_1334_0) );
na02f80 g752539 ( .a(n_27599), .b(n_27550), .o(n_27672) );
in01f80 g747941 ( .a(n_33226), .o(n_33238) );
in01f80 FE_OCPC1043_n_20307 ( .a(n_20307), .o(FE_OCPN1043_n_20307) );
no02f80 g756281 ( .a(n_23976), .b(n_23667), .o(n_24072) );
in01f80 FE_OCP_RBC2537_n_3645 ( .a(n_3645), .o(FE_OCP_RBN2537_n_3645) );
no02f80 g755873 ( .a(n_25193), .b(n_25220), .o(n_25839) );
na03f80 g737727 ( .a(n_42360), .b(n_42328), .c(n_42359), .o(n_42361) );
ao12f80 g767250 ( .a(n_13681), .b(n_13680), .c(n_13679), .o(n_14168) );
no02f80 g776930 ( .a(n_3764), .b(FE_OCP_RBN2623_n_3631), .o(n_3863) );
no02f80 g784774 ( .a(n_9724), .b(n_8750), .o(n_47260) );
na02f80 g771756 ( .a(n_9110), .b(n_44575), .o(n_9330) );
in01f80 FE_OCP_RBC2670_n_20249 ( .a(FE_OCP_RBN1333_n_20249), .o(FE_OCP_RBN2670_n_20249) );
na02f80 g770566 ( .a(n_10278), .b(n_9041), .o(n_10699) );
in01f80 g758215 ( .a(n_22877), .o(n_22878) );
na02f80 g781127 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_6_), .o(n_236) );
na02f80 g777267 ( .a(n_3578), .b(n_2913), .o(n_3668) );
in01f80 g774806 ( .a(n_6394), .o(n_6279) );
no02f80 g758062 ( .a(n_22918), .b(n_22917), .o(n_23382) );
in01f80 g766018 ( .a(n_14808), .o(n_14843) );
in01f80 newInst_1364 ( .a(newNet_1363), .o(newNet_1364) );
ao22s80 FE_RC_816_0 ( .a(n_8731), .b(n_8926), .c(FE_OCP_RBN2475_n_8664), .d(n_8960), .o(n_9125) );
na02f80 g749631 ( .a(n_31433), .b(n_31460), .o(n_31461) );
no02f80 g736801 ( .a(n_43266), .b(n_43265), .o(n_43267) );
in01f80 g748267 ( .a(n_31863), .o(n_31898) );
na02f80 g779127 ( .a(n_2015), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_12_), .o(n_2032) );
in01f80 g748453 ( .a(n_31718), .o(n_31765) );
in01f80 newInst_1841 ( .a(newNet_978), .o(newNet_1841) );
na02f80 g775148 ( .a(n_5989), .b(n_5988), .o(n_6012) );
no02f80 g750431 ( .a(n_30519), .b(n_30034), .o(n_30634) );
ao22s80 g780856 ( .a(n_457), .b(n_193), .c(n_420), .d(FE_OCPN1386_n_470), .o(n_539) );
in01f80 g751349 ( .a(n_29935), .o(n_29490) );
ao12f80 g743067 ( .a(n_37046), .b(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n_37500) );
na02f80 g755119 ( .a(n_25315), .b(n_25316), .o(n_25350) );
in01f80 newInst_3509 ( .a(newNet_3508), .o(newNet_3509) );
in01f80 newInst_2910 ( .a(newNet_2909), .o(newNet_2910) );
in01f80 fopt782750 ( .a(n_44166), .o(n_44165) );
in01f80 g770014 ( .a(n_10944), .o(n_10962) );
in01f80 FE_OCPC1795_n_30546 ( .a(n_30546), .o(FE_OCPN1795_n_30546) );
in01f80 g758821 ( .a(n_21581), .o(n_21582) );
ao12f80 g766988 ( .a(n_13771), .b(n_13770), .c(n_13769), .o(n_14259) );
in01f80 newInst_1567 ( .a(newNet_825), .o(newNet_1567) );
in01f80 g749228 ( .a(n_32158), .o(n_32176) );
na02f80 g766730 ( .a(n_13829), .b(FE_OCP_RBN3484_n_13667), .o(n_13851) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_23_ ( .ck(newNet_1312), .d(n_1261), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_) );
no02f80 g776437 ( .a(n_4104), .b(n_4006), .o(n_4185) );
no02f80 g743239 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_1_), .b(delay_add_ln22_unr23_stage9_stallmux_q_1_), .o(n_36847) );
in01f80 g746559 ( .a(n_33306), .o(n_33272) );
na02f80 g775240 ( .a(n_5952), .b(n_5940), .o(n_6008) );
na02f80 g757100 ( .a(n_23547), .b(n_23085), .o(n_23643) );
na02f80 g739319 ( .a(n_45153), .b(n_40891), .o(n_40889) );
no02f80 g747996 ( .a(n_31997), .b(n_31934), .o(n_32081) );
na02f80 g760047 ( .a(n_20413), .b(n_20342), .o(n_20439) );
no02f80 g779624 ( .a(n_1800), .b(delay_xor_ln21_unr3_stage2_stallmux_q_25_), .o(n_2082) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_12_ ( .ck(newNet_2494), .d(n_32251), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_) );
no02f80 g754432 ( .a(n_25726), .b(n_25457), .o(n_25727) );
oa12f80 g770399 ( .a(n_10153), .b(n_10243), .c(n_10197), .o(n_10405) );
in01f80 FE_OCP_RBC2372_n_8221 ( .a(FE_OCP_RBN2371_n_8221), .o(FE_OCP_RBN2372_n_8221) );
ao12f80 g755600 ( .a(n_25062), .b(n_25093), .c(n_24953), .o(n_25172) );
na02f80 g756371 ( .a(n_23795), .b(n_23794), .o(n_23796) );
na02f80 g766963 ( .a(n_13529), .b(n_13534), .o(n_13599) );
oa12f80 g774982 ( .a(n_5823), .b(n_6082), .c(n_5681), .o(n_6138) );
in01f80 g756614 ( .a(n_23738), .o(n_23675) );
na02f80 g768579 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_24_), .b(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_12892) );
na02f80 g757039 ( .a(n_23700), .b(n_23746), .o(n_23834) );
no02f80 g763259 ( .a(n_16953), .b(n_17045), .o(n_17046) );
no02f80 g777615 ( .a(n_3456), .b(n_3448), .o(n_3449) );
in01f80 g744092 ( .a(n_35693), .o(n_35694) );
no02f80 g767693 ( .a(n_12807), .b(n_12869), .o(n_12864) );
na02f80 g773767 ( .a(n_7150), .b(n_7077), .o(n_7186) );
na02f80 FE_RC_2467_0 ( .a(n_14042), .b(FE_RN_991_0), .o(FE_RN_992_0) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_27_ ( .ck(newNet_2082), .d(n_6643), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_) );
no02f80 g777185 ( .a(n_3998), .b(n_4108), .o(n_4269) );
na02f80 FE_RC_2612_0 ( .a(n_1426), .b(FE_RN_1086_0), .o(n_1491) );
no02f80 g774324 ( .a(FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_4_), .o(n_6715) );
no02f80 g771466 ( .a(n_9442), .b(n_7979), .o(n_9609) );
in01f80 g778191 ( .a(n_3494), .o(n_2784) );
oa12f80 g759032 ( .a(n_21408), .b(n_21977), .c(n_21377), .o(n_22058) );
no02f80 g741040 ( .a(n_38833), .b(n_38862), .o(n_38863) );
in01f80 g764981 ( .a(FE_OCP_RBN2812_n_15433), .o(n_15479) );
na02f80 g738242 ( .a(n_41899), .b(n_41898), .o(n_41900) );
in01f80 g757214 ( .a(n_23546), .o(n_23547) );
na02f80 g764504 ( .a(n_16216), .b(n_16215), .o(n_16267) );
no02f80 g738392 ( .a(n_41453), .b(n_41428), .o(n_41454) );
no02f80 g778920 ( .a(n_2189), .b(n_1957), .o(n_2190) );
in01f80 newInst_2805 ( .a(newNet_2804), .o(newNet_2805) );
in01f80 newInst_84 ( .a(newNet_83), .o(newNet_84) );
in01f80 FE_OCP_RBC3562_n_29857 ( .a(n_29857), .o(FE_OCP_RBN3562_n_29857) );
in01f80 g776008 ( .a(n_5244), .o(n_5210) );
na02f80 g740526 ( .a(n_39676), .b(n_39675), .o(n_39689) );
in01f80 g742943 ( .a(n_37187), .o(n_37113) );
na02f80 g754820 ( .a(n_25511), .b(n_25451), .o(n_25782) );
in01f80 newInst_3258 ( .a(newNet_3257), .o(newNet_3258) );
no02f80 g753196 ( .a(n_27207), .b(n_25962), .o(n_27391) );
oa22f80 FE_RC_409_0 ( .a(n_13207), .b(n_14280), .c(n_13206), .d(n_14279), .o(n_14444) );
in01f80 g755511 ( .a(n_24799), .o(n_24819) );
no02f80 g770051 ( .a(n_10765), .b(n_10470), .o(n_10793) );
in01f80 FE_OCP_RBC2970_n_42896 ( .a(n_42896), .o(FE_OCP_RBN2970_n_42896) );
in01f80 FE_OCP_RBC2589_n_9492 ( .a(n_9492), .o(FE_OCP_RBN2589_n_9492) );
oa12f80 g780098 ( .a(n_1097), .b(n_1119), .c(n_1096), .o(n_1136) );
na02f80 g771566 ( .a(n_9395), .b(n_9394), .o(n_9519) );
no02f80 g741596 ( .a(n_38648), .b(n_38649), .o(n_38660) );
in01f80 g739571 ( .a(n_40627), .o(n_40628) );
no02f80 g747733 ( .a(n_33258), .b(n_33242), .o(n_33298) );
in01f80 g749499 ( .a(n_30465), .o(n_30499) );
na02f80 g740972 ( .a(n_39109), .b(n_39271), .o(n_39281) );
na02f80 g743203 ( .a(n_37032), .b(n_36917), .o(n_36985) );
in01f80 g760408 ( .a(n_20127), .o(n_20128) );
na02f80 g750467 ( .a(n_30475), .b(n_29990), .o(n_30518) );
in01f80 g737776 ( .a(n_42348), .o(n_42349) );
in01f80 g757020 ( .a(n_23747), .o(n_23721) );
in01f80 g753961 ( .a(n_26253), .o(n_26254) );
no02f80 g772463 ( .a(n_8463), .b(n_8455), .o(n_8540) );
na02f80 g753556 ( .a(n_27406), .b(n_26897), .o(n_27451) );
in01f80 g752839 ( .a(n_28314), .o(n_28315) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_10_ ( .ck(newNet_2596), .d(n_27059), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_10_) );
no02f80 g739240 ( .a(n_40781), .b(n_40733), .o(n_41016) );
in01f80 g746869 ( .a(n_33178), .o(n_33179) );
in01f80 g754287 ( .a(n_25915), .o(n_25914) );
na02f80 g772716 ( .a(n_8202), .b(n_8217), .o(n_8318) );
in01f80 g773236 ( .a(n_7596), .o(n_7597) );
oa12f80 g749893 ( .a(FE_OCP_RBN3013_n_31117), .b(n_31211), .c(n_31172), .o(n_31212) );
ao12f80 g738277 ( .a(n_41786), .b(n_41888), .c(n_41825), .o(n_41870) );
na02f80 g767388 ( .a(n_13406), .b(n_13405), .o(n_13407) );
in01f80 newInst_1764 ( .a(newNet_1763), .o(newNet_1764) );
in01f80 g757859 ( .a(n_22479), .o(n_22443) );
na02f80 g745399 ( .a(n_34653), .b(n_34590), .o(n_34675) );
na02f80 g769862 ( .a(n_11180), .b(n_10240), .o(n_11211) );
oa12f80 g752457 ( .a(n_27469), .b(n_27648), .c(n_27371), .o(n_27695) );
oa12f80 g768991 ( .a(n_11769), .b(n_11659), .c(FE_OCP_RBN3266_n_45224), .o(n_11983) );
in01f80 g771489 ( .a(n_9400), .o(n_9401) );
na02f80 g753442 ( .a(n_26880), .b(n_26963), .o(n_26964) );
oa22f80 FE_RC_1193_0 ( .a(n_13172), .b(n_13711), .c(FE_OCP_RBN3480_n_13664), .d(n_13180), .o(n_13751) );
in01f80 newInst_265 ( .a(newNet_264), .o(newNet_265) );
no02f80 FE_RC_3520_0 ( .a(FE_RN_1520_0), .b(n_23110), .o(n_23176) );
in01f80 newInst_1299 ( .a(newNet_1298), .o(newNet_1299) );
no02f80 g761315 ( .a(n_19789), .b(n_19830), .o(n_19852) );
no02f80 g761784 ( .a(n_18821), .b(n_18743), .o(n_18850) );
no03m80 FE_RC_1088_0 ( .a(n_37090), .b(n_36981), .c(n_37173), .o(n_37209) );
in01f80 g776938 ( .a(n_4019), .o(n_4020) );
in01f80 FE_OCPC3788_n_15708 ( .a(n_15708), .o(FE_OCPN3788_n_15708) );
in01f80 g768652 ( .a(n_12287), .o(n_12288) );
na02f80 FE_RC_1787_0 ( .a(FE_RN_524_0), .b(n_28399), .o(FE_RN_525_0) );
in01f80 g746049 ( .a(n_34004), .o(n_34005) );
na02f80 g775239 ( .a(n_5837), .b(n_5857), .o(n_5917) );
na02f80 g768863 ( .a(n_11777), .b(n_11609), .o(n_11853) );
na02f80 g784788 ( .a(FE_OCP_RBN3085_n_31819), .b(FE_OCP_RBN2912_n_30908), .o(n_47274) );
na02f80 g761394 ( .a(n_18831), .b(n_18875), .o(n_18987) );
na02f80 g755330 ( .a(n_24918), .b(n_24876), .o(n_24971) );
na02f80 g764481 ( .a(n_16113), .b(n_16037), .o(n_16160) );
in01f80 FE_OCPC1529_n_26090 ( .a(n_26090), .o(FE_OCPN1529_n_26090) );
na02f80 g743312 ( .a(n_37857), .b(n_37856), .o(n_37858) );
oa12f80 g773990 ( .a(n_6898), .b(n_6897), .c(n_6896), .o(n_7795) );
ao12f80 g756059 ( .a(n_25139), .b(n_25133), .c(n_25129), .o(n_25195) );
in01f80 g738894 ( .a(n_41254), .o(n_41255) );
no02f80 g742219 ( .a(n_44887), .b(n_38325), .o(n_38326) );
ao12f80 g745567 ( .a(n_34249), .b(n_34248), .c(n_34250), .o(n_35427) );
in01f80 g737141 ( .a(n_43046), .o(n_43082) );
in01f80 newInst_824 ( .a(newNet_823), .o(newNet_824) );
in01f80 FE_OCP_DRV_C1584_n_30917 ( .a(FE_OCP_DRV_N1583_n_30917), .o(FE_OCP_DRV_N1584_n_30917) );
na02f80 g774788 ( .a(n_45474), .b(FE_OCP_RBN2978_n_5555), .o(n_6327) );
in01f80 g778523 ( .a(n_2566), .o(n_2567) );
in01f80 g776004 ( .a(n_5321), .o(n_5322) );
na02f80 g744645 ( .a(n_35342), .b(FE_OCP_RBN3664_n_35326), .o(n_35358) );
no02f80 g756402 ( .a(n_24162), .b(n_23740), .o(n_23858) );
in01f80 g743192 ( .a(n_37030), .o(n_36930) );
ao22s80 g750842 ( .a(FE_OCP_RBN1325_n_29056), .b(FE_OFN811_n_29140), .c(FE_OCP_RBN1324_n_29056), .d(n_27961), .o(n_29228) );
no02f80 g779383 ( .a(n_1551), .b(n_1545), .o(n_1546) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_8_ ( .ck(newNet_1893), .d(n_36891), .o(n_46254) );
no03m80 FE_RC_171_0 ( .a(n_17192), .b(n_17084), .c(n_17133), .o(n_17401) );
no02f80 g771417 ( .a(n_9340), .b(n_9274), .o(n_9513) );
in01f80 g739612 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_1_), .o(n_40614) );
in01f80 FE_OCP_RBC3075_FE_OFN807_n_46195 ( .a(FE_OFN807_n_46195), .o(FE_OCP_RBN3075_FE_OFN807_n_46195) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_9_ ( .ck(newNet_3183), .d(n_35990), .o(delay_add_ln22_unr23_stage9_stallmux_q_9_) );
oa12f80 g746425 ( .a(n_34617), .b(n_34473), .c(n_34646), .o(n_35020) );
in01f80 g755785 ( .a(n_24369), .o(n_24370) );
in01f80 g778915 ( .a(n_2271), .o(n_2272) );
oa22f80 g747971 ( .a(n_32079), .b(n_32163), .c(n_32060), .d(FE_OCP_RBN3103_n_32163), .o(n_32234) );
in01f80 newInst_548 ( .a(newNet_547), .o(newNet_548) );
oa22f80 g745114 ( .a(n_36252), .b(n_36114), .c(n_36253), .d(n_36113), .o(n_36330) );
na02f80 g779819 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_28_), .o(n_2115) );
in01f80 newInst_426 ( .a(newNet_405), .o(newNet_426) );
oa22f80 g746562 ( .a(n_34810), .b(FE_RN_876_0), .c(n_34666), .d(n_34733), .o(n_35337) );
oa22f80 g779874 ( .a(n_44659), .b(n_886), .c(n_44661), .d(n_822), .o(n_1291) );
oa12f80 g777978 ( .a(n_2866), .b(n_3056), .c(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(n_3122) );
na02f80 g759515 ( .a(n_20853), .b(n_20852), .o(n_20883) );
in01f80 fopt783812 ( .a(FE_OCP_RBN1195_n_22542), .o(n_45497) );
oa12f80 g743618 ( .a(n_37435), .b(n_37437), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37517) );
in01f80 g749083 ( .a(n_30863), .o(n_30864) );
in01f80 newInst_2015 ( .a(newNet_2014), .o(newNet_2015) );
oa22f80 g784562 ( .a(FE_OFN800_n_46285), .b(n_46988), .c(FE_OCP_RBN3709_n_46337), .d(n_10980), .o(n_46383) );
in01f80 g774471 ( .a(n_6630), .o(n_6688) );
in01f80 g746204 ( .a(n_33807), .o(n_33773) );
no02f80 FE_RC_2088_0 ( .a(FE_OCP_RBN1146_n_13098), .b(n_14372), .o(FE_RN_716_0) );
in01f80 g776751 ( .a(n_3981), .o(n_4009) );
na02f80 FE_RC_2728_0 ( .a(FE_RN_1153_0), .b(FE_RN_1154_0), .o(FE_RN_1155_0) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_16_ ( .ck(newNet_2872), .d(n_11297), .o(delay_add_ln22_unr8_stage4_stallmux_q_16_) );
in01f80 g754138 ( .a(n_26069), .o(n_26029) );
oa12f80 g770524 ( .a(n_10492), .b(n_10527), .c(n_10491), .o(n_10549) );
na02f80 g755742 ( .a(n_24492), .b(n_24491), .o(n_24493) );
no02f80 g746727 ( .a(n_34212), .b(n_34211), .o(n_34252) );
ao12f80 g741460 ( .a(n_38782), .b(n_38781), .c(n_38780), .o(n_39747) );
in01f80 g779741 ( .a(n_1629), .o(n_1596) );
in01f80 newInst_3385 ( .a(newNet_3307), .o(newNet_3385) );
in01f80 g737744 ( .a(n_42449), .o(n_42433) );
in01f80 g753312 ( .a(n_27326), .o(n_27371) );
na02f80 g746963 ( .a(n_32876), .b(n_32875), .o(n_32877) );
oa12f80 g778502 ( .a(n_2817), .b(n_2834), .c(n_2768), .o(n_2880) );
na02f80 g758766 ( .a(n_22210), .b(n_21566), .o(n_22247) );
in01f80 g763183 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_), .o(n_18291) );
ao12f80 g780745 ( .a(n_589), .b(n_590), .c(n_411), .o(n_594) );
no02f80 g779387 ( .a(n_1547), .b(n_1542), .o(n_1577) );
no02f80 g763730 ( .a(n_17310), .b(n_17309), .o(n_17614) );
in01f80 FE_OCP_DRV_C1538_n_13646 ( .a(FE_OCP_DRV_N1537_n_13646), .o(FE_OCP_DRV_N1538_n_13646) );
in01f80 FE_RC_2412_0 ( .a(FE_RN_952_0), .o(n_45488) );
no02f80 g780898 ( .a(n_403), .b(n_417), .o(n_442) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_17_ ( .ck(newNet_1531), .d(n_32229), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_17_) );
no02f80 g770027 ( .a(n_10884), .b(n_10883), .o(n_10917) );
na02f80 FE_RC_2126_0 ( .a(n_24429), .b(FE_OCP_RBN2596_n_25181), .o(FE_RN_741_0) );
no02f80 g743844 ( .a(n_35673), .b(n_35575), .o(n_35714) );
no02f80 g753819 ( .a(n_26373), .b(n_23353), .o(n_26407) );
in01f80 g775354 ( .a(FE_OCP_RBN2978_n_5555), .o(n_5636) );
no03m80 FE_RC_1116_0 ( .a(n_40738), .b(n_40749), .c(n_40750), .o(n_40751) );
in01f80 newInst_286 ( .a(newNet_285), .o(newNet_286) );
ms00f80 delay_sub_ln23_0_unr7_stage4_stallmux_q_reg ( .ck(newNet_1157), .d(n_167), .o(cordic_combinational_sub_ln23_0_unr12_z_0_) );
oa12f80 g752310 ( .a(n_27887), .b(n_27888), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(n_29140) );
in01f80 g742201 ( .a(n_37887), .o(n_37888) );
oa22f80 FE_RC_2981_0 ( .a(n_25775), .b(n_26502), .c(n_25776), .d(n_26503), .o(n_26622) );
no02f80 g776974 ( .a(n_3760), .b(n_3846), .o(n_3773) );
in01f80 fopt782790 ( .a(n_44180), .o(n_44174) );
in01f80 g762832 ( .a(n_17940), .o(n_17941) );
in01f80 FE_OCP_RBC2789_n_4294 ( .a(n_4294), .o(FE_OCP_RBN2789_n_4294) );
in01f80 newInst_2159 ( .a(newNet_2158), .o(newNet_2159) );
in01f80 g762443 ( .a(n_18107), .o(n_18108) );
na02f80 g747384 ( .a(n_33578), .b(n_33702), .o(n_33842) );
in01f80 g747859 ( .a(n_33227), .o(n_33670) );
in01f80 newInst_801 ( .a(newNet_507), .o(newNet_801) );
na02f80 g751860 ( .a(n_28191), .b(n_27971), .o(n_28230) );
in01f80 g758024 ( .a(n_22106), .o(n_22132) );
in01f80 g781157 ( .a(n_516), .o(n_200) );
na02f80 g761663 ( .a(n_18756), .b(n_18276), .o(n_18757) );
na02f80 g772763 ( .a(n_47242), .b(n_8109), .o(n_8227) );
in01f80 FE_OFC792_n_25938 ( .a(n_25938), .o(FE_OFN792_n_25938) );
na02f80 g748761 ( .a(n_31139), .b(n_31138), .o(n_31140) );
in01f80 g749694 ( .a(n_30079), .o(n_30152) );
in01f80 g757098 ( .a(n_23144), .o(n_23145) );
in01f80 g763542 ( .a(n_16793), .o(n_16811) );
na02f80 FE_RC_3012_0 ( .a(n_14274), .b(FE_OCP_RBN2709_n_15135), .o(FE_RN_1320_0) );
no02f80 g766506 ( .a(n_14092), .b(n_12877), .o(n_14154) );
na02f80 g777195 ( .a(n_5189), .b(n_5387), .o(n_5415) );
no02f80 g752996 ( .a(n_27226), .b(n_27110), .o(n_27307) );
na02f80 g762134 ( .a(n_18164), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_15_), .o(n_18222) );
oa22f80 g780864 ( .a(n_286), .b(n_145), .c(n_285), .d(n_144), .o(n_504) );
in01f80 newInst_1431 ( .a(newNet_1430), .o(newNet_1431) );
ao12f80 g778934 ( .a(n_2135), .b(n_2143), .c(n_2134), .o(n_2562) );
oa12f80 g780693 ( .a(n_511), .b(n_647), .c(n_645), .o(n_648) );
in01f80 g748161 ( .a(n_32057), .o(n_32058) );
in01f80 g740229 ( .a(n_39773), .o(n_39796) );
na02f80 g745337 ( .a(n_35929), .b(n_35841), .o(n_35930) );
na02f80 g777359 ( .a(n_4219), .b(n_4686), .o(n_4862) );
oa12f80 g755254 ( .a(n_24851), .b(n_24974), .c(n_24892), .o(n_25049) );
no02f80 g766585 ( .a(n_13953), .b(n_13926), .o(n_14072) );
in01f80 newInst_3701 ( .a(newNet_3700), .o(newNet_3701) );
in01f80 g773968 ( .a(n_6960), .o(n_6961) );
no02f80 g738869 ( .a(n_41294), .b(n_41293), .o(n_41295) );
in01f80 newInst_450 ( .a(newNet_2), .o(newNet_450) );
no02f80 g741124 ( .a(n_38957), .b(n_38877), .o(n_38991) );
na02f80 g776555 ( .a(n_4307), .b(n_3297), .o(n_4327) );
in01f80 g762839 ( .a(n_17846), .o(n_17799) );
in01f80 g743301 ( .a(n_36767), .o(n_36780) );
in01f80 g739158 ( .a(n_40913), .o(n_41041) );
na02f80 g773893 ( .a(n_7031), .b(n_6623), .o(n_7083) );
no02f80 g758522 ( .a(n_22145), .b(n_22063), .o(n_22183) );
in01f80 g774447 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_1_), .o(n_6507) );
in01f80 newInst_1280 ( .a(newNet_334), .o(newNet_1280) );
in01f80 drc28 ( .a(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46204) );
no02f80 g773919 ( .a(n_6883), .b(n_6758), .o(n_6941) );
no02f80 g770992 ( .a(n_9742), .b(FE_OCPN903_n_44581), .o(n_9803) );
in01f80 FE_OCP_RBC3694_n_26409 ( .a(n_26409), .o(FE_OCP_RBN3694_n_26409) );
in01f80 g751468 ( .a(n_28914), .o(n_28915) );
na02f80 g769791 ( .a(n_11137), .b(n_11138), .o(n_11254) );
in01f80 g756154 ( .a(FE_OCP_RBN2307_n_24288), .o(n_25386) );
in01f80 g739602 ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_3_), .o(n_40602) );
in01f80 g759797 ( .a(n_21857), .o(n_21858) );
in01f80 g763977 ( .a(FE_OFN779_n_17093), .o(n_17783) );
in01f80 g773022 ( .a(n_7747), .o(n_7748) );
no02f80 g744851 ( .a(FE_OCP_RBN2615_n_35005), .b(n_34932), .o(n_35060) );
na02f80 g756004 ( .a(n_25160), .b(n_25251), .o(n_25307) );
in01f80 g767245 ( .a(n_13639), .o(n_13640) );
in01f80 g747404 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_2_), .o(n_32615) );
no02f80 g766315 ( .a(n_14333), .b(n_14369), .o(n_14403) );
in01f80 newInst_1691 ( .a(newNet_1690), .o(newNet_1691) );
ao22s80 FE_RC_1176_0 ( .a(FE_OCP_RBN3463_n_7886), .b(FE_OCP_RBN3515_n_8498), .c(FE_OCP_RBN2302_n_7817), .d(n_8498), .o(n_8608) );
no02f80 g747666 ( .a(n_32150), .b(n_32149), .o(n_32151) );
na02f80 g736716 ( .a(n_43313), .b(n_43230), .o(n_43473) );
in01f80 g744702 ( .a(n_35251), .o(n_35252) );
na02f80 g759596 ( .a(n_20549), .b(n_45066), .o(n_20594) );
no02f80 g776784 ( .a(n_4030), .b(FE_OCP_RBN2690_FE_OCPN843_n_3912), .o(n_4115) );
na02f80 g769663 ( .a(n_11314), .b(n_11281), .o(n_11381) );
in01f80 newInst_1021 ( .a(newNet_723), .o(newNet_1021) );
na02f80 g779037 ( .a(n_2123), .b(n_2098), .o(n_2154) );
in01f80 FE_OCP_RBC3037_n_47269 ( .a(n_47269), .o(FE_OCP_RBN3037_n_47269) );
na02f80 g769124 ( .a(n_11511), .b(n_11550), .o(n_11731) );
na02f80 g776448 ( .a(n_4614), .b(n_4619), .o(n_4615) );
no02f80 g756485 ( .a(n_23970), .b(n_23945), .o(n_23967) );
no02f80 g758244 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_19_), .o(n_22846) );
no02f80 g744483 ( .a(n_35444), .b(n_35282), .o(n_35448) );
no02f80 g745224 ( .a(n_34570), .b(n_34569), .o(n_34571) );
no02f80 g738742 ( .a(n_41483), .b(n_41254), .o(n_41687) );
in01f80 newInst_1804 ( .a(newNet_976), .o(newNet_1804) );
na02f80 g770559 ( .a(n_10192), .b(FE_OCP_RBN3597_FE_OCPN1243_n_44460), .o(n_10319) );
no02f80 g772458 ( .a(n_8503), .b(n_8061), .o(n_8517) );
in01f80 g772733 ( .a(n_8291), .o(n_8292) );
in01f80 g774744 ( .a(n_6438), .o(n_6439) );
no02f80 g745947 ( .a(n_35278), .b(n_34777), .o(n_35356) );
in01f80 FE_OCPC968_n_19342 ( .a(FE_OCPN967_n_19342), .o(FE_OCPN968_n_19342) );
in01f80 g761576 ( .a(n_20231), .o(n_22833) );
no02f80 g743624 ( .a(n_36397), .b(n_36011), .o(n_36431) );
na02f80 g744950 ( .a(n_34975), .b(n_34953), .o(n_35077) );
na02f80 g743217 ( .a(n_35506), .b(delay_sub_ln21_unr24_stage9_stallmux_q_4_), .o(n_37175) );
ao12f80 g768984 ( .a(n_11975), .b(n_45685), .c(delay_xor_ln22_unr9_stage4_stallmux_q_11_), .o(n_12017) );
in01f80 g775708 ( .a(n_5545), .o(n_5546) );
in01f80 newInst_2374 ( .a(newNet_2373), .o(newNet_2374) );
na02f80 g751448 ( .a(n_28474), .b(n_28473), .o(n_28475) );
no02f80 FE_RC_2233_0 ( .a(FE_RN_813_0), .b(n_17863), .o(n_17939) );
ao22s80 FE_RC_1389_0 ( .a(n_30545), .b(n_34983), .c(delay_sub_ln23_0_unr22_stage8_stallmux_q), .d(n_34960), .o(n_35107) );
na02f80 g749689 ( .a(n_31412), .b(n_31391), .o(n_31542) );
in01f80 g745688 ( .a(n_34261), .o(n_34297) );
in01f80 g773654 ( .a(n_7848), .o(n_7356) );
na02f80 g746464 ( .a(n_34844), .b(n_34776), .o(n_34845) );
in01f80 g764605 ( .a(n_16179), .o(n_16269) );
na02f80 g763358 ( .a(n_17708), .b(n_17467), .o(n_17709) );
in01f80 newInst_991 ( .a(newNet_647), .o(newNet_991) );
oa12f80 g759085 ( .a(n_21958), .b(n_21909), .c(n_21957), .o(n_21994) );
na02f80 g762125 ( .a(n_18174), .b(n_18173), .o(n_18175) );
in01f80 newInst_691 ( .a(newNet_199), .o(newNet_691) );
in01f80 g779047 ( .a(n_2173), .o(n_2174) );
na02f80 g778675 ( .a(n_2365), .b(n_2929), .o(n_2412) );
no02f80 g764582 ( .a(n_16154), .b(n_16111), .o(n_16112) );
in01f80 newInst_2093 ( .a(newNet_1013), .o(newNet_2093) );
in01f80 FE_OCP_RBC2291_n_2438 ( .a(n_2438), .o(FE_OCP_RBN2291_n_2438) );
na02f80 g743027 ( .a(n_37102), .b(n_36435), .o(n_37103) );
in01f80 newInst_204 ( .a(newNet_17), .o(newNet_204) );
in01f80 FE_OCP_RBC2702_n_4041 ( .a(n_4041), .o(FE_OCP_RBN2702_n_4041) );
oa12f80 g745077 ( .a(n_34241), .b(n_34714), .c(n_34687), .o(n_34715) );
na02f80 g762263 ( .a(n_18582), .b(n_18495), .o(n_19485) );
na02f80 g754809 ( .a(n_25362), .b(n_25361), .o(n_25457) );
ao12f80 g761842 ( .a(n_18704), .b(n_18741), .c(n_17748), .o(n_18743) );
na02f80 g778124 ( .a(n_2873), .b(n_2679), .o(n_2917) );
in01f80 FE_RC_2417_0 ( .a(n_7132), .o(FE_RN_955_0) );
in01f80 g780138 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_21_), .o(n_1177) );
in01f80 g761627 ( .a(n_19607), .o(n_19900) );
in01f80 newInst_788 ( .a(newNet_787), .o(newNet_788) );
no02f80 g777067 ( .a(n_3667), .b(n_3705), .o(n_3742) );
na02f80 g774973 ( .a(n_6165), .b(FE_OCP_RBN2931_n_5307), .o(n_6235) );
na02f80 g745579 ( .a(n_34291), .b(n_34292), .o(n_34344) );
no02f80 g755688 ( .a(n_24372), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24412) );
in01f80 g754703 ( .a(n_26271), .o(n_26690) );
in01f80 g737270 ( .a(n_46939), .o(n_43243) );
na02f80 g748283 ( .a(FE_OCP_RBN3732_n_31819), .b(n_30955), .o(n_32017) );
no02f80 g756009 ( .a(n_25160), .b(n_25250), .o(n_25679) );
ao22s80 FE_RC_260_0 ( .a(n_19264), .b(n_19748), .c(n_19749), .d(n_19301), .o(n_19894) );
na02f80 g742796 ( .a(n_37314), .b(n_37313), .o(n_37315) );
no02f80 g756232 ( .a(n_24122), .b(n_23679), .o(n_24164) );
in01f80 g778274 ( .a(n_2739), .o(n_2740) );
ao12f80 g768849 ( .a(n_11836), .b(n_11835), .c(n_11834), .o(n_12699) );
in01f80 newInst_709 ( .a(newNet_708), .o(newNet_709) );
oa12f80 g759245 ( .a(n_21043), .b(n_21042), .c(n_21041), .o(n_21124) );
no02f80 g776172 ( .a(FE_OCP_RBN2816_n_4459), .b(FE_OCP_RBN2723_n_4219), .o(n_4570) );
in01f80 g755077 ( .a(n_25747), .o(n_25748) );
na02f80 g736757 ( .a(n_43273), .b(n_43260), .o(n_43366) );
na02f80 g738346 ( .a(n_41792), .b(n_41746), .o(n_41816) );
in01f80 newInst_3208 ( .a(newNet_1171), .o(newNet_3208) );
no02f80 g780846 ( .a(n_448), .b(n_447), .o(n_449) );
in01f80 newInst_2179 ( .a(newNet_2178), .o(newNet_2179) );
na02f80 g772588 ( .a(n_8484), .b(n_8424), .o(n_8511) );
no02f80 FE_RC_3472_0 ( .a(FE_RN_1491_0), .b(n_39081), .o(FE_RN_1492_0) );
in01f80 g762107 ( .a(n_18261), .o(n_18262) );
in01f80 g741013 ( .a(n_39139), .o(n_39104) );
in01f80 g742740 ( .a(n_37395), .o(n_37396) );
no02f80 g763284 ( .a(n_17230), .b(n_17229), .o(n_17272) );
no02f80 g779592 ( .a(n_1364), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1406) );
no02f80 FE_RC_2382_0 ( .a(FE_RN_929_0), .b(n_12281), .o(FE_RN_930_0) );
in01f80 g750849 ( .a(n_29115), .o(n_29141) );
na02f80 g767822 ( .a(n_13084), .b(n_12255), .o(n_13381) );
na02f80 g744498 ( .a(n_35444), .b(n_35327), .o(n_35442) );
in01f80 g776063 ( .a(n_4751), .o(n_5988) );
na02f80 g771420 ( .a(n_9140), .b(n_9193), .o(n_9342) );
in01f80 g760875 ( .a(n_19465), .o(n_19466) );
no02f80 g737682 ( .a(FE_OCPN885_n_42216), .b(n_42052), .o(n_42549) );
no02f80 g742000 ( .a(n_38016), .b(n_37980), .o(n_38261) );
in01f80 g758411 ( .a(FE_OCPN1494_n_23398), .o(n_23447) );
in01f80 FE_OCP_RBC2881_n_21272 ( .a(n_21272), .o(FE_OCP_RBN2881_n_21272) );
oa22f80 FE_RC_1669_0 ( .a(n_17584), .b(n_17550), .c(n_17753), .d(n_17475), .o(n_17585) );
na02f80 g737758 ( .a(n_42310), .b(n_42309), .o(n_42311) );
na02f80 g750060 ( .a(n_29869), .b(FE_OCP_RBN2265_n_29033), .o(n_30120) );
oa12f80 g742886 ( .a(n_46254), .b(n_37071), .c(delay_add_ln22_unr23_stage9_stallmux_q_23_), .o(n_37130) );
na02f80 g743938 ( .a(n_36915), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_0_), .o(n_36925) );
in01f80 g744901 ( .a(n_36450), .o(n_36451) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_11_ ( .ck(newNet_593), .d(n_17647), .o(delay_xor_ln22_unr12_stage5_stallmux_q_11_) );
na02f80 FE_RC_814_0 ( .a(FE_RN_245_0), .b(n_29122), .o(n_46960) );
in01f80 newInst_558 ( .a(newNet_557), .o(newNet_558) );
ao12f80 g784611 ( .a(n_42890), .b(n_42869), .c(n_42616), .o(n_46939) );
na02f80 g748877 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_5_), .o(n_32481) );
oa22f80 g776685 ( .a(n_3993), .b(n_3106), .c(n_4017), .d(n_3082), .o(n_4307) );
oa12f80 g761060 ( .a(n_20116), .b(n_20115), .c(n_20114), .o(n_21454) );
no02f80 g761733 ( .a(n_18566), .b(n_18437), .o(n_18681) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_26_ ( .ck(newNet_2271), .d(n_40553), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_) );
na02f80 g749366 ( .a(n_30622), .b(n_30671), .o(n_30944) );
na02f80 g739972 ( .a(n_40295), .b(n_40134), .o(n_40398) );
in01f80 g739693 ( .a(n_40574), .o(n_40585) );
na02f80 g751737 ( .a(FE_OCPN987_n_28402), .b(n_28354), .o(n_28512) );
no02f80 g771160 ( .a(n_9879), .b(n_9817), .o(n_10029) );
ao12f80 g767480 ( .a(n_13185), .b(FE_OCP_RBN2230_n_13141), .c(n_12881), .o(n_13332) );
in01f80 FE_OCP_RBC2760_n_15180 ( .a(n_15180), .o(FE_OCP_RBN2760_n_15180) );
in01f80 g773668 ( .a(n_7341), .o(n_7342) );
no02f80 g739116 ( .a(n_40945), .b(n_40789), .o(n_41017) );
in01f80 FE_OCP_DRV_C1595_n_21458 ( .a(n_21458), .o(FE_OCP_DRV_N1595_n_21458) );
in01f80 g751022 ( .a(n_30001), .o(n_29910) );
ao12f80 g756947 ( .a(n_23747), .b(n_23803), .c(n_23800), .o(n_24194) );
no02f80 g769869 ( .a(n_11074), .b(n_11048), .o(n_11134) );
oa12f80 g767464 ( .a(n_13302), .b(n_13394), .c(n_13357), .o(n_13448) );
ao12f80 g745083 ( .a(n_34849), .b(n_34848), .c(n_34847), .o(n_34947) );
in01f80 newInst_1997 ( .a(newNet_1508), .o(newNet_1997) );
in01f80 FE_OCP_RBC2322_n_2638 ( .a(n_2638), .o(FE_OCP_RBN2322_n_2638) );
na02f80 g749786 ( .a(n_31570), .b(n_31528), .o(n_31627) );
no02f80 FE_RC_185_0 ( .a(FE_RN_62_0), .b(n_354), .o(n_355) );
na02f80 g769180 ( .a(n_11571), .b(n_11570), .o(n_11728) );
na02f80 g778527 ( .a(n_2551), .b(delay_add_ln22_unr2_stage2_stallmux_q_24_), .o(n_2630) );
in01f80 g737232 ( .a(n_42968), .o(n_42980) );
ao12f80 g774052 ( .a(n_7195), .b(n_7172), .c(delay_xor_ln22_unr6_stage3_stallmux_q_21_), .o(n_7328) );
no03m80 g773449 ( .a(n_7515), .b(n_7529), .c(n_6828), .o(n_7624) );
in01f80 FE_OCP_RBC2514_n_8739 ( .a(n_8739), .o(FE_OCP_RBN2514_n_8739) );
no02f80 g749311 ( .a(n_30655), .b(n_30343), .o(n_30676) );
ao12f80 g757524 ( .a(n_22342), .b(n_22686), .c(n_22220), .o(n_22687) );
in01f80 g771215 ( .a(n_9757), .o(n_9758) );
oa22f80 FE_RC_2650_0 ( .a(n_2759), .b(FE_OCP_RBN2576_n_47017), .c(n_3615), .d(n_47017), .o(n_3761) );
in01f80 newInst_387 ( .a(newNet_30), .o(newNet_387) );
in01f80 FE_RC_1310_0 ( .a(n_3613), .o(FE_RN_384_0) );
in01f80 g755693 ( .a(n_24467), .o(n_24468) );
no02f80 g759946 ( .a(n_21406), .b(n_21625), .o(n_21772) );
oa12f80 g764671 ( .a(n_16481), .b(n_16480), .c(n_16479), .o(n_16523) );
in01f80 g778968 ( .a(n_2151), .o(n_2152) );
in01f80 g742073 ( .a(n_38328), .o(n_38329) );
no02f80 g753889 ( .a(n_26185), .b(n_24591), .o(n_26338) );
in01f80 g755733 ( .a(n_25311), .o(n_25312) );
na02f80 g773585 ( .a(n_7417), .b(n_7416), .o(n_7418) );
ao12f80 g745165 ( .a(n_34220), .b(n_34542), .c(n_34203), .o(n_34663) );
in01f80 g758289 ( .a(n_22213), .o(n_22253) );
in01f80 g780311 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_8_), .o(n_946) );
na02f80 g768280 ( .a(n_12561), .b(n_12560), .o(n_12562) );
oa12f80 g769104 ( .a(n_45685), .b(n_12076), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n_12168) );
na02f80 g750565 ( .a(n_29401), .b(n_29241), .o(n_29481) );
no02f80 g761693 ( .a(n_18824), .b(n_18713), .o(n_18825) );
ao22s80 FE_RC_1265_0 ( .a(n_2905), .b(n_3595), .c(n_2904), .d(n_3636), .o(n_3807) );
na02f80 g744149 ( .a(n_35776), .b(FE_OCP_RBN2645_n_34980), .o(n_35819) );
oa12f80 g751529 ( .a(n_29253), .b(n_29252), .c(n_29251), .o(n_29359) );
oa12f80 g738200 ( .a(n_41964), .b(n_41977), .c(n_41963), .o(n_42500) );
oa22f80 g739856 ( .a(n_40377), .b(n_40386), .c(n_40378), .d(n_40387), .o(n_40440) );
no02f80 FE_RC_364_0 ( .a(FE_RN_108_0), .b(FE_RN_109_0), .o(FE_RN_110_0) );
no02f80 g765201 ( .a(n_15270), .b(n_15269), .o(n_15271) );
na02f80 g768408 ( .a(n_12383), .b(n_12376), .o(n_12464) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_6_ ( .ck(newNet_2238), .d(n_40198), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_) );
in01f80 g737856 ( .a(n_42620), .o(n_42621) );
in01f80 newInst_2998 ( .a(newNet_1599), .o(newNet_2998) );
na02f80 g775630 ( .a(n_5459), .b(n_5424), .o(n_5497) );
no02f80 g740227 ( .a(n_40098), .b(FE_OCP_RBN3022_n_39942), .o(n_40251) );
oa12f80 g772986 ( .a(n_7407), .b(n_7754), .c(n_7388), .o(n_7938) );
in01f80 g741707 ( .a(n_38573), .o(n_38550) );
na02f80 g748242 ( .a(n_31783), .b(n_31804), .o(n_31847) );
na02f80 g756934 ( .a(n_23700), .b(n_23810), .o(n_23867) );
no02f80 FE_RC_2638_0 ( .a(n_2288), .b(n_2289), .o(FE_RN_1100_0) );
in01f80 g771654 ( .a(n_8939), .o(n_8940) );
no02f80 g743795 ( .a(n_35923), .b(n_35879), .o(n_36015) );
na02f80 g762337 ( .a(n_18050), .b(n_18006), .o(n_18075) );
in01f80 g768028 ( .a(n_13621), .o(n_12917) );
na02f80 g766814 ( .a(n_14346), .b(n_14351), .o(n_14431) );
na02f80 g773471 ( .a(n_7500), .b(delay_add_ln22_unr5_stage3_stallmux_q_24_), .o(n_7530) );
in01f80 g767760 ( .a(n_13099), .o(n_13173) );
oa12f80 g757268 ( .a(n_22732), .b(n_23468), .c(n_22843), .o(n_23488) );
na02f80 g768546 ( .a(n_12316), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .o(n_12389) );
na02f80 g778988 ( .a(n_2107), .b(n_1952), .o(n_2158) );
in01f80 FE_OCP_RBC2907_n_16230 ( .a(n_16230), .o(FE_OCP_RBN2907_n_16230) );
in01f80 g740394 ( .a(n_40206), .o(n_40207) );
na02f80 g739305 ( .a(n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_18_), .o(n_40790) );
na02f80 FE_RC_1790_0 ( .a(n_7016), .b(n_7209), .o(FE_RN_527_0) );
in01f80 FE_OCPC1525_n_26587 ( .a(n_26587), .o(FE_OCPN1525_n_26587) );
no02f80 g755273 ( .a(n_24986), .b(n_24965), .o(n_25067) );
no02f80 g764936 ( .a(n_15393), .b(n_15354), .o(n_15557) );
in01f80 newInst_761 ( .a(newNet_300), .o(newNet_761) );
in01f80 g769095 ( .a(n_11713), .o(n_11714) );
in01f80 newInst_518 ( .a(newNet_517), .o(newNet_518) );
no02f80 g773664 ( .a(n_7323), .b(n_7143), .o(n_7358) );
in01f80 FE_OCP_RBC2512_n_19884 ( .a(n_19884), .o(FE_OCP_RBN2512_n_19884) );
no02f80 g768097 ( .a(n_12670), .b(n_12086), .o(n_12741) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_2_ ( .ck(newNet_305), .d(n_1335), .o(delay_xor_ln22_unr3_stage2_stallmux_q_2_) );
in01f80 g749589 ( .a(n_30424), .o(n_30425) );
in01f80 g765310 ( .a(n_15959), .o(n_15960) );
na02f80 g771224 ( .a(n_9535), .b(FE_OCPN903_n_44581), .o(n_9635) );
no02f80 g749705 ( .a(n_31147), .b(n_31088), .o(n_31191) );
no02f80 FE_RC_2788_0 ( .a(n_34224), .b(n_34164), .o(FE_RN_1191_0) );
in01f80 g768961 ( .a(n_11788), .o(n_11789) );
in01f80 newInst_701 ( .a(newNet_135), .o(newNet_701) );
oa22f80 g746876 ( .a(FE_OCP_RBN3389_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_17_), .c(n_33108), .d(n_32171), .o(n_33519) );
no02f80 g774285 ( .a(n_6863), .b(n_6850), .o(n_6942) );
na02f80 FE_RC_141_0 ( .a(n_18050), .b(n_18226), .o(FE_RN_40_0) );
na02f80 g743096 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_29_), .o(n_37150) );
ao12f80 g757906 ( .a(n_23055), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n_23568) );
no02f80 g774819 ( .a(n_6247), .b(n_6213), .o(n_6308) );
no02f80 FE_RC_2265_0 ( .a(FE_RN_840_0), .b(n_25119), .o(FE_RN_841_0) );
in01f80 g742969 ( .a(n_36975), .o(n_36976) );
no02f80 g737564 ( .a(n_42261), .b(n_42285), .o(n_42317) );
no02f80 g761078 ( .a(n_19141), .b(FE_OCP_RBN1687_n_18986), .o(n_19209) );
ao12f80 g763500 ( .a(n_16777), .b(n_16784), .c(n_16752), .o(n_16904) );
no02f80 g767594 ( .a(n_12950), .b(n_12797), .o(n_13290) );
na02f80 g772364 ( .a(n_8571), .b(n_7957), .o(n_8660) );
na02f80 g743186 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_4_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .o(n_36936) );
in01f80 FE_RC_3817_0 ( .a(n_24562), .o(FE_RN_1665_0) );
in01f80 g736851 ( .a(n_43545), .o(n_43546) );
in01f80 newInst_1203 ( .a(newNet_922), .o(newNet_1203) );
in01f80 g739024 ( .a(n_41545), .o(n_41180) );
ao12f80 g741743 ( .a(n_38428), .b(n_38427), .c(n_38426), .o(n_38498) );
in01f80 g765882 ( .a(n_14901), .o(n_14902) );
in01f80 g780126 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_22_), .o(n_2379) );
in01f80 g747422 ( .a(n_32634), .o(n_32621) );
no02f80 g741178 ( .a(FE_OCP_RBN2637_n_38806), .b(n_38884), .o(n_39081) );
in01f80 g778206 ( .a(n_2861), .o(n_2862) );
in01f80 g745051 ( .a(n_35785), .o(n_34772) );
no02f80 g748646 ( .a(n_32608), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n_32609) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_7_ ( .ck(newNet_3474), .d(n_21702), .o(delay_add_ln22_unr14_stage6_stallmux_q_7_) );
in01f80 g765547 ( .a(n_15144), .o(n_15182) );
in01f80 g770491 ( .a(n_10243), .o(n_10320) );
ao12f80 g757280 ( .a(n_23449), .b(n_23468), .c(n_23448), .o(n_23804) );
in01f80 fopt783584 ( .a(n_6328), .o(n_45214) );
na02f80 g756022 ( .a(n_25139), .b(n_25135), .o(n_25253) );
na02f80 g777009 ( .a(n_3842), .b(n_3928), .o(n_4006) );
oa12f80 g759027 ( .a(n_21528), .b(n_21527), .c(n_21526), .o(n_21602) );
ao22s80 FE_RC_249_0 ( .a(n_14747), .b(n_14821), .c(FE_OCPN3767_n_14439), .d(n_14746), .o(n_14865) );
na02f80 g745056 ( .a(n_34730), .b(n_34755), .o(n_34828) );
oa22f80 g752600 ( .a(n_27555), .b(n_27542), .c(n_27556), .d(n_27543), .o(n_27584) );
ao12f80 g773866 ( .a(n_6989), .b(n_6997), .c(n_6988), .o(n_7053) );
in01f80 newInst_2425 ( .a(newNet_197), .o(newNet_2425) );
na02f80 g779554 ( .a(n_1366), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1455) );
oa22f80 g739736 ( .a(n_40496), .b(n_40408), .c(n_40497), .d(n_40407), .o(n_40530) );
na02f80 g758788 ( .a(n_21556), .b(n_21554), .o(n_21588) );
in01f80 newInst_891 ( .a(newNet_890), .o(newNet_891) );
in01f80 g741296 ( .a(n_38906), .o(n_38994) );
in01f80 FE_OCP_RBC3701_n_31064 ( .a(n_31064), .o(FE_OCP_RBN3701_n_31064) );
in01f80 FE_OCP_RBC2466_n_8393 ( .a(n_8393), .o(FE_OCP_RBN2466_n_8393) );
na02f80 g746037 ( .a(n_33828), .b(n_33697), .o(n_33859) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_9_ ( .ck(newNet_1356), .d(n_36454), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_9_) );
ao12f80 g746529 ( .a(n_34473), .b(n_34640), .c(n_34582), .o(n_34641) );
in01f80 g753527 ( .a(n_26839), .o(n_26840) );
na02f80 g752007 ( .a(n_28897), .b(n_28203), .o(n_29201) );
in01f80 g746239 ( .a(n_33595), .o(n_33596) );
in01f80 g748842 ( .a(n_31058), .o(n_31059) );
na02f80 g753161 ( .a(n_27420), .b(n_27456), .o(n_27544) );
no02f80 g755295 ( .a(n_25065), .b(n_25064), .o(n_25246) );
no02f80 g777277 ( .a(n_3698), .b(n_3697), .o(n_3699) );
in01f80 FE_OCPC848_n_3597 ( .a(FE_OCPN847_n_3597), .o(FE_OCPN848_n_3597) );
no02f80 g743948 ( .a(n_36098), .b(n_36148), .o(n_36199) );
in01f80 fopt782682 ( .a(n_44084), .o(n_44083) );
in01f80 g739680 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n_40545) );
no02f80 g753327 ( .a(n_27100), .b(n_27099), .o(n_27151) );
in01f80 newInst_1734 ( .a(newNet_1733), .o(newNet_1734) );
in01f80 g774353 ( .a(n_6570), .o(n_6831) );
in01f80 newInst_803 ( .a(newNet_273), .o(newNet_803) );
na02f80 g780613 ( .a(n_662), .b(n_553), .o(n_664) );
na02f80 g756872 ( .a(n_24028), .b(n_23803), .o(n_24091) );
in01f80 g767679 ( .a(n_13463), .o(n_13464) );
no02f80 g767780 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_23_), .o(n_12807) );
oa12f80 g754976 ( .a(n_25108), .b(n_25118), .c(n_25107), .o(n_26801) );
oa12f80 g740501 ( .a(n_39735), .b(n_39734), .c(FE_OCP_RBN2866_n_39640), .o(n_39736) );
no02f80 g754260 ( .a(n_26717), .b(n_26454), .o(n_26795) );
in01f80 fopt784019 ( .a(n_45755), .o(n_45754) );
in01f80 FE_RC_2463_0 ( .a(n_13898), .o(FE_RN_989_0) );
in01f80 g751427 ( .a(n_28476), .o(n_29737) );
in01f80 newInst_2862 ( .a(newNet_2861), .o(newNet_2862) );
no02f80 g774314 ( .a(FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .o(n_6716) );
no02f80 FE_RC_502_0 ( .a(FE_RN_152_0), .b(n_23329), .o(n_23315) );
na02f80 g745411 ( .a(FE_OCP_RBN3697_n_35543), .b(n_35559), .o(n_35560) );
in01f80 g748331 ( .a(n_31953), .o(n_31861) );
oa12f80 g759726 ( .a(n_20637), .b(n_20636), .c(n_20635), .o(n_20715) );
ao12f80 g756522 ( .a(n_23874), .b(n_23783), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_), .o(n_23941) );
no02f80 g778129 ( .a(n_2932), .b(n_2774), .o(n_2950) );
no02f80 g744848 ( .a(n_35092), .b(n_30633), .o(n_35117) );
na02f80 g775094 ( .a(n_6026), .b(n_5792), .o(n_6053) );
no02f80 g761003 ( .a(n_19184), .b(n_18425), .o(n_19185) );
in01f80 newInst_89 ( .a(newNet_37), .o(newNet_89) );
in01f80 newInst_2304 ( .a(newNet_2303), .o(newNet_2304) );
in01f80 g744814 ( .a(n_36477), .o(n_36478) );
na02f80 g754938 ( .a(n_25884), .b(n_25883), .o(n_25885) );
na02f80 g744612 ( .a(n_36603), .b(n_36283), .o(n_36623) );
na02f80 g768029 ( .a(n_12910), .b(n_12909), .o(n_13621) );
in01f80 g754496 ( .a(n_26905), .o(n_26906) );
no02f80 g761545 ( .a(n_18758), .b(n_18264), .o(n_18864) );
na02f80 g763831 ( .a(n_17421), .b(n_17300), .o(n_17980) );
no02f80 g743106 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_19_), .o(n_37046) );
in01f80 FE_RC_3375_0 ( .a(n_18629), .o(FE_RN_1465_0) );
in01f80 g769743 ( .a(n_11223), .o(n_11256) );
no02f80 g738590 ( .a(n_41560), .b(n_41687), .o(n_42141) );
no02f80 g768344 ( .a(n_12590), .b(n_12581), .o(n_12582) );
no02f80 g744153 ( .a(n_36063), .b(n_36062), .o(n_36064) );
na02f80 g747244 ( .a(n_32655), .b(n_32654), .o(n_32668) );
in01f80 g757355 ( .a(n_23124), .o(n_23125) );
in01f80 g774927 ( .a(n_6191), .o(n_6192) );
in01f80 FE_OCP_RBC2903_n_44174 ( .a(FE_OCP_RBN2901_n_44174), .o(FE_OCP_RBN2903_n_44174) );
na02f80 g767043 ( .a(FE_OCP_RBN3529_n_13765), .b(n_13893), .o(n_13973) );
in01f80 FE_OCPC3179_FE_OCP_RBN2744_n_15319 ( .a(FE_OCP_RBN2744_n_15319), .o(FE_OCPN3179_FE_OCP_RBN2744_n_15319) );
in01f80 g751474 ( .a(n_28601), .o(n_28602) );
na02f80 g738024 ( .a(n_42144), .b(n_42196), .o(n_42146) );
na02f80 g759428 ( .a(n_20937), .b(n_20570), .o(n_20998) );
in01f80 FE_RC_1516_0 ( .a(n_31738), .o(FE_RN_426_0) );
no02f80 g747628 ( .a(n_33297), .b(n_33241), .o(n_33361) );
ao12f80 g771700 ( .a(n_7584), .b(n_44057), .c(n_8699), .o(n_8746) );
no02f80 g755049 ( .a(n_25445), .b(n_25375), .o(n_25479) );
in01f80 g738932 ( .a(n_41217), .o(n_41482) );
in01f80 newInst_2248 ( .a(newNet_2247), .o(newNet_2248) );
no02f80 g780415 ( .a(n_803), .b(n_802), .o(n_1208) );
no02f80 g752187 ( .a(n_28096), .b(n_28095), .o(n_28061) );
in01f80 FE_OCP_RBC2737_n_15300 ( .a(n_15300), .o(FE_OCP_RBN2737_n_15300) );
in01f80 g750872 ( .a(n_29091), .o(n_29111) );
oa12f80 g770343 ( .a(n_10658), .b(n_10689), .c(n_10657), .o(n_10717) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_5_ ( .ck(newNet_696), .d(n_46176), .o(delay_xor_ln21_unr6_stage3_stallmux_q_5_) );
in01f80 newInst_495 ( .a(newNet_494), .o(newNet_495) );
in01f80 g781329 ( .a(n_69), .o(n_155) );
no02f80 g775869 ( .a(n_5283), .b(n_5228), .o(n_5229) );
oa22f80 FE_RC_885_0 ( .a(n_24757), .b(n_24899), .c(n_24756), .d(n_24898), .o(n_25023) );
no02f80 g773091 ( .a(n_7980), .b(n_8012), .o(n_8013) );
no02f80 g777108 ( .a(n_3677), .b(FE_OCP_RBN2582_n_3734), .o(n_3777) );
in01f80 g748883 ( .a(n_32416), .o(n_32486) );
in01f80 g764157 ( .a(n_16889), .o(n_16890) );
in01f80 newInst_2605 ( .a(newNet_2604), .o(newNet_2605) );
in01f80 FE_OCP_RBC2502_n_13896 ( .a(FE_OCP_RBN3528_n_13765), .o(FE_OCP_RBN2502_n_13896) );
in01f80 g744449 ( .a(n_35512), .o(n_35513) );
in01f80 newInst_3273 ( .a(newNet_1742), .o(newNet_3273) );
in01f80 FE_OCPC897_n_44776 ( .a(FE_OCPN896_n_44776), .o(FE_OCPN897_n_44776) );
in01f80 FE_OCP_RBC2185_FE_RN_464_0 ( .a(FE_RN_464_0), .o(FE_OCP_RBN2185_FE_RN_464_0) );
ao12f80 g739198 ( .a(n_45153), .b(n_40888), .c(n_40891), .o(n_40939) );
in01f80 g773180 ( .a(n_7665), .o(n_7666) );
in01f80 g749944 ( .a(n_30369), .o(n_30370) );
na02f80 g775983 ( .a(n_5243), .b(n_5242), .o(n_5274) );
na02f80 g761011 ( .a(n_19206), .b(n_17900), .o(n_19253) );
na02f80 FE_RC_4023_0 ( .a(FE_RN_1747_0), .b(n_25912), .o(FE_RN_1573_0) );
oa12f80 g754594 ( .a(n_26601), .b(n_26896), .c(n_26643), .o(n_26924) );
na02f80 g739353 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n_41040) );
ao12f80 g750033 ( .a(n_30903), .b(n_30925), .c(n_30902), .o(n_30970) );
in01f80 fopt782732 ( .a(n_29316), .o(n_44139) );
ao22s80 g756220 ( .a(n_24093), .b(FE_OCPN1780_n_24097), .c(n_24098), .d(n_22752), .o(n_24218) );
ao12f80 g742161 ( .a(n_37892), .b(n_44887), .c(n_37852), .o(n_38382) );
na02f80 g741317 ( .a(FE_OCP_RBN2546_n_44944), .b(n_38529), .o(n_39131) );
no02f80 g770200 ( .a(n_10595), .b(n_10553), .o(n_10676) );
no02f80 g747218 ( .a(n_32718), .b(n_32669), .o(n_32758) );
in01f80 g765952 ( .a(n_14790), .o(n_14791) );
in01f80 FE_OCP_RBC2885_n_35517 ( .a(n_35517), .o(FE_OCP_RBN2885_n_35517) );
na02f80 g755806 ( .a(n_25259), .b(n_25160), .o(n_25221) );
ao12f80 g772508 ( .a(n_8432), .b(n_8431), .c(n_8430), .o(n_9587) );
na02f80 g775328 ( .a(n_5888), .b(n_5649), .o(n_5901) );
in01f80 g743686 ( .a(n_36347), .o(n_36348) );
na02f80 g738209 ( .a(n_41953), .b(n_41952), .o(n_41954) );
oa12f80 g765799 ( .a(n_14353), .b(n_15289), .c(n_14491), .o(n_15446) );
no02f80 g777362 ( .a(n_4556), .b(n_4693), .o(n_4721) );
in01f80 g761749 ( .a(n_18600), .o(n_18605) );
oa22f80 FE_RC_4137_0 ( .a(n_22819), .b(n_22801), .c(n_22793), .d(n_22792), .o(n_22893) );
in01f80 g771784 ( .a(n_8966), .o(n_8967) );
na02f80 g759510 ( .a(n_20878), .b(n_20842), .o(n_20966) );
in01f80 newInst_1453 ( .a(newNet_1452), .o(newNet_1453) );
na02f80 g772925 ( .a(n_7836), .b(FE_OCPN1396_n_7881), .o(n_7882) );
na02f80 g759103 ( .a(n_21191), .b(n_21192), .o(n_21224) );
na02f80 g764375 ( .a(n_16190), .b(n_14805), .o(n_16283) );
no02f80 g764424 ( .a(n_16169), .b(n_14420), .o(n_16168) );
in01f80 g779346 ( .a(n_1653), .o(n_1654) );
no02f80 g746485 ( .a(n_34668), .b(n_34698), .o(n_34742) );
in01f80 newInst_3203 ( .a(newNet_3202), .o(newNet_3203) );
in01f80 newInst_1946 ( .a(newNet_1945), .o(newNet_1946) );
in01f80 g762724 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_26_), .o(n_17806) );
in01f80 FE_RC_2340_0 ( .a(n_11756), .o(FE_RN_896_0) );
in01f80 g767395 ( .a(n_13453), .o(n_13404) );
oa12f80 g765109 ( .a(n_16258), .b(n_16175), .c(n_15874), .o(n_16308) );
oa12f80 g750774 ( .a(n_29291), .b(n_29313), .c(n_29290), .o(n_29364) );
in01f80 g776367 ( .a(n_4774), .o(n_4821) );
no02f80 g739080 ( .a(n_41444), .b(n_41028), .o(n_41063) );
in01f80 g745766 ( .a(n_34180), .o(n_34181) );
no02f80 g769996 ( .a(n_10934), .b(n_10954), .o(n_11055) );
in01f80 FE_RC_52_0 ( .a(n_4140), .o(FE_RN_12_0) );
no02f80 g745428 ( .a(FE_OCP_RBN2993_n_35539), .b(n_35217), .o(n_36154) );
in01f80 g758727 ( .a(n_22395), .o(n_22426) );
oa22f80 g749170 ( .a(n_32174), .b(n_31389), .c(n_32175), .d(n_31388), .o(n_32247) );
in01f80 g775587 ( .a(n_5791), .o(n_5792) );
na02f80 g759934 ( .a(n_21374), .b(n_21371), .o(n_21519) );
in01f80 g738825 ( .a(n_41357), .o(n_41358) );
in01f80 g771807 ( .a(n_8964), .o(n_8965) );
oa12f80 g780078 ( .a(n_1214), .b(n_1213), .c(n_1212), .o(n_1219) );
in01f80 newInst_2526 ( .a(newNet_2525), .o(newNet_2526) );
in01f80 newInst_2495 ( .a(newNet_852), .o(newNet_2495) );
na02f80 g745977 ( .a(n_34033), .b(n_33981), .o(n_34064) );
in01f80 g755300 ( .a(n_24921), .o(n_24922) );
in01f80 g756569 ( .a(n_23632), .o(n_23633) );
no02f80 FE_RC_1740_0 ( .a(FE_RN_485_0), .b(FE_RN_486_0), .o(FE_RN_487_0) );
na02f80 g766689 ( .a(n_13779), .b(n_13238), .o(n_13838) );
na02f80 g748977 ( .a(n_31127), .b(n_27246), .o(n_31131) );
in01f80 FE_OCPC953_n_41540 ( .a(FE_OCPN951_n_41540), .o(FE_OCPN953_n_41540) );
in01f80 g780368 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_2_), .o(n_756) );
no02f80 g739393 ( .a(n_45155), .b(n_40340), .o(n_40919) );
na02f80 g776110 ( .a(n_4995), .b(n_4596), .o(n_5046) );
na02f80 g738722 ( .a(n_41435), .b(n_41447), .o(n_41485) );
oa12f80 g768239 ( .a(n_12588), .b(n_12591), .c(n_12587), .o(n_13721) );
in01f80 g760500 ( .a(n_20059), .o(n_20060) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_17_ ( .ck(newNet_2575), .d(n_27584), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_17_) );
no02f80 FE_RC_3142_0 ( .a(FE_RN_1394_0), .b(n_16622), .o(n_16682) );
na02f80 g748110 ( .a(n_31990), .b(n_47274), .o(n_32023) );
no02f80 g748137 ( .a(n_31953), .b(n_32103), .o(n_32104) );
oa22f80 g781277 ( .a(n_46055), .b(beta_12), .c(n_7), .d(n_27), .o(n_210) );
na02f80 g780469 ( .a(n_855), .b(n_759), .o(n_804) );
in01f80 g762816 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_24_), .o(n_18329) );
na02f80 g776792 ( .a(n_4212), .b(n_4211), .o(n_4365) );
na02f80 g779367 ( .a(n_1571), .b(n_1107), .o(n_1656) );
na02f80 g736864 ( .a(n_43343), .b(n_43455), .o(n_43541) );
na02f80 g764950 ( .a(n_15387), .b(FE_OCPN1007_n_13962), .o(n_15437) );
ao12f80 g765058 ( .a(n_15239), .b(n_15276), .c(n_15205), .o(n_15385) );
in01f80 FE_RC_3255_0 ( .a(FE_RN_1436_0), .o(FE_RN_1435_0) );
na02f80 FE_RC_582_0 ( .a(FE_RN_177_0), .b(FE_RN_178_0), .o(FE_RN_179_0) );
no02f80 g745655 ( .a(n_35454), .b(n_34841), .o(n_35477) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_2_ ( .ck(newNet_452), .d(n_27687), .o(delay_xor_ln22_unr18_stage7_stallmux_q_2_) );
in01f80 g760360 ( .a(n_20214), .o(n_20222) );
in01f80 g737367 ( .a(n_42956), .o(n_42878) );
ao12f80 g756631 ( .a(n_23559), .b(n_23558), .c(n_23557), .o(n_23627) );
in01f80 FE_OFC2_n_43918 ( .a(FE_OFN0_n_43918), .o(FE_OFN2_n_43918) );
in01f80 FE_OCP_RBC2511_n_19884 ( .a(n_19884), .o(FE_OCP_RBN2511_n_19884) );
na02f80 g751793 ( .a(n_28299), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_8_), .o(n_28316) );
in01f80 g763415 ( .a(n_16910), .o(n_16911) );
no02f80 g745962 ( .a(n_34061), .b(n_34060), .o(n_34062) );
no02f80 g776165 ( .a(n_4861), .b(n_4476), .o(n_4941) );
in01f80 g768795 ( .a(n_12092), .o(n_12093) );
in01f80 FE_OCP_RBC2103_n_44962 ( .a(FE_OCP_RBN3334_n_44962), .o(FE_OCP_RBN2103_n_44962) );
in01f80 FE_OCPC997_n_44460 ( .a(FE_OCP_RBN3573_n_44563), .o(FE_OCPN997_n_44460) );
na02f80 g746536 ( .a(n_34775), .b(n_34776), .o(n_34806) );
ao12f80 g759579 ( .a(n_20841), .b(n_20877), .c(n_20876), .o(n_20961) );
in01f80 newInst_2315 ( .a(newNet_2314), .o(newNet_2315) );
oa12f80 g748617 ( .a(n_31441), .b(n_31438), .c(n_31356), .o(n_31544) );
na02f80 FE_RC_2784_0 ( .a(n_18140), .b(n_19599), .o(FE_RN_1188_0) );
in01f80 g766276 ( .a(n_14447), .o(n_14408) );
in01f80 FE_RC_765_0 ( .a(n_33213), .o(FE_RN_237_0) );
no02f80 g771749 ( .a(n_9830), .b(n_9876), .o(n_9915) );
in01f80 g743358 ( .a(n_36675), .o(n_36676) );
na02f80 FE_RC_3132_0 ( .a(n_22064), .b(n_22154), .o(FE_RN_1388_0) );
in01f80 g744928 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_7_), .o(n_36784) );
na02f80 g769729 ( .a(n_11238), .b(n_11044), .o(n_11270) );
oa22f80 FE_RC_2529_0 ( .a(n_37141), .b(n_37461), .c(n_37140), .d(n_37462), .o(n_37581) );
no02f80 g769612 ( .a(n_11366), .b(FE_OCP_RBN3063_n_11325), .o(n_11387) );
na02f80 g775628 ( .a(n_5627), .b(n_4289), .o(n_5728) );
in01f80 g754206 ( .a(n_26077), .o(n_26078) );
oa12f80 g760675 ( .a(n_19721), .b(n_19720), .c(n_19719), .o(n_21493) );
ao12f80 g746717 ( .a(n_33111), .b(n_33145), .c(n_33110), .o(n_33968) );
na02f80 g740915 ( .a(n_39284), .b(n_39268), .o(n_39341) );
in01f80 newInst_682 ( .a(newNet_681), .o(newNet_682) );
in01f80 newInst_1420 ( .a(newNet_1321), .o(newNet_1420) );
ao12f80 g764214 ( .a(n_15928), .b(n_16798), .c(n_15922), .o(n_16816) );
in01f80 g765936 ( .a(n_14851), .o(n_14795) );
no02f80 g774489 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_7_), .o(n_6683) );
na02f80 g740169 ( .a(FE_OCP_RBN3719_n_39913), .b(n_39978), .o(n_40181) );
ao12f80 g784436 ( .a(n_46210), .b(n_46204), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_22_), .o(n_46248) );
na02f80 g773503 ( .a(n_7496), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .o(n_7536) );
ao12f80 g736476 ( .a(n_43372), .b(FE_OCP_RBN3110_n_43711), .c(n_43273), .o(n_43750) );
in01f80 g777113 ( .a(n_4058), .o(n_4059) );
no02f80 g780685 ( .a(n_657), .b(n_655), .o(n_656) );
no02f80 FE_RC_3493_0 ( .a(n_12709), .b(n_12902), .o(FE_RN_1506_0) );
in01f80 FE_OCP_RBC3270_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3270_n_45224) );
no02f80 g752010 ( .a(n_28073), .b(n_28068), .o(n_28192) );
na03f80 FE_RC_1872_0 ( .a(n_32439), .b(FE_RN_578_0), .c(n_32641), .o(n_32699) );
in01f80 g761345 ( .a(n_18984), .o(n_18985) );
no02f80 g762869 ( .a(n_17797), .b(n_17796), .o(n_17798) );
in01f80 FE_OCP_RBC3370_n_32436 ( .a(FE_OCP_RBN3368_n_32436), .o(FE_OCP_RBN3370_n_32436) );
no02f80 FE_RC_4044_0 ( .a(FE_RN_1757_0), .b(n_21503), .o(n_21659) );
in01f80 newInst_2599 ( .a(newNet_2598), .o(newNet_2599) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_13_ ( .ck(newNet_1253), .d(n_5498), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_) );
in01f80 FE_OCP_RBC2816_n_4459 ( .a(n_4459), .o(FE_OCP_RBN2816_n_4459) );
in01f80 newInst_1970 ( .a(newNet_1969), .o(newNet_1970) );
in01f80 g757050 ( .a(n_23808), .o(n_23778) );
na02f80 g741513 ( .a(n_38704), .b(n_38695), .o(n_38734) );
no02f80 g772951 ( .a(n_7838), .b(n_7793), .o(n_7974) );
na02f80 g761166 ( .a(n_20015), .b(n_20053), .o(n_20054) );
in01f80 newInst_1964 ( .a(newNet_1901), .o(newNet_1964) );
na02f80 g766117 ( .a(n_14682), .b(n_14681), .o(n_14706) );
in01f80 g742923 ( .a(n_37219), .o(n_37220) );
no02f80 g754468 ( .a(n_25675), .b(n_25459), .o(n_25726) );
in01f80 g759691 ( .a(n_20719), .o(n_20720) );
na02f80 g776251 ( .a(n_47006), .b(n_47341), .o(n_5017) );
oa12f80 g746112 ( .a(n_33776), .b(n_33775), .c(n_33774), .o(n_35312) );
no02f80 g765636 ( .a(n_15446), .b(n_15398), .o(n_15399) );
na02f80 g767072 ( .a(n_13591), .b(n_13590), .o(n_13618) );
ao12f80 g741716 ( .a(n_38503), .b(n_38502), .c(n_38501), .o(n_38919) );
in01f80 g749559 ( .a(n_30492), .o(n_30507) );
no02f80 g779185 ( .a(n_1880), .b(n_1909), .o(n_2487) );
na02f80 g757057 ( .a(n_23671), .b(n_23670), .o(n_23722) );
in01f80 newInst_3292 ( .a(newNet_1578), .o(newNet_3292) );
in01f80 g776074 ( .a(n_5056), .o(n_5057) );
no02f80 g743339 ( .a(n_36704), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36735) );
in01f80 FE_OCP_RBC2139_n_17547 ( .a(n_17547), .o(FE_OCP_RBN2139_n_17547) );
in01f80 g736875 ( .a(n_43605), .o(n_43606) );
no02f80 g741337 ( .a(FE_OCP_RBN2553_n_44921), .b(n_38518), .o(n_38973) );
no02f80 g764623 ( .a(n_15861), .b(n_14588), .o(n_15917) );
no02f80 g761942 ( .a(n_18284), .b(n_17773), .o(n_18548) );
in01f80 g740409 ( .a(n_40030), .o(n_40133) );
in01f80 newInst_2958 ( .a(newNet_271), .o(newNet_2958) );
in01f80 newInst_1492 ( .a(newNet_1491), .o(newNet_1492) );
na02f80 g748937 ( .a(n_31101), .b(n_27366), .o(n_31200) );
no04s80 FE_RC_1288_0 ( .a(n_3041), .b(n_3138), .c(n_3170), .d(n_3237), .o(n_3292) );
na02f80 g740358 ( .a(n_39741), .b(n_39740), .o(n_39753) );
in01f80 g779494 ( .a(n_1436), .o(n_1437) );
na02f80 g749573 ( .a(n_30302), .b(n_30046), .o(n_30354) );
ao22s80 g768855 ( .a(n_44355), .b(n_11714), .c(n_44354), .d(n_11713), .o(n_12058) );
ao12f80 g752113 ( .a(n_28157), .b(n_28636), .c(n_28174), .o(n_28751) );
in01f80 g739044 ( .a(n_41124), .o(n_41501) );
no02f80 g749031 ( .a(n_31075), .b(n_31074), .o(n_31076) );
in01f80 g765676 ( .a(n_15664), .o(n_15719) );
na02f80 g745457 ( .a(n_34352), .b(FE_OCP_RBN2471_n_34285), .o(n_34411) );
no02f80 g752298 ( .a(n_28092), .b(n_27891), .o(n_27964) );
in01f80 newInst_879 ( .a(newNet_85), .o(newNet_879) );
in01f80 g739985 ( .a(n_39987), .o(n_40024) );
no02f80 g743644 ( .a(n_37477), .b(n_46239), .o(n_37478) );
in01f80 g759216 ( .a(n_20983), .o(n_21014) );
no02f80 g757664 ( .a(n_23221), .b(n_22764), .o(n_23242) );
in01f80 FE_OCP_RBC1131_n_24179 ( .a(FE_OCP_RBN1130_n_24179), .o(FE_OCP_RBN1131_n_24179) );
na02f80 FE_RC_1534_0 ( .a(FE_RN_432_0), .b(FE_RN_433_0), .o(FE_RN_434_0) );
in01f80 FE_OCP_RBC1351_n_19148 ( .a(FE_OCP_RBN1350_n_19148), .o(FE_OCP_RBN1351_n_19148) );
na02f80 g768784 ( .a(n_11956), .b(n_11766), .o(n_11957) );
na02f80 g741692 ( .a(n_38523), .b(n_38217), .o(n_38539) );
na02f80 g758722 ( .a(n_21657), .b(n_20060), .o(n_21792) );
in01f80 newInst_743 ( .a(newNet_742), .o(newNet_743) );
no02f80 g737255 ( .a(n_42905), .b(n_42401), .o(n_42975) );
na02f80 g740236 ( .a(n_39811), .b(n_39859), .o(n_39860) );
no02f80 g744019 ( .a(n_36882), .b(n_36880), .o(n_36881) );
na02f80 g780785 ( .a(n_429), .b(n_373), .o(n_455) );
oa22f80 g758562 ( .a(n_22526), .b(n_21859), .c(n_22525), .d(n_21860), .o(n_22606) );
na02f80 FE_RC_1966_0 ( .a(FE_RN_635_0), .b(n_24323), .o(FE_RN_636_0) );
no02f80 g774299 ( .a(n_6621), .b(n_6620), .o(n_6899) );
no02f80 FE_RC_3842_0 ( .a(FE_RN_1673_0), .b(FE_RN_1674_0), .o(FE_RN_1675_0) );
no02f80 g762206 ( .a(n_18773), .b(n_45002), .o(n_18882) );
na02f80 g747160 ( .a(n_33888), .b(n_33553), .o(n_33953) );
in01f80 g749418 ( .a(n_30601), .o(n_30602) );
na02f80 g752798 ( .a(n_27951), .b(n_27575), .o(n_27993) );
oa22f80 g752591 ( .a(n_27578), .b(n_27544), .c(FE_OCP_RBN3125_n_27578), .d(n_27545), .o(n_27617) );
na02f80 g736925 ( .a(FE_OCP_RBN3699_n_43015), .b(n_43021), .o(n_43054) );
in01f80 FE_RC_3844_0 ( .a(n_23330), .o(FE_RN_1676_0) );
na02f80 g742067 ( .a(n_38007), .b(n_37588), .o(n_38089) );
no02f80 g743993 ( .a(n_36331), .b(n_36294), .o(n_36365) );
in01f80 g759920 ( .a(n_21252), .o(n_21205) );
no02f80 g761255 ( .a(FE_OCP_RBN3825_n_18951), .b(n_18323), .o(n_19013) );
in01f80 newInst_2944 ( .a(newNet_2943), .o(newNet_2944) );
na02f80 FE_RC_3045_0 ( .a(n_35375), .b(FE_RN_1333_0), .o(n_35467) );
oa22f80 FE_RC_1475_0 ( .a(n_24059), .b(n_27785), .c(n_27796), .d(n_27758), .o(n_27843) );
in01f80 g754827 ( .a(n_26007), .o(n_26008) );
in01f80 FE_OCP_RBC1210_n_16814 ( .a(FE_OCP_RBN1207_n_16814), .o(FE_OCP_RBN1210_n_16814) );
in01f80 g753841 ( .a(n_26399), .o(n_26400) );
ao12f80 g773989 ( .a(n_6947), .b(n_6946), .c(n_6945), .o(n_7026) );
in01f80 FE_RC_601_0 ( .a(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .o(FE_RN_189_0) );
na02f80 g745994 ( .a(n_33956), .b(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33981) );
oa12f80 g743055 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .c(delay_add_ln22_unr23_stage9_stallmux_q_9_), .o(n_37008) );
na02f80 FE_RC_2397_0 ( .a(FE_RN_942_0), .b(n_42590), .o(FE_RN_943_0) );
in01f80 g778064 ( .a(n_3038), .o(n_3329) );
no02f80 g773680 ( .a(n_7332), .b(n_7316), .o(n_7317) );
no02f80 g773617 ( .a(n_7347), .b(n_7195), .o(n_7363) );
na02f80 g781022 ( .a(cos_out_2), .b(FE_OFN2_n_43918), .o(n_343) );
na02f80 g744800 ( .a(n_35143), .b(FE_OCPN1434_n_30614), .o(n_35223) );
in01f80 g773275 ( .a(n_7730), .o(n_7802) );
in01f80 g752258 ( .a(n_28669), .o(n_28555) );
na02f80 g773880 ( .a(n_6952), .b(n_5511), .o(n_7048) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_30_ ( .ck(newNet_2359), .d(n_36615), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_30_) );
na02f80 g753143 ( .a(n_27338), .b(n_27382), .o(n_27490) );
no02f80 g754839 ( .a(n_25418), .b(n_25393), .o(n_25454) );
in01f80 g777307 ( .a(n_4612), .o(n_4613) );
no02f80 g770463 ( .a(n_10572), .b(n_10560), .o(n_10561) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_20_ ( .ck(newNet_3621), .d(n_17294), .o(delay_add_ln22_unr11_stage5_stallmux_q_20_) );
oa22f80 FE_RC_716_0 ( .a(n_7399), .b(n_8139), .c(n_7400), .d(n_8138), .o(n_8242) );
in01f80 FE_OCP_RBC3465_n_7886 ( .a(FE_OCP_RBN3459_n_7886), .o(FE_OCP_RBN3465_n_7886) );
in01f80 newInst_2784 ( .a(newNet_2783), .o(newNet_2784) );
ao12f80 g748756 ( .a(n_27246), .b(n_31061), .c(n_30889), .o(n_31063) );
no02f80 g745240 ( .a(n_35968), .b(n_35937), .o(n_35970) );
na02f80 g737955 ( .a(n_42201), .b(n_42047), .o(n_42339) );
in01f80 newInst_1518 ( .a(newNet_1517), .o(newNet_1518) );
na02f80 g779399 ( .a(n_1525), .b(n_1556), .o(n_1662) );
na02f80 FE_RC_673_0 ( .a(FE_RN_213_0), .b(FE_RN_214_0), .o(FE_RN_215_0) );
in01f80 FE_OCP_RBC2988_n_35539 ( .a(FE_OCP_RBN3698_n_35543), .o(FE_OCP_RBN2988_n_35539) );
no02f80 g752507 ( .a(n_28328), .b(n_27955), .o(n_28378) );
in01f80 g776803 ( .a(n_4334), .o(n_4335) );
no02f80 g773078 ( .a(n_7914), .b(n_7913), .o(n_8430) );
no02f80 g757223 ( .a(n_23490), .b(n_23060), .o(n_23549) );
no02f80 g756863 ( .a(n_23750), .b(n_23702), .o(n_23753) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_8_ ( .ck(newNet_1463), .d(n_31856), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_) );
in01f80 g748379 ( .a(n_31793), .o(n_31794) );
oa12f80 g774272 ( .a(n_6414), .b(n_6487), .c(n_6295), .o(n_6493) );
na02f80 g762653 ( .a(n_18017), .b(n_18066), .o(n_18168) );
na02f80 g742402 ( .a(n_37759), .b(n_37738), .o(n_37817) );
no02f80 g761326 ( .a(n_19953), .b(n_19871), .o(n_20741) );
no02f80 g740150 ( .a(FE_OCP_RBN3055_n_39913), .b(n_39869), .o(n_40220) );
in01f80 FE_RC_4244_0 ( .a(n_26467), .o(FE_RN_1866_0) );
in01f80 g774764 ( .a(n_6465), .o(n_6466) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_10_ ( .ck(newNet_2980), .d(n_5569), .o(delay_add_ln22_unr5_stage3_stallmux_q_10_) );
in01f80 FE_OCP_RBC3047_n_6013 ( .a(n_6013), .o(FE_OCP_RBN3047_n_6013) );
na02f80 g780540 ( .a(n_700), .b(n_697), .o(n_727) );
no02f80 g774512 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .o(n_6755) );
in01f80 g748860 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_1_), .o(n_32684) );
ao12f80 g763433 ( .a(n_17366), .b(n_17576), .c(n_17614), .o(n_17615) );
na02f80 g779009 ( .a(n_2077), .b(n_1628), .o(n_2093) );
in01f80 g743447 ( .a(n_36615), .o(n_36585) );
in01f80 g745232 ( .a(n_34573), .o(n_34518) );
oa12f80 g780433 ( .a(n_1110), .b(n_1109), .c(n_1108), .o(n_1140) );
no02f80 g767523 ( .a(n_13224), .b(n_13183), .o(n_13291) );
ao12f80 g750747 ( .a(n_30307), .b(n_30306), .c(n_29850), .o(n_30359) );
in01f80 g758569 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_), .o(n_23403) );
na02f80 g757384 ( .a(n_23036), .b(n_23035), .o(n_23037) );
in01f80 g754064 ( .a(n_26198), .o(n_26240) );
na02f80 g778516 ( .a(n_2484), .b(n_2483), .o(n_2582) );
in01f80 g736840 ( .a(n_43040), .o(n_43041) );
no02f80 g736544 ( .a(n_43651), .b(n_43285), .o(n_43686) );
no02f80 g762212 ( .a(n_18734), .b(FE_OFN750_n_45003), .o(n_18771) );
ao22s80 g776897 ( .a(n_47014), .b(n_3788), .c(FE_OCP_RBN3589_n_47014), .d(n_3912), .o(n_4030) );
na02f80 g760241 ( .a(FE_OCPN1261_n_20242), .b(n_20430), .o(n_20489) );
in01f80 g745614 ( .a(n_34486), .o(n_34535) );
ao22s80 g747288 ( .a(n_32616), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .c(n_32638), .d(n_31260), .o(n_32693) );
na02f80 g754097 ( .a(n_26079), .b(FE_OCPN1440_n_23339), .o(n_26149) );
in01f80 g745788 ( .a(n_34334), .o(n_34335) );
in01f80 g747545 ( .a(n_33672), .o(n_33705) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_9_ ( .ck(newNet_2797), .d(n_10705), .o(delay_add_ln22_unr8_stage4_stallmux_q_9_) );
in01f80 g751488 ( .a(n_28885), .o(n_28886) );
in01f80 newInst_436 ( .a(newNet_435), .o(newNet_436) );
in01f80 g761603 ( .a(n_19787), .o(n_19980) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_5_ ( .ck(newNet_2243), .d(n_40410), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_5_) );
in01f80 FE_OCP_RBC3372_n_6745 ( .a(FE_OCP_RBN2127_n_6745), .o(FE_OCP_RBN3372_n_6745) );
no02f80 g743767 ( .a(n_37284), .b(n_36793), .o(n_37285) );
in01f80 g751398 ( .a(n_29311), .o(n_29312) );
in01f80 g748560 ( .a(n_31449), .o(n_31476) );
in01f80 newInst_2076 ( .a(newNet_65), .o(newNet_2076) );
in01f80 g772395 ( .a(n_8619), .o(n_8620) );
oa12f80 g740852 ( .a(n_39223), .b(n_39222), .c(n_39221), .o(n_39832) );
oa22f80 g737650 ( .a(n_42392), .b(n_41983), .c(FE_OCPN888_n_42367), .d(n_41993), .o(n_42728) );
in01f80 g770768 ( .a(n_10355), .o(n_10254) );
no02f80 g761861 ( .a(n_18595), .b(n_18594), .o(n_18596) );
ao12f80 g778458 ( .a(n_2407), .b(n_2406), .c(FE_OFN812_n_2405), .o(n_2488) );
in01f80 g768735 ( .a(n_12148), .o(n_12149) );
no02f80 FE_RC_1944_0 ( .a(FE_RN_619_0), .b(FE_RN_620_0), .o(FE_RN_621_0) );
na02f80 g756590 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_28_), .o(n_23817) );
in01f80 FE_OCP_RBC2679_n_14768 ( .a(n_14768), .o(FE_OCP_RBN2679_n_14768) );
in01f80 g737285 ( .a(n_42898), .o(n_42899) );
na02f80 g749841 ( .a(FE_OCP_RBN3009_n_31117), .b(n_30416), .o(n_31221) );
no02f80 g766032 ( .a(n_14611), .b(n_14610), .o(n_14693) );
na02f80 g774337 ( .a(n_6697), .b(n_6737), .o(n_7297) );
in01f80 g747934 ( .a(n_33372), .o(n_33392) );
in01f80 g775837 ( .a(n_5501), .o(n_5502) );
no02f80 g755145 ( .a(n_25070), .b(n_25116), .o(n_25244) );
in01f80 g758828 ( .a(n_21804), .o(n_21805) );
na02f80 g736730 ( .a(n_43213), .b(n_43226), .o(n_43692) );
in01f80 g755900 ( .a(n_24311), .o(n_24312) );
oa12f80 g757928 ( .a(n_22812), .b(n_22731), .c(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(n_22887) );
in01f80 g768668 ( .a(n_12217), .o(n_12190) );
in01f80 g764346 ( .a(n_16454), .o(n_16455) );
in01f80 g772528 ( .a(n_8590), .o(n_8617) );
na02f80 g736888 ( .a(n_43493), .b(n_43529), .o(n_43593) );
ao12f80 g779022 ( .a(n_2055), .b(n_2054), .c(n_2053), .o(n_2596) );
no02f80 FE_RC_2431_0 ( .a(FE_RN_966_0), .b(n_6826), .o(FE_RN_967_0) );
in01f80 FE_OCP_RBC2604_n_39126 ( .a(n_39126), .o(FE_OCP_RBN2604_n_39126) );
in01f80 g749002 ( .a(n_31101), .o(n_31102) );
ao12f80 g757220 ( .a(n_23124), .b(n_23191), .c(n_23187), .o(n_23235) );
no02f80 g761491 ( .a(n_19647), .b(n_19790), .o(n_19822) );
in01f80 FE_OCP_RBC2287_n_2268 ( .a(n_2268), .o(FE_OCP_RBN2287_n_2268) );
no02f80 g766791 ( .a(n_13661), .b(FE_OCP_RBN2244_n_13017), .o(n_13690) );
in01f80 newInst_3000 ( .a(newNet_2999), .o(newNet_3000) );
no02f80 g766206 ( .a(n_14447), .b(n_14369), .o(n_14483) );
na02f80 g753493 ( .a(FE_OCP_RBN2983_n_26767), .b(n_26762), .o(n_26763) );
no02f80 g774480 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .o(n_6687) );
in01f80 g748301 ( .a(n_31608), .o(n_31609) );
in01f80 g764306 ( .a(n_16374), .o(n_16375) );
in01f80 newInst_358 ( .a(newNet_324), .o(newNet_358) );
in01f80 g782638 ( .a(n_44032), .o(n_44033) );
ao12f80 g768761 ( .a(n_12035), .b(n_12034), .c(n_12033), .o(n_12789) );
in01f80 g741621 ( .a(n_38626), .o(n_38639) );
oa22f80 g747446 ( .a(n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_0_), .c(FE_OCP_RBN3332_n_44962), .d(n_32387), .o(n_32525) );
in01f80 newInst_2788 ( .a(newNet_2660), .o(newNet_2788) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_23_ ( .ck(newNet_1606), .d(n_27479), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_) );
in01f80 FE_OCPC1494_n_23398 ( .a(FE_OCPN1493_n_23398), .o(FE_OCPN1494_n_23398) );
in01f80 newInst_2408 ( .a(newNet_2407), .o(newNet_2408) );
na02f80 g737539 ( .a(n_42290), .b(n_42254), .o(n_42337) );
na02f80 g766122 ( .a(n_14545), .b(n_44850), .o(n_14580) );
in01f80 g754424 ( .a(n_25757), .o(n_25777) );
in01f80 fopt784701 ( .a(n_47180), .o(n_47181) );
no02f80 g738550 ( .a(n_41689), .b(n_41537), .o(n_41742) );
in01f80 FE_RC_1720_0 ( .a(n_28219), .o(FE_RN_475_0) );
na02f80 g741498 ( .a(n_38739), .b(n_38738), .o(n_38744) );
no02f80 g756566 ( .a(n_23563), .b(n_22669), .o(n_23664) );
na02f80 g746492 ( .a(n_34529), .b(n_34525), .o(n_34552) );
in01f80 g761580 ( .a(n_20252), .o(n_22961) );
in01f80 newInst_2201 ( .a(newNet_660), .o(newNet_2201) );
ao12f80 g761307 ( .a(n_19029), .b(n_19028), .c(n_19027), .o(n_19098) );
oa12f80 g784670 ( .a(n_5468), .b(n_5452), .c(n_4908), .o(n_47000) );
ao12f80 g761219 ( .a(n_19984), .b(n_20036), .c(n_19980), .o(n_21140) );
in01f80 newInst_2819 ( .a(newNet_2818), .o(newNet_2819) );
in01f80 FE_RC_3649_0 ( .a(n_21955), .o(FE_RN_1601_0) );
in01f80 g766430 ( .a(n_14268), .o(n_14269) );
oa12f80 g772548 ( .a(n_8558), .b(n_8557), .c(n_8556), .o(n_9367) );
in01f80 g780188 ( .a(n_1090), .o(n_1091) );
no02f80 g762088 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_28_), .o(n_18541) );
no02f80 g764791 ( .a(n_15510), .b(n_15274), .o(n_15559) );
in01f80 g753913 ( .a(n_27210), .o(n_26323) );
na02f80 g758840 ( .a(n_21476), .b(n_45026), .o(n_21556) );
oa12f80 g772286 ( .a(n_8723), .b(n_8722), .c(n_8721), .o(n_9913) );
no02f80 g760911 ( .a(n_19380), .b(n_17881), .o(n_19469) );
in01f80 g761837 ( .a(n_18322), .o(n_18379) );
oa12f80 g766197 ( .a(n_14998), .b(n_14677), .c(n_14676), .o(n_14732) );
no02f80 g744982 ( .a(n_34827), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34882) );
na02f80 g754728 ( .a(n_26541), .b(n_26643), .o(n_26601) );
no02f80 g740803 ( .a(n_39293), .b(n_39142), .o(n_39294) );
no02f80 g743554 ( .a(n_36472), .b(n_36066), .o(n_36473) );
na02f80 g749420 ( .a(n_30513), .b(n_30297), .o(n_30582) );
in01f80 newInst_2825 ( .a(newNet_2824), .o(newNet_2825) );
no02f80 g760788 ( .a(n_19563), .b(FE_OCP_DRV_N1562_n_19562), .o(n_19594) );
na02f80 g767928 ( .a(n_12651), .b(n_12455), .o(n_12686) );
oa22f80 FE_RC_3969_0 ( .a(n_24207), .b(n_25228), .c(n_24125), .d(n_24269), .o(n_24291) );
na02f80 g751564 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_27_), .o(n_28720) );
na02f80 g752750 ( .a(n_27512), .b(n_27352), .o(n_27549) );
no02f80 g761680 ( .a(n_18794), .b(n_18750), .o(n_18948) );
in01f80 g764221 ( .a(n_16601), .o(n_16578) );
ao12f80 g756882 ( .a(n_23743), .b(n_23834), .c(n_23897), .o(n_23958) );
in01f80 g775932 ( .a(n_5534), .o(n_5374) );
na02f80 g739888 ( .a(n_40298), .b(n_39975), .o(n_40345) );
no02f80 g750128 ( .a(FE_OCP_RBN2573_n_29922), .b(n_30310), .o(n_30343) );
no02f80 g771007 ( .a(n_9763), .b(n_9663), .o(n_9847) );
in01f80 g771724 ( .a(n_8983), .o(n_8992) );
na02f80 g779754 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_1731) );
in01f80 FE_OCP_DRV_C1603_n_19961 ( .a(n_19961), .o(FE_OCP_DRV_N1603_n_19961) );
no02f80 FE_RC_3066_0 ( .a(n_20654), .b(FE_RN_1347_0), .o(FE_RN_1348_0) );
oa22f80 g764355 ( .a(n_16653), .b(n_16060), .c(n_16673), .d(n_16061), .o(n_16767) );
oa12f80 g751410 ( .a(n_29256), .b(n_29255), .c(n_29254), .o(n_29838) );
ao12f80 g750591 ( .a(n_30434), .b(n_30440), .c(n_30433), .o(n_31172) );
in01f80 g749321 ( .a(n_30865), .o(n_30866) );
no02f80 g777971 ( .a(n_3154), .b(n_3178), .o(n_3179) );
oa12f80 g753692 ( .a(n_26325), .b(n_26506), .c(n_26403), .o(n_26599) );
na02f80 g767798 ( .a(n_12823), .b(n_12215), .o(n_12956) );
na02f80 g744252 ( .a(FE_OCPN1510_n_44174), .b(n_35554), .o(n_36183) );
no02f80 g757854 ( .a(n_22422), .b(n_22145), .o(n_22475) );
no02f80 g757053 ( .a(n_23700), .b(n_23860), .o(n_24007) );
oa12f80 g757729 ( .a(n_22298), .b(n_22556), .c(n_22333), .o(n_22598) );
in01f80 g776078 ( .a(n_4998), .o(n_5018) );
na03f80 g751754 ( .a(n_28063), .b(n_28271), .c(n_28270), .o(n_28295) );
ao22s80 g757283 ( .a(n_23417), .b(n_23201), .c(n_23416), .d(n_23202), .o(n_23985) );
na02f80 g750703 ( .a(n_29234), .b(n_28826), .o(n_29300) );
in01f80 g745012 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_6_), .o(n_36358) );
na02f80 g777093 ( .a(n_3751), .b(n_3734), .o(n_3879) );
na02f80 FE_RC_2937_0 ( .a(n_29417), .b(n_29697), .o(FE_RN_1281_0) );
na02f80 g749958 ( .a(n_30021), .b(n_29985), .o(n_30376) );
na02f80 g752689 ( .a(n_28202), .b(n_28156), .o(n_28157) );
in01f80 g751331 ( .a(n_28656), .o(n_28657) );
na02f80 g781031 ( .a(cos_out_17), .b(FE_OFN2_n_43918), .o(n_329) );
in01f80 newInst_951 ( .a(newNet_950), .o(newNet_951) );
no02f80 g764500 ( .a(n_16542), .b(n_15878), .o(n_16615) );
in01f80 FE_OCPC903_n_44581 ( .a(FE_OCPN902_n_44581), .o(FE_OCPN903_n_44581) );
no02f80 g745881 ( .a(n_34015), .b(n_34017), .o(n_34016) );
na02f80 g778919 ( .a(n_2284), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_), .o(n_2358) );
in01f80 g757885 ( .a(n_22237), .o(n_22316) );
no02f80 g766216 ( .a(n_14468), .b(FE_OCP_RBN2249_n_13017), .o(n_14469) );
in01f80 g773086 ( .a(n_8086), .o(n_8087) );
in01f80 newInst_3368 ( .a(newNet_3367), .o(newNet_3368) );
no02f80 FE_RC_2359_0 ( .a(FE_RN_909_0), .b(FE_RN_910_0), .o(FE_RN_911_0) );
na02f80 g741213 ( .a(n_38818), .b(n_38817), .o(n_38894) );
oa12f80 g758596 ( .a(n_21883), .b(n_22489), .c(n_21832), .o(n_22549) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_16_ ( .ck(newNet_357), .d(n_1350), .o(delay_xor_ln22_unr3_stage2_stallmux_q_16_) );
oa22f80 FE_RC_852_0 ( .a(FE_OCP_RBN3546_n_44575), .b(n_9182), .c(n_44563), .d(FE_OCP_RBN2719_n_9182), .o(n_9400) );
in01f80 g761464 ( .a(n_19905), .o(n_19872) );
ao12f80 g751919 ( .a(n_29308), .b(n_28919), .c(n_28689), .o(n_29741) );
na02f80 g754105 ( .a(n_26118), .b(n_23353), .o(n_26204) );
in01f80 g737495 ( .a(n_42597), .o(n_42598) );
na02f80 g763406 ( .a(FE_OCP_RBN3724_n_16975), .b(n_16003), .o(n_17178) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_2_ ( .ck(newNet_2073), .d(n_4590), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_2_) );
no02f80 g739225 ( .a(n_40674), .b(delay_add_ln22_unr27_stage10_stallmux_q_11_), .o(n_40680) );
ao22s80 FE_RC_4130_0 ( .a(n_32473), .b(n_32625), .c(n_32472), .d(n_32596), .o(n_32667) );
in01f80 g744246 ( .a(n_35531), .o(n_36243) );
in01f80 g746619 ( .a(n_34638), .o(n_34608) );
na02f80 g770744 ( .a(n_9819), .b(FE_OCP_RBN2478_n_8599), .o(n_9974) );
in01f80 g737449 ( .a(n_42716), .o(n_42717) );
na02f80 g739301 ( .a(n_40720), .b(n_40545), .o(n_40764) );
na02f80 g759131 ( .a(n_21909), .b(n_21376), .o(n_21977) );
no02f80 g778036 ( .a(n_3036), .b(n_2994), .o(n_3098) );
in01f80 FE_OCP_RBC2343_FE_OCPN870_n_2737 ( .a(FE_OCP_RBN2342_FE_OCPN870_n_2737), .o(FE_OCP_RBN2343_FE_OCPN870_n_2737) );
in01f80 g760591 ( .a(n_19818), .o(n_19819) );
na02f80 g736939 ( .a(n_43242), .b(n_43147), .o(n_43460) );
oa12f80 g760442 ( .a(n_20044), .b(n_20078), .c(n_20077), .o(n_20145) );
no02f80 g757845 ( .a(n_22446), .b(n_22448), .o(n_22476) );
in01f80 FE_OCPC1044_n_20307 ( .a(FE_OCPN1043_n_20307), .o(FE_OCPN1044_n_20307) );
na02f80 g747376 ( .a(FE_OCP_RBN3332_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_2_), .o(n_32437) );
no02f80 g736613 ( .a(n_43481), .b(n_43364), .o(n_43626) );
na02f80 g772997 ( .a(n_7718), .b(n_8389), .o(n_7746) );
in01f80 g752690 ( .a(n_28216), .o(n_28261) );
in01f80 fopt783562 ( .a(n_45180), .o(n_45181) );
na02f80 g740248 ( .a(n_39851), .b(n_39889), .o(n_39890) );
ao12f80 g737640 ( .a(n_42527), .b(n_42392), .c(n_42112), .o(n_42825) );
na02f80 g770182 ( .a(n_10670), .b(n_10735), .o(n_10757) );
in01f80 newInst_2829 ( .a(newNet_2828), .o(newNet_2829) );
na02f80 FE_RC_1079_0 ( .a(FE_RN_318_0), .b(FE_RN_319_0), .o(FE_RN_320_0) );
in01f80 g757682 ( .a(n_22818), .o(n_22791) );
no02f80 g778693 ( .a(n_2289), .b(FE_OCPN3759_n_2346), .o(n_2282) );
oa22f80 FE_RC_886_0 ( .a(FE_OFN802_n_46285), .b(n_12114), .c(FE_OFN771_n_46337), .d(n_12037), .o(n_46357) );
no02f80 g758187 ( .a(n_44268), .b(FE_OCP_DRV_N3162_n_21419), .o(n_22194) );
in01f80 g761164 ( .a(n_19112), .o(n_19140) );
na02f80 g778102 ( .a(n_2951), .b(n_3006), .o(n_3007) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_27_ ( .ck(newNet_2543), .d(n_27785), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_) );
na02f80 g769650 ( .a(n_11308), .b(FE_OCP_RBN2821_n_10023), .o(n_11375) );
na02f80 g739210 ( .a(n_40788), .b(n_40787), .o(n_40789) );
na02f80 FE_RC_3635_0 ( .a(FE_RN_1593_0), .b(n_31518), .o(n_31549) );
in01f80 g775666 ( .a(n_5442), .o(n_5443) );
in01f80 g752240 ( .a(n_28005), .o(n_28006) );
in01f80 g769720 ( .a(n_11242), .o(n_11243) );
na02f80 g756599 ( .a(n_23631), .b(n_23578), .o(n_23894) );
no02f80 g769744 ( .a(n_11148), .b(n_11121), .o(n_11223) );
no02f80 g776267 ( .a(n_4733), .b(n_4713), .o(n_4887) );
in01f80 FE_OCP_RBC3087_n_36535 ( .a(n_36535), .o(FE_OCP_RBN3087_n_36535) );
na02f80 g740048 ( .a(n_39918), .b(n_39953), .o(n_39954) );
in01f80 g749371 ( .a(n_32035), .o(n_32063) );
no02f80 g740999 ( .a(n_39133), .b(n_39134), .o(n_39191) );
in01f80 newInst_3659 ( .a(newNet_2198), .o(newNet_3659) );
na02f80 g743224 ( .a(n_36801), .b(n_36756), .o(n_36846) );
in01f80 g745861 ( .a(n_34135), .o(n_34136) );
na02f80 g766914 ( .a(n_13582), .b(n_13589), .o(n_13615) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_23_ ( .ck(newNet_3044), .d(n_1205), .o(delay_add_ln22_unr2_stage2_stallmux_q_23_) );
no02f80 g768832 ( .a(n_11942), .b(n_9949), .o(n_12097) );
no04s80 g747295 ( .a(n_32599), .b(n_32595), .c(n_32522), .d(n_32602), .o(n_32641) );
no02f80 g751371 ( .a(n_28536), .b(n_28514), .o(n_28515) );
in01f80 g759171 ( .a(n_21192), .o(n_21126) );
oa22f80 g784364 ( .a(FE_OFN775_n_46137), .b(n_5708), .c(FE_OFN805_n_46196), .d(n_5724), .o(n_46170) );
na02f80 g779232 ( .a(n_1865), .b(n_946), .o(n_1953) );
in01f80 FE_RC_1277_0 ( .a(n_2914), .o(FE_RN_376_0) );
no02f80 g745046 ( .a(n_34860), .b(n_34826), .o(n_34923) );
no02f80 g772745 ( .a(n_8128), .b(n_8071), .o(n_8179) );
no02f80 g745152 ( .a(n_34576), .b(n_34575), .o(n_34577) );
no02f80 g773797 ( .a(n_7188), .b(n_7006), .o(n_7218) );
no02f80 FE_RC_2040_0 ( .a(FE_RN_682_0), .b(n_27120), .o(n_27146) );
oa12f80 g747291 ( .a(n_33631), .b(n_33630), .c(n_33629), .o(n_34645) );
in01f80 g770427 ( .a(n_10634), .o(n_10635) );
oa22f80 FE_RC_417_0 ( .a(n_13010), .b(n_13144), .c(n_13146), .d(FE_OCP_RBN2221_n_13010), .o(n_13225) );
in01f80 newInst_524 ( .a(newNet_523), .o(newNet_524) );
na03f80 FE_RC_2519_0 ( .a(FE_RN_1025_0), .b(n_37366), .c(n_37353), .o(n_37369) );
in01f80 newInst_1500 ( .a(newNet_1499), .o(newNet_1500) );
in01f80 FE_OCP_RBC2486_n_3498 ( .a(n_3498), .o(FE_OCP_RBN2486_n_3498) );
na02f80 g754846 ( .a(n_25275), .b(n_24332), .o(n_25303) );
in01f80 FE_OCP_RBC2312_n_41420 ( .a(n_41420), .o(FE_OCP_RBN2312_n_41420) );
in01f80 FE_OCP_RBC2482_n_14326 ( .a(n_14326), .o(FE_OCP_RBN2482_n_14326) );
na02f80 g737602 ( .a(n_42464), .b(n_42448), .o(n_42489) );
na02f80 g759723 ( .a(n_20612), .b(n_20587), .o(n_20678) );
oa12f80 g755636 ( .a(n_25188), .b(n_25286), .c(n_24979), .o(n_25345) );
na02f80 g772960 ( .a(n_7813), .b(n_7509), .o(n_7825) );
in01f80 g739848 ( .a(n_40300), .o(n_40349) );
no02f80 g742489 ( .a(n_37597), .b(n_37709), .o(n_37627) );
in01f80 g755973 ( .a(FE_OFN788_n_25834), .o(n_25738) );
in01f80 g769216 ( .a(n_11451), .o(n_11520) );
oa12f80 g756350 ( .a(n_23517), .b(n_23827), .c(n_23556), .o(n_23930) );
no02f80 g757506 ( .a(n_22799), .b(n_22821), .o(n_22930) );
no02f80 g747801 ( .a(n_33372), .b(n_32901), .o(n_33421) );
in01f80 g739707 ( .a(n_40519), .o(n_40520) );
no02f80 g765267 ( .a(n_15576), .b(n_15575), .o(n_15577) );
in01f80 g775650 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_9_), .o(n_5511) );
na02f80 g774750 ( .a(n_6369), .b(n_6269), .o(n_6417) );
in01f80 newInst_771 ( .a(newNet_770), .o(newNet_771) );
in01f80 FE_OCP_RBC2303_n_7817 ( .a(FE_OCP_RBN2302_n_7817), .o(FE_OCP_RBN2303_n_7817) );
no02f80 g745528 ( .a(n_34764), .b(n_34321), .o(n_34819) );
na02f80 g751989 ( .a(n_28781), .b(n_28835), .o(n_28991) );
in01f80 g751484 ( .a(n_28826), .o(n_28827) );
in01f80 FE_OCPC1786_n_30134 ( .a(FE_OCPN1785_n_30134), .o(FE_OCPN1786_n_30134) );
ao22s80 FE_RC_830_0 ( .a(n_22089), .b(FE_OCP_RBN2422_n_24501), .c(n_22280), .d(n_24501), .o(n_24618) );
na02f80 g745445 ( .a(n_35926), .b(n_35525), .o(n_35526) );
na02f80 g754721 ( .a(n_26541), .b(n_26509), .o(n_26710) );
na02f80 g746027 ( .a(n_35191), .b(n_34669), .o(n_35243) );
na02f80 g767056 ( .a(FE_OCP_RBN2503_n_13896), .b(n_14107), .o(n_14212) );
no03m80 FE_RC_76_0 ( .a(n_17339), .b(n_17436), .c(n_17442), .o(n_17579) );
no02f80 g755261 ( .a(n_24986), .b(n_24819), .o(n_25015) );
in01f80 g776970 ( .a(n_3849), .o(n_3897) );
no02f80 g769686 ( .a(n_11256), .b(n_44511), .o(n_11257) );
in01f80 g741079 ( .a(n_39502), .o(n_39503) );
no02f80 g750792 ( .a(n_29258), .b(n_29096), .o(n_29316) );
in01f80 g760306 ( .a(n_20285), .o(n_20243) );
ao22s80 FE_RC_1345_0 ( .a(n_43828), .b(n_43397), .c(n_43396), .d(n_43827), .o(n_43862) );
na02f80 g774296 ( .a(FE_OCP_RBN3250_delay_xor_ln22_unr6_stage3_stallmux_q_0_), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6546) );
no02f80 g756744 ( .a(n_23426), .b(n_23114), .o(n_23482) );
in01f80 FE_OCP_RBC3602_n_3913 ( .a(n_3913), .o(FE_OCP_RBN3602_n_3913) );
na02f80 g759563 ( .a(n_20447), .b(n_20341), .o(n_20595) );
oa12f80 g759584 ( .a(n_21882), .b(n_21881), .c(n_21880), .o(n_21930) );
na02f80 g772666 ( .a(n_45828), .b(n_8346), .o(n_8316) );
in01f80 newInst_3413 ( .a(newNet_501), .o(newNet_3413) );
in01f80 g747199 ( .a(n_34614), .o(n_34579) );
in01f80 newInst_3594 ( .a(newNet_3593), .o(newNet_3594) );
na02f80 g779290 ( .a(n_1742), .b(n_1741), .o(n_1743) );
na02f80 g751575 ( .a(n_28447), .b(n_27475), .o(n_28491) );
na02f80 g764869 ( .a(n_45502), .b(n_14420), .o(n_15556) );
na02f80 g739243 ( .a(n_40933), .b(n_40903), .o(n_40954) );
na02f80 g763677 ( .a(n_17365), .b(n_17428), .o(n_17429) );
in01f80 g749390 ( .a(n_46959), .o(n_30646) );
no02f80 g745447 ( .a(n_35540), .b(n_34965), .o(n_35541) );
in01f80 g757577 ( .a(n_22901), .o(n_22861) );
oa12f80 g746360 ( .a(n_33490), .b(n_33489), .c(n_33488), .o(n_33541) );
in01f80 FE_OCP_RBC3459_n_7886 ( .a(n_7886), .o(FE_OCP_RBN3459_n_7886) );
no02f80 g766324 ( .a(n_14496), .b(FE_OCP_RBN2509_n_13896), .o(n_14568) );
no02f80 g769252 ( .a(FE_OCP_RBN3094_n_11475), .b(n_10676), .o(n_11623) );
no02f80 g752777 ( .a(n_27356), .b(n_27437), .o(n_27436) );
no02f80 g777087 ( .a(n_3803), .b(n_3698), .o(n_3852) );
no02f80 g766885 ( .a(n_13846), .b(n_14340), .o(n_14454) );
no02f80 g777289 ( .a(n_3639), .b(n_3118), .o(n_3567) );
in01f80 g774833 ( .a(n_6345), .o(n_6346) );
no02f80 g756481 ( .a(n_23884), .b(n_23853), .o(n_23923) );
in01f80 g760861 ( .a(n_19393), .o(n_19479) );
in01f80 FE_OCPC939_n_7712 ( .a(n_7712), .o(FE_OCPN939_n_7712) );
in01f80 g740347 ( .a(n_40304), .o(n_40305) );
no02f80 g767638 ( .a(n_13392), .b(n_13369), .o(n_13442) );
in01f80 g780351 ( .a(n_972), .o(n_1017) );
in01f80 fopt783139 ( .a(n_1282), .o(n_44636) );
in01f80 FE_RC_3669_0 ( .a(n_21289), .o(FE_RN_1612_0) );
oa12f80 g759399 ( .a(n_20459), .b(n_20973), .c(FE_OCP_RBN2739_n_20432), .o(n_21002) );
in01f80 g737056 ( .a(n_43126), .o(n_43168) );
in01f80 FE_RC_2901_0 ( .a(n_19497), .o(FE_RN_1258_0) );
no02f80 g750109 ( .a(n_29857), .b(n_29167), .o(n_30195) );
na02f80 g771658 ( .a(n_8969), .b(n_8971), .o(n_8972) );
in01f80 g757169 ( .a(n_23646), .o(n_23671) );
na02f80 g756508 ( .a(n_23608), .b(n_23583), .o(n_23680) );
in01f80 g761137 ( .a(n_19173), .o(n_19174) );
no02f80 g771796 ( .a(n_9049), .b(n_8988), .o(n_9240) );
in01f80 g739015 ( .a(n_41198), .o(n_41142) );
no02f80 g758010 ( .a(n_22262), .b(n_22301), .o(n_22387) );
oa22f80 g747756 ( .a(FE_OCP_RBN3099_n_32001), .b(n_31912), .c(n_32001), .d(n_31913), .o(n_32085) );
in01f80 g762893 ( .a(n_17728), .o(n_17682) );
ao22s80 g736480 ( .a(n_43735), .b(n_43344), .c(n_43722), .d(n_43345), .o(n_43761) );
oa22f80 g764277 ( .a(n_16675), .b(n_16303), .c(n_16676), .d(n_16302), .o(n_16744) );
in01f80 g761870 ( .a(n_18513), .o(n_18514) );
in01f80 FE_OCP_RBC2469_n_19806 ( .a(n_19806), .o(FE_OCP_RBN2469_n_19806) );
in01f80 g741539 ( .a(n_38726), .o(n_38727) );
in01f80 g762299 ( .a(FE_OCPUNCON1804_n_18111), .o(n_18112) );
in01f80 g764302 ( .a(n_16376), .o(n_16402) );
no02f80 g760153 ( .a(n_20456), .b(n_19654), .o(n_20778) );
na02f80 g765098 ( .a(n_15527), .b(n_15526), .o(n_15528) );
no02f80 g767035 ( .a(FE_OCP_RBN2459_n_13765), .b(n_13936), .o(n_13974) );
ao12f80 g772454 ( .a(n_45212), .b(n_8386), .c(n_8406), .o(n_8461) );
in01f80 g778454 ( .a(n_2685), .o(n_2686) );
in01f80 g775377 ( .a(n_5717), .o(n_5718) );
no02f80 g778334 ( .a(n_2585), .b(n_2473), .o(n_2586) );
na02f80 g749153 ( .a(n_30774), .b(n_30749), .o(n_30888) );
in01f80 FE_RC_2668_0 ( .a(n_4953), .o(FE_RN_1115_0) );
na02f80 g762418 ( .a(n_45118), .b(n_18521), .o(n_18568) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_9_ ( .ck(newNet_2891), .d(n_5483), .o(delay_add_ln22_unr5_stage3_stallmux_q_9_) );
no02f80 g747989 ( .a(n_33043), .b(n_33042), .o(n_33044) );
no02f80 g748178 ( .a(n_31992), .b(n_32049), .o(n_32128) );
in01f80 FE_OCP_RBC2696_n_14814 ( .a(FE_OCP_RBN2695_n_14814), .o(FE_OCP_RBN2696_n_14814) );
na02f80 g744654 ( .a(n_35345), .b(n_35310), .o(n_35311) );
in01f80 g756294 ( .a(n_24070), .o(n_24098) );
in01f80 newInst_2039 ( .a(newNet_295), .o(newNet_2039) );
no02f80 g744519 ( .a(n_35364), .b(n_35231), .o(n_35404) );
na02f80 g770456 ( .a(n_10473), .b(n_10503), .o(n_10562) );
na02f80 g780762 ( .a(n_565), .b(n_564), .o(n_566) );
in01f80 FE_OCP_RBC1323_n_29056 ( .a(n_29056), .o(FE_OCP_RBN1323_n_29056) );
na02f80 g760657 ( .a(n_19752), .b(FE_OCP_DRV_N1568_n_19751), .o(n_19775) );
no02f80 g763301 ( .a(n_17388), .b(n_16996), .o(n_17389) );
oa12f80 g779411 ( .a(n_1407), .b(n_1515), .c(n_1456), .o(n_1551) );
ao22s80 FE_RC_585_0 ( .a(n_23439), .b(n_23167), .c(n_23453), .d(n_23168), .o(n_23539) );
in01f80 g738129 ( .a(FE_OCP_RBN2443_n_42051), .o(n_42069) );
in01f80 g750065 ( .a(n_30077), .o(n_30171) );
no02f80 g746911 ( .a(n_33034), .b(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(n_33159) );
ao12f80 g762657 ( .a(n_17851), .b(FE_OCP_RBN2142_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .o(n_17897) );
na02f80 g745265 ( .a(n_35851), .b(n_35849), .o(n_35940) );
na02f80 g751912 ( .a(n_28881), .b(n_28904), .o(n_29225) );
oa22f80 FE_RC_1585_0 ( .a(n_17336), .b(n_17812), .c(n_16339), .d(n_17809), .o(n_17879) );
in01f80 g764476 ( .a(n_16231), .o(n_16190) );
na02f80 g746010 ( .a(n_33881), .b(n_33880), .o(n_33926) );
in01f80 g766682 ( .a(n_13757), .o(n_13758) );
na02f80 g770419 ( .a(n_10542), .b(n_44463), .o(n_10444) );
na02f80 g736884 ( .a(n_43452), .b(n_43497), .o(n_43597) );
oa22f80 g763625 ( .a(n_46976), .b(FE_OFN767_n_15670), .c(n_16774), .d(n_16339), .o(n_16863) );
no02f80 g776175 ( .a(n_4894), .b(n_4321), .o(n_4944) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_22_ ( .ck(newNet_2941), .d(n_46994), .o(delay_add_ln22_unr5_stage3_stallmux_q_22_) );
no02f80 g780624 ( .a(n_679), .b(n_678), .o(n_684) );
oa12f80 g736349 ( .a(n_291), .b(n_43847), .c(FE_OFN1_n_43918), .o(n_43884) );
na02f80 g745301 ( .a(n_36081), .b(n_36171), .o(n_36219) );
no02f80 g765348 ( .a(n_15127), .b(n_47261), .o(n_15192) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_19_ ( .ck(newNet_1015), .d(n_17878), .o(delay_xor_ln21_unr12_stage5_stallmux_q_19_) );
in01f80 g764483 ( .a(n_16123), .o(n_16124) );
na02f80 g764723 ( .a(n_15850), .b(n_15897), .o(n_16071) );
no02f80 g752198 ( .a(n_44825), .b(n_28615), .o(n_28667) );
na02f80 g757392 ( .a(n_23034), .b(n_44071), .o(n_23160) );
na02f80 g781056 ( .a(sin_out_15), .b(FE_OFN3_n_43918), .o(n_340) );
na02f80 g772966 ( .a(n_7747), .b(n_7026), .o(n_7844) );
in01f80 g751073 ( .a(n_30412), .o(n_30413) );
in01f80 g754028 ( .a(n_26976), .o(n_26977) );
na02f80 g756775 ( .a(n_23411), .b(n_23145), .o(n_23412) );
oa22f80 g754000 ( .a(n_26974), .b(n_26903), .c(n_26949), .d(n_26904), .o(n_27016) );
no02f80 g768127 ( .a(n_12620), .b(n_12619), .o(n_12647) );
ao22s80 g771736 ( .a(n_9035), .b(FE_OCP_RBN3547_n_44575), .c(n_9064), .d(FE_OCP_RBN2606_FE_OCPN899_n_44593), .o(n_9332) );
no02f80 g761040 ( .a(n_19213), .b(n_19114), .o(n_19214) );
in01f80 g776515 ( .a(n_4054), .o(n_4103) );
in01f80 FE_OCP_RBC2517_n_8762 ( .a(n_8762), .o(FE_OCP_RBN2517_n_8762) );
no03m80 FE_RC_2224_0 ( .a(FE_RN_806_0), .b(n_32936), .c(n_33273), .o(FE_RN_807_0) );
no02f80 g748707 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_30_), .o(n_32561) );
in01f80 g764419 ( .a(n_16200), .o(n_16201) );
no02f80 g771836 ( .a(n_9602), .b(n_9695), .o(n_10237) );
ao12f80 g755918 ( .a(n_25340), .b(n_25188), .c(n_25285), .o(n_25739) );
in01f80 g758706 ( .a(n_22396), .o(n_22428) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_23_ ( .ck(newNet_3137), .d(n_40530), .o(delay_add_ln22_unr27_stage10_stallmux_q_23_) );
in01f80 newInst_2939 ( .a(newNet_2938), .o(newNet_2939) );
in01f80 g770683 ( .a(n_9982), .o(n_9983) );
in01f80 FE_RC_2944_0 ( .a(FE_RN_1285_0), .o(n_15494) );
ao12f80 g768099 ( .a(n_12214), .b(n_12663), .c(n_12119), .o(n_12707) );
in01f80 g778511 ( .a(n_2475), .o(n_2410) );
oa22f80 g779863 ( .a(n_44652), .b(n_1211), .c(n_44623), .d(n_1204), .o(n_1317) );
in01f80 g765291 ( .a(n_16060), .o(n_16061) );
na02f80 FE_RC_2367_0 ( .a(n_1596), .b(n_1597), .o(FE_RN_918_0) );
no02f80 g769759 ( .a(n_46423), .b(n_44453), .o(n_11200) );
oa12f80 g745206 ( .a(n_34355), .b(n_34492), .c(n_34384), .o(n_34572) );
in01f80 FE_RC_3841_0 ( .a(n_17247), .o(FE_RN_1674_0) );
oa12f80 g761709 ( .a(n_19400), .b(n_19401), .c(n_18694), .o(n_19486) );
na02f80 g766384 ( .a(n_14268), .b(n_14267), .o(n_14360) );
na02f80 g781026 ( .a(sin_out_18), .b(FE_OFN3_n_43918), .o(n_288) );
na02f80 g752614 ( .a(n_27568), .b(n_27403), .o(n_27614) );
oa22f80 g773696 ( .a(n_7226), .b(n_7161), .c(n_7236), .d(n_7162), .o(n_7288) );
ao12f80 g768320 ( .a(n_12515), .b(n_12514), .c(n_12513), .o(n_12965) );
na02f80 g739142 ( .a(n_40957), .b(n_40822), .o(n_40978) );
na02f80 g741264 ( .a(FE_OCP_RBN3579_n_44944), .b(n_38908), .o(n_39326) );
no02f80 g771543 ( .a(n_8796), .b(n_7657), .o(n_8845) );
na02f80 g745848 ( .a(n_34138), .b(n_34137), .o(n_34197) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_31_ ( .ck(newNet_3382), .d(n_27799), .o(delay_add_ln22_unr17_stage7_stallmux_q_31_) );
na02f80 FE_RC_4170_0 ( .a(FE_RN_1816_0), .b(FE_RN_1818_0), .o(n_18682) );
na02f80 g779033 ( .a(n_2163), .b(n_1883), .o(n_2195) );
no02f80 g781249 ( .a(n_100), .b(n_86), .o(n_270) );
oa12f80 g740873 ( .a(n_39326), .b(n_44309), .c(n_38940), .o(n_39374) );
no02f80 g778488 ( .a(n_2392), .b(n_2288), .o(n_2401) );
na02f80 g738315 ( .a(n_41833), .b(n_41832), .o(n_41834) );
in01f80 newInst_921 ( .a(newNet_920), .o(newNet_921) );
no02f80 g766997 ( .a(n_13558), .b(n_13017), .o(n_13592) );
na02f80 g769207 ( .a(n_11601), .b(n_11634), .o(n_12029) );
in01f80 FE_OCP_RBC2286_n_2433 ( .a(n_2433), .o(FE_OCP_RBN2286_n_2433) );
in01f80 g765917 ( .a(n_14872), .o(n_14932) );
ao22s80 g766401 ( .a(n_14355), .b(FE_OCP_RBN2503_n_13896), .c(n_16143), .d(FE_OCP_RBN2504_n_13896), .o(n_14533) );
no02f80 g742465 ( .a(n_37667), .b(n_37709), .o(n_37690) );
ao12f80 g783818 ( .a(n_8531), .b(n_8471), .c(n_7594), .o(n_45503) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_17_ ( .ck(newNet_3155), .d(n_40490), .o(delay_add_ln22_unr27_stage10_stallmux_q_17_) );
na02f80 g777303 ( .a(n_3564), .b(n_3563), .o(n_3565) );
ao22s80 FE_RC_3907_0 ( .a(n_30276), .b(n_30736), .c(n_30275), .d(n_30735), .o(n_30849) );
na02f80 g778231 ( .a(n_2775), .b(n_2740), .o(n_2826) );
no02f80 g739103 ( .a(n_41017), .b(n_41016), .o(n_41018) );
na02f80 g738029 ( .a(n_42151), .b(n_42102), .o(n_42152) );
no02f80 g745421 ( .a(FE_OCP_RBN2993_n_35539), .b(n_35629), .o(n_35630) );
in01f80 g762407 ( .a(n_18722), .o(n_18723) );
na02f80 g774929 ( .a(n_6139), .b(n_5900), .o(n_6190) );
in01f80 g760370 ( .a(n_20081), .o(n_20151) );
oa22f80 FE_RC_2474_0 ( .a(n_39247), .b(n_39477), .c(n_39478), .d(n_39248), .o(n_39559) );
in01f80 g780034 ( .a(n_1253), .o(n_1254) );
in01f80 newInst_1238 ( .a(newNet_652), .o(newNet_1238) );
in01f80 g779539 ( .a(n_1397), .o(n_1398) );
in01f80 g771891 ( .a(n_8786), .o(n_8787) );
ao22s80 FE_RC_1062_0 ( .a(n_1462), .b(n_1558), .c(n_792), .d(n_1780), .o(n_1590) );
no02f80 g770364 ( .a(n_10547), .b(n_10508), .o(n_10548) );
no02f80 g779599 ( .a(n_1852), .b(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .o(n_1882) );
na02f80 g765788 ( .a(n_14979), .b(n_14758), .o(n_15043) );
in01f80 g770764 ( .a(n_10290), .o(n_10347) );
ao12f80 g762455 ( .a(n_17975), .b(FE_OCP_RBN2142_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_14_), .o(n_18003) );
in01f80 FE_RC_1093_0 ( .a(n_17802), .o(FE_RN_322_0) );
no02f80 g751406 ( .a(n_28610), .b(n_28534), .o(n_28682) );
na02f80 g755544 ( .a(n_24719), .b(n_24497), .o(n_24778) );
in01f80 g760641 ( .a(n_19803), .o(n_19804) );
in01f80 newInst_3716 ( .a(newNet_3715), .o(newNet_3716) );
no02f80 g738737 ( .a(n_41483), .b(n_41228), .o(n_41530) );
ao12f80 g768479 ( .a(n_12372), .b(n_45659), .c(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .o(n_12642) );
in01f80 newInst_182 ( .a(newNet_181), .o(newNet_182) );
in01f80 FE_OCPC3751_n_44222 ( .a(FE_OCPN3750_n_44222), .o(FE_OCPN3751_n_44222) );
in01f80 g749230 ( .a(n_30847), .o(n_30910) );
oa12f80 g760413 ( .a(n_20034), .b(n_20033), .c(n_20032), .o(n_21788) );
oa12f80 g742150 ( .a(FE_OCP_RBN3452_n_37945), .b(n_37574), .c(n_37567), .o(n_38156) );
in01f80 g736526 ( .a(n_43701), .o(n_43711) );
na02f80 g745073 ( .a(n_34711), .b(n_34281), .o(n_34730) );
no02f80 g770158 ( .a(n_10902), .b(FE_OCP_RBN2704_n_9411), .o(n_10927) );
no02f80 g737415 ( .a(n_42734), .b(n_42712), .o(n_42752) );
in01f80 g768745 ( .a(n_12182), .o(n_12183) );
in01f80 FE_OCP_RBC2175_n_37559 ( .a(FE_OCP_RBN2174_n_37559), .o(FE_OCP_RBN2175_n_37559) );
in01f80 FE_OCPC1436_n_19855 ( .a(FE_OCPN1435_n_19855), .o(FE_OCPN1436_n_19855) );
in01f80 newInst_1311 ( .a(newNet_911), .o(newNet_1311) );
na02f80 g778109 ( .a(FE_OCP_RBN2414_n_2922), .b(n_2977), .o(n_3004) );
na02f80 g765083 ( .a(n_15275), .b(FE_OCPN1007_n_13962), .o(n_15425) );
no02f80 g769325 ( .a(FE_OCPN858_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(n_11970) );
no02f80 g754407 ( .a(n_25753), .b(n_25510), .o(n_25778) );
in01f80 g770193 ( .a(n_10821), .o(n_10788) );
in01f80 g754617 ( .a(FE_OCPN1410_n_27014), .o(n_27130) );
na02f80 g742232 ( .a(n_44887), .b(n_37929), .o(n_38247) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_5_ ( .ck(newNet_1568), .d(n_27000), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_) );
no02f80 g767627 ( .a(n_12949), .b(n_12769), .o(n_12950) );
ao12f80 g755465 ( .a(n_24781), .b(n_24780), .c(n_24779), .o(n_24848) );
oa12f80 g777948 ( .a(n_3073), .b(n_3072), .c(n_3071), .o(n_4632) );
in01f80 g775879 ( .a(n_5359), .o(n_5395) );
no02f80 g745418 ( .a(FE_OCP_RBN2993_n_35539), .b(n_34988), .o(n_35718) );
no02f80 g764637 ( .a(n_15945), .b(n_15937), .o(n_16154) );
in01f80 g763754 ( .a(n_16825), .o(n_16826) );
no02f80 g767061 ( .a(FE_OCP_RBN2458_n_13765), .b(n_13288), .o(n_13892) );
in01f80 g780226 ( .a(n_1065), .o(n_1049) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_28_ ( .ck(newNet_3507), .d(n_22857), .o(delay_add_ln22_unr14_stage6_stallmux_q_28_) );
no02f80 g741026 ( .a(n_39030), .b(n_39056), .o(n_39080) );
in01f80 g775732 ( .a(n_5340), .o(n_5382) );
in01f80 FE_OCP_RBC1204_n_26121 ( .a(n_26121), .o(FE_OCP_RBN1204_n_26121) );
in01f80 g742992 ( .a(n_36966), .o(n_36967) );
in01f80 g763288 ( .a(n_17043), .o(n_17044) );
in01f80 newInst_3531 ( .a(newNet_3530), .o(newNet_3531) );
no02f80 g742086 ( .a(FE_OCP_RBN3445_n_37945), .b(n_38235), .o(n_38255) );
na02f80 FE_RC_2300_0 ( .a(FE_RN_866_0), .b(FE_RN_867_0), .o(FE_RN_868_0) );
in01f80 g743190 ( .a(n_36923), .o(n_36888) );
in01f80 FE_OCP_RBC1699_n_19353 ( .a(n_19353), .o(FE_OCP_RBN1699_n_19353) );
ao12f80 g758957 ( .a(n_21448), .b(n_22011), .c(n_21516), .o(n_22061) );
no02f80 g761126 ( .a(n_19146), .b(n_19171), .o(n_19285) );
no02f80 g757965 ( .a(n_22660), .b(n_22649), .o(n_22738) );
ao12f80 g770292 ( .a(n_10571), .b(n_10478), .c(n_10548), .o(n_10667) );
na02f80 FE_RC_1058_0 ( .a(FE_RN_309_0), .b(FE_RN_310_0), .o(FE_RN_311_0) );
na02f80 g761462 ( .a(n_19609), .b(n_19608), .o(n_19709) );
na02f80 g764972 ( .a(n_15674), .b(n_15673), .o(n_15675) );
oa22f80 g778407 ( .a(n_2410), .b(n_2461), .c(n_2475), .d(n_2442), .o(n_2554) );
na02f80 FE_RC_1546_0 ( .a(FE_RN_435_0), .b(FE_RN_436_0), .o(FE_RN_437_0) );
in01f80 FE_OCPC1762_n_37877 ( .a(FE_OCPN1761_n_37877), .o(FE_OCPN1762_n_37877) );
no02f80 g753461 ( .a(n_27541), .b(n_26794), .o(n_27589) );
in01f80 g747830 ( .a(n_33601), .o(n_33572) );
in01f80 newInst_218 ( .a(newNet_30), .o(newNet_218) );
in01f80 newInst_3154 ( .a(newNet_3153), .o(newNet_3154) );
na02f80 g773675 ( .a(n_7314), .b(n_7313), .o(n_7315) );
in01f80 g765734 ( .a(n_15599), .o(n_15670) );
no02f80 FE_RC_2911_0 ( .a(n_13054), .b(n_13221), .o(FE_RN_1266_0) );
oa12f80 g780432 ( .a(n_872), .b(n_1203), .c(FE_OFN50_n_1045), .o(n_921) );
in01f80 g744718 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_12_), .o(n_36541) );
no02f80 g745943 ( .a(n_34086), .b(n_34085), .o(n_34134) );
oa12f80 g743774 ( .a(n_37262), .b(n_37283), .c(n_46230), .o(n_37304) );
no02f80 g760615 ( .a(n_19753), .b(n_19779), .o(n_19838) );
oa12f80 g736307 ( .a(n_308), .b(n_43867), .c(FE_OFN1_n_43918), .o(n_43906) );
na02f80 g781232 ( .a(n_107), .b(n_106), .o(n_108) );
in01f80 g748714 ( .a(n_31268), .o(n_31183) );
na02f80 FE_RC_2000_0 ( .a(n_19580), .b(FE_RN_655_0), .o(FE_RN_656_0) );
no02f80 g759123 ( .a(n_21367), .b(n_45026), .o(n_21389) );
oa12f80 g755518 ( .a(n_25469), .b(n_25468), .c(n_25467), .o(n_26307) );
ao22s80 FE_RC_3257_0 ( .a(n_9611), .b(n_9426), .c(n_9425), .d(n_9612), .o(n_9788) );
in01f80 g759895 ( .a(n_21379), .o(n_21298) );
na02f80 g769834 ( .a(n_11081), .b(n_10987), .o(n_11095) );
in01f80 g748921 ( .a(n_32491), .o(n_32405) );
oa22f80 FE_RC_431_0 ( .a(n_16423), .b(n_16419), .c(n_14577), .d(n_16426), .o(n_16526) );
in01f80 g767200 ( .a(n_14419), .o(n_14588) );
oa12f80 g772982 ( .a(n_7787), .b(n_7803), .c(n_7786), .o(n_7861) );
na02f80 g748821 ( .a(n_32377), .b(n_32423), .o(n_32503) );
no02f80 g740449 ( .a(n_39718), .b(n_39725), .o(n_39761) );
ao12f80 g746859 ( .a(n_33186), .b(FE_OCP_RBN3387_n_33108), .c(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n_33560) );
in01f80 newInst_2849 ( .a(newNet_2848), .o(newNet_2849) );
ao12f80 g762701 ( .a(n_17920), .b(FE_OCPN854_n_45450), .c(delay_xor_ln22_unr12_stage5_stallmux_q_17_), .o(n_17944) );
no02f80 g781173 ( .a(n_175), .b(n_170), .o(n_182) );
no02f80 g765032 ( .a(n_15285), .b(n_15241), .o(n_15387) );
in01f80 FE_OCPC1498_n_26360 ( .a(FE_OCPN1497_n_26360), .o(FE_OCPN1498_n_26360) );
no02f80 g765006 ( .a(n_15321), .b(n_15112), .o(n_15389) );
in01f80 g750018 ( .a(n_30218), .o(n_30219) );
oa12f80 g756835 ( .a(n_24034), .b(n_23989), .c(n_24188), .o(n_24736) );
na02f80 g773209 ( .a(n_7743), .b(n_7769), .o(n_7815) );
no02f80 FE_RC_3010_0 ( .a(FE_RN_1318_0), .b(n_20913), .o(n_20932) );
in01f80 newInst_364 ( .a(newNet_363), .o(newNet_364) );
in01f80 FE_OFC794_n_45813 ( .a(FE_OFN793_n_45813), .o(FE_OFN794_n_45813) );
ao12f80 g752205 ( .a(n_27916), .b(FE_OCPN877_n_44734), .c(delay_xor_ln22_unr18_stage7_stallmux_q_10_), .o(n_28290) );
oa12f80 g749110 ( .a(n_31016), .b(n_31046), .c(n_31045), .o(n_31123) );
in01f80 newInst_2623 ( .a(newNet_2622), .o(newNet_2623) );
in01f80 g740121 ( .a(n_40320), .o(n_40321) );
in01f80 g737188 ( .a(n_43003), .o(n_42997) );
na02f80 g745070 ( .a(n_34873), .b(n_34850), .o(n_34851) );
na02f80 g753252 ( .a(n_27098), .b(n_25808), .o(n_27143) );
no02f80 g773760 ( .a(n_7258), .b(n_7045), .o(n_7260) );
na02f80 g736919 ( .a(n_43038), .b(n_43037), .o(n_43385) );
in01f80 g741591 ( .a(n_38651), .o(n_38662) );
in01f80 FE_OCPC1446_n_31473 ( .a(FE_OCPN1445_n_31473), .o(FE_OCPN1446_n_31473) );
in01f80 g764601 ( .a(n_16003), .o(n_16038) );
na02f80 g763945 ( .a(n_16604), .b(n_16641), .o(n_16661) );
ao12f80 g747699 ( .a(n_33392), .b(n_33390), .c(n_33441), .o(n_33442) );
na02f80 g749126 ( .a(n_46957), .b(n_27246), .o(n_30861) );
ao12f80 g781266 ( .a(n_60), .b(n_46055), .c(beta_10), .o(n_96) );
oa12f80 g752720 ( .a(n_27068), .b(n_27128), .c(n_27073), .o(n_27239) );
in01f80 FE_OCPC955_n_44460 ( .a(FE_OCPN954_n_44460), .o(FE_OCPN955_n_44460) );
in01f80 g755710 ( .a(n_24471), .o(n_24567) );
na02f80 g751040 ( .a(n_30065), .b(n_30028), .o(n_30066) );
no02f80 g754012 ( .a(n_26129), .b(n_26128), .o(n_26158) );
na02f80 g737011 ( .a(FE_OCP_RBN3072_n_43230), .b(n_46935), .o(n_43430) );
na02f80 g740797 ( .a(n_39354), .b(n_38984), .o(n_39384) );
no02f80 g755795 ( .a(n_25256), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25257) );
ao12f80 g755372 ( .a(FE_OCPN1512_n_22280), .b(n_24875), .c(n_24874), .o(n_24896) );
ao12f80 g769240 ( .a(n_11863), .b(n_11707), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_), .o(n_12485) );
ms00f80 sin_out_reg_8_ ( .ck(newNet_11), .d(n_43746), .o(sin_out_8) );
na02f80 g745546 ( .a(n_34167), .b(n_34153), .o(n_34154) );
in01f80 g768981 ( .a(n_11817), .o(n_11818) );
in01f80 FE_OCPC1410_n_27014 ( .a(FE_OCPN1409_n_27014), .o(FE_OCPN1410_n_27014) );
oa22f80 g745344 ( .a(n_35956), .b(n_36111), .c(FE_OCP_RBN2995_n_35539), .d(n_35602), .o(n_36229) );
na02f80 g737572 ( .a(n_42449), .b(n_42448), .o(n_42450) );
oa12f80 g747635 ( .a(n_32052), .b(n_47205), .c(n_32326), .o(n_32345) );
ao12f80 g747975 ( .a(n_33047), .b(n_33046), .c(n_33045), .o(n_33552) );
na02f80 g765926 ( .a(n_14785), .b(n_14758), .o(n_14880) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_0_ ( .ck(newNet_3571), .d(n_20715), .o(delay_add_ln22_unr14_stage6_stallmux_q_0_) );
in01f80 g737912 ( .a(n_42545), .o(n_42546) );
na02f80 g780744 ( .a(n_594), .b(n_593), .o(n_595) );
in01f80 g753742 ( .a(n_26522), .o(n_26523) );
no02f80 g773578 ( .a(n_7456), .b(n_7455), .o(n_7457) );
no02f80 g745034 ( .a(n_34853), .b(n_34372), .o(n_34900) );
in01f80 g751503 ( .a(n_28732), .o(n_28733) );
in01f80 FE_OCPC1055_n_14098 ( .a(FE_OCPN1053_n_14098), .o(FE_OCPN1055_n_14098) );
no02f80 g763770 ( .a(n_17105), .b(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17210) );
no02f80 g758758 ( .a(n_21660), .b(n_21659), .o(n_21682) );
in01f80 g761780 ( .a(n_18562), .o(n_18563) );
oa12f80 g775463 ( .a(n_4746), .b(n_5716), .c(n_4921), .o(n_5775) );
na02f80 g745980 ( .a(n_33962), .b(n_33836), .o(n_33983) );
in01f80 g755228 ( .a(n_25178), .o(n_25173) );
no02f80 g767282 ( .a(n_13456), .b(n_13388), .o(n_13488) );
in01f80 FE_OCPC973_n_15900 ( .a(FE_OCPN972_n_15900), .o(FE_OCPN973_n_15900) );
in01f80 g777355 ( .a(n_4622), .o(n_4746) );
na03f80 g755620 ( .a(n_24498), .b(n_24500), .c(n_23943), .o(n_24527) );
ao12f80 g779424 ( .a(n_1705), .b(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_7_), .o(n_1711) );
na02f80 g740543 ( .a(n_39697), .b(n_39694), .o(n_39715) );
in01f80 g740089 ( .a(n_40136), .o(n_40189) );
ao12f80 g751066 ( .a(n_28501), .b(n_28852), .c(n_28547), .o(n_28869) );
na02f80 g781175 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_2_), .o(n_177) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_1_ ( .ck(newNet_1013), .d(n_16700), .o(n_44721) );
na02f80 g767303 ( .a(n_13675), .b(n_13674), .o(n_13676) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_15_ ( .ck(newNet_2309), .d(n_40405), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_) );
no02f80 g740188 ( .a(FE_OCP_RBN3052_n_39913), .b(n_40005), .o(n_40110) );
na02f80 g749024 ( .a(n_31048), .b(n_30931), .o(n_31078) );
no02f80 g741235 ( .a(n_39149), .b(n_39091), .o(n_39173) );
in01f80 newInst_1541 ( .a(newNet_583), .o(newNet_1541) );
in01f80 g747606 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_19_), .o(n_32222) );
in01f80 g769844 ( .a(n_11213), .o(n_11214) );
na02f80 g779228 ( .a(n_1845), .b(n_1844), .o(n_2008) );
in01f80 g741118 ( .a(n_39205), .o(n_39206) );
in01f80 g749782 ( .a(n_31429), .o(n_31430) );
in01f80 g755612 ( .a(FE_OCP_RBN2405_n_24638), .o(n_24959) );
no02f80 g749831 ( .a(n_31044), .b(n_31043), .o(n_31118) );
no02f80 g763240 ( .a(n_17127), .b(n_17188), .o(n_17241) );
no02f80 g760836 ( .a(n_20056), .b(n_20058), .o(n_20137) );
no02f80 g777369 ( .a(n_3638), .b(n_2359), .o(n_3725) );
na02f80 FE_RC_3653_0 ( .a(FE_RN_1603_0), .b(n_22037), .o(n_22064) );
in01f80 newInst_3391 ( .a(newNet_3390), .o(newNet_3391) );
in01f80 g751897 ( .a(n_29070), .o(n_29128) );
no02f80 g778671 ( .a(n_2289), .b(n_2292), .o(n_2348) );
no02f80 g748220 ( .a(FE_OCP_RBN3732_n_31819), .b(n_32076), .o(n_32077) );
na02f80 g780288 ( .a(n_910), .b(n_1159), .o(n_911) );
oa12f80 g747848 ( .a(n_31611), .b(n_32003), .c(n_31605), .o(n_32061) );
in01f80 g776998 ( .a(n_4198), .o(n_4199) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_25_ ( .ck(newNet_2088), .d(n_6500), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_25_) );
in01f80 FE_OCP_RBC2545_n_44944 ( .a(n_44944), .o(FE_OCP_RBN2545_n_44944) );
in01f80 g771486 ( .a(n_9523), .o(n_9524) );
no02f80 g759749 ( .a(n_21479), .b(n_21403), .o(n_22060) );
in01f80 newInst_1226 ( .a(newNet_520), .o(newNet_1226) );
in01f80 g737612 ( .a(n_42487), .o(n_42488) );
in01f80 FE_OCP_RBC2454_n_14157 ( .a(n_14157), .o(FE_OCP_RBN2454_n_14157) );
in01f80 g770996 ( .a(n_10031), .o(n_10164) );
oa12f80 g755156 ( .a(n_24961), .b(n_25049), .c(n_24913), .o(n_25118) );
na02f80 g739206 ( .a(n_40687), .b(n_40689), .o(n_40708) );
no02f80 g747951 ( .a(n_33092), .b(n_33091), .o(n_33093) );
in01f80 g765166 ( .a(n_15275), .o(n_15347) );
no02f80 g753635 ( .a(n_26597), .b(n_26596), .o(n_26628) );
oa22f80 g739754 ( .a(n_40425), .b(n_40079), .c(n_40426), .d(n_40078), .o(n_40464) );
na02f80 g740002 ( .a(n_40141), .b(n_40073), .o(n_40192) );
in01f80 g759672 ( .a(n_20721), .o(n_20722) );
no02f80 g766892 ( .a(n_13847), .b(n_14210), .o(n_14455) );
no02f80 g743342 ( .a(n_36715), .b(n_36750), .o(n_36777) );
oa22f80 g758197 ( .a(n_22604), .b(n_21867), .c(n_22605), .d(n_21868), .o(n_22689) );
na03f80 g779261 ( .a(n_1550), .b(n_1806), .c(n_1527), .o(n_1820) );
oa22f80 g776460 ( .a(n_4158), .b(n_3029), .c(FE_OCP_RBN2667_n_4158), .d(n_4093), .o(n_4346) );
oa22f80 g746872 ( .a(FE_OCP_RBN2169_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_31_), .c(FE_OCP_RBN2172_n_32892), .d(n_32542), .o(n_33213) );
na02f80 FE_RC_1206_0 ( .a(FE_RN_365_0), .b(n_16902), .o(n_17522) );
na02f80 g760536 ( .a(n_19896), .b(n_19895), .o(n_19897) );
in01f80 g775885 ( .a(n_5323), .o(n_5285) );
no02f80 g776533 ( .a(n_4138), .b(n_4125), .o(n_4294) );
na02f80 g739564 ( .a(n_40622), .b(n_40647), .o(n_40651) );
no02f80 g745287 ( .a(n_35805), .b(n_35804), .o(n_35806) );
in01f80 g772975 ( .a(n_7835), .o(n_7836) );
na02f80 g746213 ( .a(n_33753), .b(n_33324), .o(n_33772) );
in01f80 g741098 ( .a(n_39500), .o(n_39501) );
in01f80 g746359 ( .a(n_33541), .o(n_34314) );
ao12f80 g741852 ( .a(n_38411), .b(n_38410), .c(n_38409), .o(n_38859) );
oa12f80 g765922 ( .a(n_14664), .b(n_14696), .c(n_14611), .o(n_14775) );
in01f80 g775679 ( .a(n_5571), .o(n_5611) );
no02f80 g753982 ( .a(n_26186), .b(n_26293), .o(n_26187) );
in01f80 g736855 ( .a(n_43617), .o(n_43618) );
na02f80 g753974 ( .a(n_26977), .b(n_26612), .o(n_27035) );
na02f80 g773554 ( .a(n_7423), .b(n_7385), .o(n_7430) );
na02f80 g761189 ( .a(FE_OCP_RBN1685_n_18986), .b(n_17783), .o(n_19044) );
in01f80 FE_RC_1813_0 ( .a(FE_RN_539_0), .o(n_17791) );
no02f80 g757718 ( .a(n_22559), .b(n_22539), .o(n_22613) );
na02f80 g763133 ( .a(n_17480), .b(n_17443), .o(n_17620) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_25_ ( .ck(newNet_321), .d(n_1356), .o(delay_xor_ln22_unr3_stage2_stallmux_q_25_) );
na02f80 g739186 ( .a(n_40911), .b(n_40860), .o(n_40912) );
in01f80 newInst_2476 ( .a(newNet_2475), .o(newNet_2476) );
oa12f80 g763027 ( .a(n_17056), .b(n_17863), .c(n_17530), .o(n_17984) );
in01f80 newInst_2043 ( .a(newNet_1681), .o(newNet_2043) );
in01f80 newInst_695 ( .a(newNet_694), .o(newNet_695) );
no02f80 g752634 ( .a(n_27554), .b(n_27168), .o(n_27590) );
oa22f80 FE_RC_4119_0 ( .a(n_22820), .b(n_22746), .c(n_22595), .d(n_22747), .o(n_22899) );
na02f80 g749852 ( .a(n_31311), .b(n_31223), .o(n_31508) );
no02f80 g764970 ( .a(n_15389), .b(n_15391), .o(n_15434) );
in01f80 fopt783254 ( .a(n_9676), .o(n_44819) );
na02f80 g750428 ( .a(FE_OCP_RBN3491_n_29553), .b(n_29630), .o(n_29579) );
in01f80 newInst_2359 ( .a(newNet_2358), .o(newNet_2359) );
no02f80 g740920 ( .a(n_39114), .b(n_38881), .o(n_39167) );
ao12f80 g746337 ( .a(n_34867), .b(n_34868), .c(n_34545), .o(n_34944) );
na02f80 g777709 ( .a(n_3413), .b(n_3384), .o(n_3474) );
in01f80 FE_OCP_RBC2553_n_44921 ( .a(n_44921), .o(FE_OCP_RBN2553_n_44921) );
in01f80 FE_OCP_RBC3387_n_33108 ( .a(FE_OCP_RBN3386_n_33108), .o(FE_OCP_RBN3387_n_33108) );
in01f80 g765870 ( .a(n_15212), .o(n_15289) );
in01f80 FE_OCP_RBC3624_n_38870 ( .a(FE_OCP_RBN2685_n_38870), .o(FE_OCP_RBN3624_n_38870) );
oa22f80 FE_RC_3267_0 ( .a(n_21132), .b(n_44718), .c(FE_OCP_RBN2880_n_21132), .d(n_44717), .o(n_21285) );
na02f80 g775021 ( .a(n_6056), .b(n_6048), .o(n_6154) );
no02f80 g748749 ( .a(n_32537), .b(n_32449), .o(n_33091) );
na02f80 g766020 ( .a(n_14638), .b(FE_OCP_RBN3528_n_13765), .o(n_14667) );
ao12f80 g773716 ( .a(n_6733), .b(n_7270), .c(n_6717), .o(n_7298) );
no02f80 g773123 ( .a(n_7627), .b(n_7613), .o(n_7693) );
in01f80 g753617 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .o(n_27285) );
oa12f80 g779806 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_8_), .o(n_1601) );
na02f80 g766832 ( .a(n_14381), .b(n_14301), .o(n_14423) );
oa22f80 FE_RC_3868_0 ( .a(n_27868), .b(n_27825), .c(n_27751), .d(n_27826), .o(n_28009) );
na02f80 g758077 ( .a(n_44267), .b(FE_OCP_RBN1723_n_21004), .o(n_22266) );
in01f80 newInst_229 ( .a(newNet_228), .o(newNet_229) );
no02f80 g740341 ( .a(n_40128), .b(n_40240), .o(n_40353) );
no02f80 g756375 ( .a(n_24016), .b(n_23738), .o(n_24017) );
in01f80 g749147 ( .a(n_30875), .o(n_30876) );
oa12f80 g767490 ( .a(n_13142), .b(n_13227), .c(n_13295), .o(n_13400) );
in01f80 g745645 ( .a(n_34151), .o(n_34152) );
no02f80 g780545 ( .a(FE_OCPN852_n_694), .b(n_46055), .o(n_831) );
in01f80 FE_RC_2510_0 ( .a(n_17891), .o(FE_RN_1021_0) );
in01f80 g774142 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .o(n_7595) );
no02f80 g764589 ( .a(n_16180), .b(n_16108), .o(n_16268) );
in01f80 newInst_3547 ( .a(newNet_2787), .o(newNet_3547) );
ao12f80 g762974 ( .a(n_17542), .b(n_17939), .c(n_17364), .o(n_17994) );
oa22f80 g743738 ( .a(n_36207), .b(n_35788), .c(n_36206), .d(n_35787), .o(n_36310) );
no02f80 g744524 ( .a(n_35421), .b(n_35420), .o(n_35465) );
in01f80 FE_OCP_DRV_C3739_n_29439 ( .a(FE_OCP_DRV_N3738_n_29439), .o(FE_OCP_DRV_N3739_n_29439) );
oa12f80 g777965 ( .a(n_2593), .b(n_3022), .c(n_2603), .o(n_3111) );
oa12f80 g743210 ( .a(n_36905), .b(n_36904), .c(n_36903), .o(n_37661) );
in01f80 FE_RC_4090_0 ( .a(FE_RN_1788_0), .o(FE_RN_1784_0) );
in01f80 g766003 ( .a(n_14783), .o(n_14784) );
in01f80 g739833 ( .a(n_40448), .o(n_40449) );
na02f80 g751999 ( .a(n_28897), .b(n_28837), .o(n_29043) );
in01f80 FE_RC_2177_0 ( .a(n_26202), .o(FE_RN_777_0) );
no02f80 g737406 ( .a(n_42737), .b(n_42429), .o(n_42811) );
na02f80 g756644 ( .a(n_23576), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .o(n_23636) );
no02f80 g773454 ( .a(n_7527), .b(n_6765), .o(n_7533) );
na02f80 g768340 ( .a(n_12509), .b(n_12508), .o(n_12510) );
ao12f80 g772739 ( .a(n_8161), .b(n_8169), .c(n_8160), .o(n_9220) );
no02f80 g747743 ( .a(n_33372), .b(n_33670), .o(n_33951) );
in01f80 g775717 ( .a(n_5313), .o(n_5314) );
in01f80 FE_OCPC874_n_44672 ( .a(FE_OCPN873_n_44672), .o(FE_OCPN874_n_44672) );
in01f80 newInst_1589 ( .a(newNet_1588), .o(newNet_1589) );
no02f80 g750825 ( .a(n_29095), .b(n_28774), .o(n_29116) );
in01f80 g770572 ( .a(n_10101), .o(n_10195) );
in01f80 g738963 ( .a(n_41191), .o(n_41194) );
in01f80 g754278 ( .a(n_25934), .o(n_25933) );
na02f80 g760735 ( .a(n_19538), .b(FE_OCPN1800_FE_OFN780_n_17093), .o(n_19568) );
in01f80 g738219 ( .a(n_41960), .o(n_41961) );
in01f80 g745976 ( .a(n_34064), .o(n_34049) );
ao12f80 g754128 ( .a(n_26812), .b(n_26947), .c(n_26866), .o(n_26952) );
in01f80 newInst_790 ( .a(newNet_789), .o(newNet_790) );
no02f80 g777907 ( .a(n_3189), .b(FE_OCP_RBN2345_FE_OCPN870_n_2737), .o(n_3241) );
no02f80 g760483 ( .a(n_20020), .b(FE_OCP_RBN1155_n_18375), .o(n_20093) );
in01f80 newInst_3248 ( .a(newNet_3247), .o(newNet_3248) );
no02f80 g769585 ( .a(n_47182), .b(n_11394), .o(n_11395) );
na02f80 g737585 ( .a(n_42747), .b(n_42726), .o(n_42769) );
na02f80 g761064 ( .a(n_19116), .b(n_18428), .o(n_19154) );
in01f80 g743990 ( .a(n_36332), .o(n_36333) );
no02f80 FE_RC_348_0 ( .a(FE_RN_101_0), .b(n_11962), .o(n_47211) );
in01f80 g776018 ( .a(n_5098), .o(n_5099) );
in01f80 fopt783338 ( .a(n_38830), .o(n_44921) );
no02f80 g743511 ( .a(FE_OCP_RBN3342_delay_add_ln22_unr23_stage9_stallmux_q_24_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .o(n_36903) );
no02f80 g743876 ( .a(n_36204), .b(n_36245), .o(n_36307) );
ao12f80 g745111 ( .a(n_34591), .b(n_34767), .c(FE_OCP_RBN3541_n_34487), .o(n_34786) );
ao12f80 g747202 ( .a(n_33914), .b(n_33913), .c(n_33912), .o(n_34472) );
in01f80 FE_RC_2335_0 ( .a(n_18524), .o(FE_RN_892_0) );
in01f80 g739804 ( .a(n_40422), .o(n_40456) );
in01f80 newInst_3573 ( .a(newNet_3572), .o(newNet_3573) );
ao12f80 g757705 ( .a(n_22345), .b(n_22513), .c(n_22046), .o(n_22566) );
in01f80 g751813 ( .a(n_29103), .o(n_29104) );
no02f80 g745963 ( .a(n_34059), .b(n_34058), .o(n_34111) );
in01f80 g763702 ( .a(n_16758), .o(n_16782) );
na02f80 g737783 ( .a(n_42302), .b(n_42321), .o(n_42303) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_4_ ( .ck(newNet_1284), .d(n_740), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_4_) );
no02f80 g766868 ( .a(n_13556), .b(n_13017), .o(n_13595) );
oa12f80 g781143 ( .a(beta_12), .b(n_206), .c(n_59), .o(n_205) );
in01f80 g748306 ( .a(n_31736), .o(n_31737) );
in01f80 newInst_372 ( .a(newNet_371), .o(newNet_372) );
in01f80 newInst_1858 ( .a(newNet_1857), .o(newNet_1858) );
no02f80 g760609 ( .a(n_19784), .b(n_19703), .o(n_19785) );
na02f80 g781012 ( .a(cos_out_7), .b(FE_OFN2_n_43918), .o(n_287) );
no02f80 FE_RC_4245_0 ( .a(FE_RN_1865_0), .b(FE_RN_1866_0), .o(FE_RN_1867_0) );
in01f80 FE_OCP_RBC2895_n_39575 ( .a(FE_OCP_RBN2894_n_39575), .o(FE_OCP_RBN2895_n_39575) );
no02f80 g746832 ( .a(n_33401), .b(n_33061), .o(n_33452) );
in01f80 FE_RC_3761_0 ( .a(n_40737), .o(FE_RN_1652_0) );
ao12f80 g746508 ( .a(n_33167), .b(n_33168), .c(n_33166), .o(n_33221) );
no02f80 g762875 ( .a(FE_OCP_RBN2141_FE_OCPN861_n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_11_), .o(n_17885) );
na02f80 g755448 ( .a(n_24826), .b(n_24825), .o(n_24851) );
na02f80 g753771 ( .a(n_26413), .b(n_26412), .o(n_26414) );
no02f80 g778170 ( .a(n_2859), .b(n_2858), .o(n_2907) );
na02f80 g773500 ( .a(n_8302), .b(n_7484), .o(n_7519) );
in01f80 g758509 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n_22620) );
na02f80 g763103 ( .a(n_17561), .b(n_17346), .o(n_17448) );
in01f80 newInst_3285 ( .a(newNet_3284), .o(newNet_3285) );
in01f80 newInst_2908 ( .a(newNet_2907), .o(newNet_2908) );
na02f80 g777260 ( .a(n_3485), .b(n_2770), .o(n_3504) );
na02f80 g748322 ( .a(n_31702), .b(FE_OCPN975_n_46956), .o(n_31705) );
no02f80 g749492 ( .a(n_30411), .b(n_30050), .o(n_30453) );
in01f80 newInst_392 ( .a(newNet_221), .o(newNet_392) );
in01f80 g748631 ( .a(n_31305), .o(n_31306) );
ao12f80 FE_RC_2560_0 ( .a(FE_RN_1048_0), .b(FE_RN_1049_0), .c(n_6835), .o(n_6945) );
no02f80 g767507 ( .a(n_13058), .b(n_13144), .o(n_13145) );
no02f80 g736978 ( .a(FE_OCPN1246_n_43120), .b(n_43070), .o(n_43507) );
na02f80 g749190 ( .a(n_30829), .b(FE_OCPN1486_n_27315), .o(n_30913) );
na02f80 g781110 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_7_), .o(n_257) );
na02f80 g761634 ( .a(n_18796), .b(n_18757), .o(n_18893) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_6_ ( .ck(newNet_212), .d(n_46164), .o(delay_xor_ln22_unr6_stage3_stallmux_q_6_) );
no02f80 g744494 ( .a(n_35425), .b(n_35344), .o(n_35455) );
no02f80 g755476 ( .a(n_24619), .b(FE_OCPN1482_n_22207), .o(n_24696) );
in01f80 g736808 ( .a(n_43462), .o(n_43463) );
in01f80 g746588 ( .a(n_34757), .o(n_34758) );
oa22f80 FE_RC_3788_0 ( .a(n_20716), .b(n_20877), .c(n_20960), .d(n_20876), .o(n_20903) );
in01f80 g765216 ( .a(n_15243), .o(n_15305) );
no02f80 g773140 ( .a(n_7617), .b(n_7881), .o(n_7689) );
in01f80 newInst_1639 ( .a(newNet_1465), .o(newNet_1639) );
oa12f80 g773926 ( .a(n_7255), .b(n_7217), .c(delay_xor_ln21_unr6_stage3_stallmux_q_25_), .o(n_7294) );
no02f80 g773562 ( .a(n_7439), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .o(n_7460) );
no02f80 g739357 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n_40909) );
in01f80 g756005 ( .a(n_25003), .o(n_24982) );
in01f80 g775537 ( .a(n_5465), .o(n_5466) );
in01f80 g746601 ( .a(n_34644), .o(n_34586) );
no02f80 g757331 ( .a(n_23067), .b(n_23066), .o(n_23068) );
no02f80 g755111 ( .a(n_25201), .b(n_25228), .o(n_25293) );
oa22f80 g765172 ( .a(n_15055), .b(n_14928), .c(n_15056), .d(n_14953), .o(n_15200) );
in01f80 g769488 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_20_), .o(n_11524) );
no02f80 FE_RC_3386_0 ( .a(FE_RN_1466_0), .b(FE_RN_1467_0), .o(FE_RN_1468_0) );
no02f80 g748887 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32483) );
na02f80 g776737 ( .a(n_4024), .b(n_4105), .o(n_4300) );
in01f80 FE_OCP_RBC3378_n_40716 ( .a(n_40716), .o(FE_OCP_RBN3378_n_40716) );
in01f80 g757894 ( .a(n_23812), .o(n_23869) );
in01f80 g765379 ( .a(n_16016), .o(n_16102) );
in01f80 g780911 ( .a(n_480), .o(n_458) );
in01f80 g762841 ( .a(n_17843), .o(n_17910) );
na02f80 g743467 ( .a(n_36505), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36539) );
in01f80 newInst_1511 ( .a(newNet_1510), .o(newNet_1511) );
in01f80 g745872 ( .a(n_35388), .o(n_35389) );
na02f80 g754158 ( .a(n_26947), .b(n_26946), .o(n_26948) );
na02f80 g764110 ( .a(n_16565), .b(n_16564), .o(n_16566) );
in01f80 newInst_305 ( .a(newNet_304), .o(newNet_305) );
in01f80 g741702 ( .a(n_38577), .o(n_38578) );
na02f80 g744146 ( .a(n_35776), .b(n_35899), .o(n_35945) );
na02f80 g753512 ( .a(n_26779), .b(n_26421), .o(n_26826) );
in01f80 g741837 ( .a(n_38420), .o(n_38388) );
in01f80 g764043 ( .a(n_17881), .o(n_17900) );
na02f80 g778742 ( .a(n_2289), .b(n_2292), .o(n_2402) );
no02f80 g740053 ( .a(n_40015), .b(n_46950), .o(n_39952) );
no02f80 g772275 ( .a(n_8736), .b(n_8735), .o(n_8737) );
in01f80 newInst_3325 ( .a(newNet_3324), .o(newNet_3325) );
in01f80 newInst_74 ( .a(newNet_60), .o(newNet_74) );
in01f80 g768034 ( .a(n_13113), .o(n_13114) );
in01f80 newInst_68 ( .a(newNet_39), .o(newNet_68) );
in01f80 newInst_2528 ( .a(newNet_2527), .o(newNet_2528) );
in01f80 newInst_998 ( .a(newNet_997), .o(newNet_998) );
oa22f80 g737863 ( .a(n_42270), .b(n_42137), .c(n_42547), .d(n_42113), .o(n_42673) );
na02f80 g745784 ( .a(n_34147), .b(n_34126), .o(n_34223) );
no02f80 g760552 ( .a(n_19868), .b(n_19861), .o(n_19944) );
na02f80 g779299 ( .a(n_1701), .b(n_1032), .o(n_1785) );
in01f80 g737550 ( .a(n_42472), .o(n_42473) );
na02f80 g754317 ( .a(n_25889), .b(n_23317), .o(n_25911) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_1_ ( .ck(newNet_726), .d(n_46174), .o(delay_xor_ln21_unr6_stage3_stallmux_q_1_) );
na02f80 g776458 ( .a(n_4464), .b(n_4327), .o(n_4465) );
no02f80 FE_RC_3515_0 ( .a(n_28342), .b(n_28343), .o(FE_RN_1518_0) );
in01f80 fopt783173 ( .a(n_44711), .o(n_44710) );
na02f80 g768401 ( .a(n_12449), .b(n_11976), .o(n_12471) );
na02f80 g763833 ( .a(n_16611), .b(n_16465), .o(n_16629) );
na02f80 g764749 ( .a(n_46981), .b(n_15935), .o(n_15980) );
no02f80 g777324 ( .a(n_4182), .b(FE_OFN818_n_4575), .o(n_4598) );
oa22f80 FE_RC_3879_0 ( .a(n_24469), .b(n_44621), .c(n_24450), .d(n_24862), .o(n_24945) );
na02f80 g757189 ( .a(n_23133), .b(n_23171), .o(n_23309) );
na02f80 g745572 ( .a(n_34297), .b(n_33539), .o(n_34351) );
in01f80 g748497 ( .a(n_31549), .o(n_31612) );
na02f80 FE_RC_2294_0 ( .a(FE_RN_862_0), .b(n_28130), .o(FE_RN_863_0) );
na02f80 g739348 ( .a(n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n_40675) );
na02f80 g774839 ( .a(n_6228), .b(n_5706), .o(n_6362) );
na02f80 g780073 ( .a(n_1215), .b(n_811), .o(n_1222) );
no02f80 g740893 ( .a(n_44309), .b(n_39049), .o(n_39380) );
in01f80 g750481 ( .a(n_29568), .o(n_29569) );
no02f80 g746243 ( .a(n_33644), .b(n_33581), .o(n_33645) );
in01f80 g745940 ( .a(n_34109), .o(n_34110) );
na02f80 g747823 ( .a(n_33238), .b(n_33294), .o(n_33417) );
in01f80 newInst_737 ( .a(newNet_736), .o(newNet_737) );
in01f80 g743295 ( .a(n_37504), .o(n_36768) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_4_ ( .ck(newNet_411), .d(n_32565), .o(delay_xor_ln22_unr21_stage8_stallmux_q_4_) );
in01f80 g740506 ( .a(n_39717), .o(n_39718) );
na02f80 g753206 ( .a(n_27204), .b(n_25928), .o(n_27426) );
ao12f80 g770395 ( .a(n_10566), .b(n_10575), .c(n_10565), .o(n_10636) );
oa22f80 FE_RC_3325_0 ( .a(n_12837), .b(n_13631), .c(n_12862), .d(n_13632), .o(n_13726) );
in01f80 drc784129 ( .a(n_45879), .o(n_45880) );
ao12f80 g751925 ( .a(n_29223), .b(n_28897), .c(n_28923), .o(n_29286) );
na02f80 g770514 ( .a(n_10230), .b(n_10153), .o(n_10318) );
na02f80 g759308 ( .a(FE_OCP_RBN1724_n_21004), .b(FE_OCP_RBN1914_n_20965), .o(n_21076) );
na02f80 g760132 ( .a(n_20456), .b(FE_OCP_RBN3839_n_19513), .o(n_20573) );
in01f80 newInst_3498 ( .a(newNet_2593), .o(newNet_3498) );
no02f80 FE_RC_3008_0 ( .a(FE_RN_713_0), .b(n_30818), .o(FE_RN_1317_0) );
no02f80 g762379 ( .a(FE_OCP_RBN3410_n_45120), .b(n_18251), .o(n_18585) );
no02f80 g746934 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_14_), .o(n_32914) );
in01f80 newInst_1257 ( .a(newNet_344), .o(newNet_1257) );
no02f80 g758283 ( .a(n_22003), .b(n_22002), .o(n_22018) );
na02f80 g780711 ( .a(n_628), .b(n_627), .o(n_629) );
in01f80 fopt783444 ( .a(n_45010), .o(n_45013) );
in01f80 newInst_2752 ( .a(newNet_1979), .o(newNet_2752) );
na02f80 g784595 ( .a(n_8493), .b(n_8346), .o(n_46418) );
in01f80 g756030 ( .a(n_25030), .o(n_25083) );
in01f80 g743608 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_17_), .o(n_36486) );
in01f80 g756261 ( .a(FE_OCP_RBN2278_n_24173), .o(n_24217) );
na02f80 g746614 ( .a(n_34473), .b(n_34474), .o(n_34760) );
in01f80 newInst_3607 ( .a(newNet_277), .o(newNet_3607) );
in01f80 g774719 ( .a(n_6376), .o(n_6365) );
na02f80 g740759 ( .a(n_39535), .b(n_40183), .o(n_39534) );
no02f80 g767553 ( .a(n_13216), .b(n_13215), .o(n_13217) );
in01f80 FE_OCP_RBC2117_n_45224 ( .a(FE_OCP_RBN3266_n_45224), .o(FE_OCP_RBN2117_n_45224) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_9_ ( .ck(newNet_1562), .d(n_27002), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_9_) );
na02f80 g738875 ( .a(n_41231), .b(n_41230), .o(n_41232) );
na02f80 g765622 ( .a(n_15074), .b(n_15040), .o(n_15224) );
in01f80 g768065 ( .a(n_12718), .o(n_12719) );
in01f80 newInst_1404 ( .a(newNet_637), .o(newNet_1404) );
in01f80 FE_OCPC1402_n_9642 ( .a(FE_OCPN1401_n_9642), .o(FE_OCPN1402_n_9642) );
na02f80 g763342 ( .a(n_17180), .b(n_17217), .o(n_17376) );
na02f80 g760955 ( .a(n_19327), .b(n_18937), .o(n_19332) );
in01f80 g774948 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_17_), .o(n_6167) );
no02f80 FE_RC_1995_0 ( .a(n_19374), .b(n_19420), .o(FE_RN_653_0) );
in01f80 g761959 ( .a(n_18405), .o(n_18397) );
na02f80 g740608 ( .a(n_39636), .b(n_45841), .o(n_39661) );
na02f80 g740620 ( .a(n_39617), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39652) );
in01f80 newInst_2011 ( .a(newNet_1353), .o(newNet_2011) );
no02f80 g751300 ( .a(n_29654), .b(n_29653), .o(n_29655) );
na02f80 g763411 ( .a(n_16838), .b(n_16874), .o(n_16950) );
in01f80 g758799 ( .a(n_21615), .o(n_21708) );
no02f80 g773150 ( .a(n_7802), .b(n_7848), .o(n_7909) );
na02f80 g756398 ( .a(n_24216), .b(n_23898), .o(n_24277) );
na02f80 FE_RC_2535_0 ( .a(n_36234), .b(n_36490), .o(FE_RN_1034_0) );
in01f80 FE_OCP_RBC3512_n_13960 ( .a(FE_OCP_RBN2411_n_13960), .o(FE_OCP_RBN3512_n_13960) );
in01f80 g772574 ( .a(n_8398), .o(n_8399) );
na02f80 g737751 ( .a(n_42341), .b(n_42384), .o(n_42385) );
in01f80 g769230 ( .a(n_11715), .o(n_11677) );
no02f80 g740403 ( .a(FE_OCP_RBN3022_n_39942), .b(n_39992), .o(n_40241) );
no02f80 g736694 ( .a(n_43234), .b(n_43150), .o(n_43235) );
in01f80 g741100 ( .a(n_39528), .o(n_39529) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_16_ ( .ck(newNet_3328), .d(n_32029), .o(delay_add_ln22_unr20_stage8_stallmux_q_16_) );
na02f80 g761071 ( .a(n_19110), .b(n_17900), .o(n_19120) );
in01f80 newInst_2539 ( .a(newNet_2538), .o(newNet_2539) );
in01f80 fopt783088 ( .a(n_44566), .o(n_44563) );
in01f80 g739299 ( .a(n_40831), .o(n_40765) );
oa22f80 g743639 ( .a(n_36424), .b(n_36332), .c(n_36425), .d(n_36333), .o(n_36469) );
ao12f80 g746843 ( .a(n_33323), .b(FE_OCP_RBN3384_n_33108), .c(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n_33366) );
oa12f80 g780335 ( .a(n_716), .b(n_715), .c(n_714), .o(n_738) );
no02f80 g748880 ( .a(n_32356), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(n_32376) );
na02f80 g751871 ( .a(n_28248), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_6_), .o(n_28293) );
ao22s80 FE_RC_1580_0 ( .a(n_33596), .b(n_33140), .c(n_33141), .d(n_33595), .o(n_33675) );
in01f80 FE_OCP_RBC2812_n_15433 ( .a(FE_OCP_RBN2811_n_15433), .o(FE_OCP_RBN2812_n_15433) );
in01f80 fopt783207 ( .a(FE_OCP_RBN3308_n_44722), .o(n_44759) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_10_ ( .ck(newNet_3264), .d(n_36387), .o(delay_add_ln22_unr23_stage9_stallmux_q_10_) );
in01f80 g762021 ( .a(n_18427), .o(n_18428) );
ao12f80 g780784 ( .a(n_454), .b(n_425), .c(n_365), .o(n_534) );
na02f80 g753584 ( .a(n_27283), .b(n_26898), .o(n_27406) );
in01f80 g749386 ( .a(n_30625), .o(n_30681) );
no02f80 g766205 ( .a(n_14408), .b(n_14270), .o(n_14474) );
in01f80 g773609 ( .a(n_7361), .o(n_7362) );
in01f80 g763425 ( .a(n_17176), .o(n_17177) );
in01f80 newInst_1916 ( .a(newNet_304), .o(newNet_1916) );
no02f80 g747580 ( .a(n_33481), .b(n_33442), .o(n_33498) );
no02f80 g748675 ( .a(n_32537), .b(n_32559), .o(n_32563) );
na02f80 g755115 ( .a(n_25315), .b(n_25318), .o(n_25352) );
in01f80 g768045 ( .a(n_12774), .o(n_12737) );
in01f80 newInst_3337 ( .a(newNet_1812), .o(newNet_3337) );
in01f80 g751827 ( .a(n_28252), .o(n_28253) );
na02f80 g784403 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_25_), .o(n_46215) );
in01f80 fopt783136 ( .a(n_44626), .o(n_44624) );
in01f80 newInst_2710 ( .a(newNet_2655), .o(newNet_2710) );
oa12f80 g749641 ( .a(n_31642), .b(FE_OCP_RBN3708_n_31396), .c(n_31640), .o(n_31690) );
na02f80 g758904 ( .a(n_22061), .b(n_22060), .o(n_22062) );
in01f80 FE_RC_13_0 ( .a(n_1871), .o(FE_RN_3_0) );
in01f80 g758149 ( .a(n_22295), .o(n_22296) );
ao12f80 g747707 ( .a(n_33991), .b(n_33372), .c(n_33743), .o(n_34329) );
in01f80 g760681 ( .a(n_19707), .o(n_19726) );
na02f80 g776118 ( .a(n_5016), .b(n_3663), .o(n_5150) );
na02f80 g760121 ( .a(n_20311), .b(n_20268), .o(n_20312) );
na02f80 g746071 ( .a(n_33853), .b(n_33366), .o(n_33903) );
in01f80 g770502 ( .a(n_10402), .o(n_10403) );
no02f80 g739362 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_20_), .o(n_40785) );
no02f80 g744869 ( .a(n_35032), .b(n_35008), .o(n_35097) );
in01f80 g777162 ( .a(n_5385), .o(n_5386) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_8_ ( .ck(newNet_2699), .d(n_15978), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_8_) );
na02f80 g737426 ( .a(n_42706), .b(n_42495), .o(n_42782) );
na02f80 g741542 ( .a(n_38680), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38721) );
na02f80 FE_RC_2685_0 ( .a(FE_RN_1122_0), .b(n_8580), .o(FE_RN_1123_0) );
no02f80 g759405 ( .a(n_20736), .b(n_20582), .o(n_20801) );
no02f80 g755028 ( .a(n_25743), .b(n_25343), .o(n_25868) );
in01f80 newInst_1754 ( .a(newNet_1753), .o(newNet_1754) );
na02f80 g751325 ( .a(n_29601), .b(n_29074), .o(n_29598) );
in01f80 g749061 ( .a(n_32295), .o(n_32269) );
na02f80 g753586 ( .a(n_26628), .b(n_26590), .o(n_26672) );
no03m80 g748001 ( .a(n_33028), .b(n_33005), .c(n_32488), .o(n_33122) );
no02f80 g775519 ( .a(n_5716), .b(n_4874), .o(n_5711) );
ao12f80 g781164 ( .a(n_77), .b(n_182), .c(n_49), .o(n_183) );
no02f80 g765195 ( .a(n_16021), .b(n_16020), .o(n_16063) );
no02f80 g759545 ( .a(n_20763), .b(n_45013), .o(n_20806) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_29_ ( .ck(newNet_3394), .d(n_27805), .o(delay_add_ln22_unr17_stage7_stallmux_q_29_) );
na02f80 g772957 ( .a(n_8046), .b(n_7999), .o(n_8082) );
na02f80 g759479 ( .a(n_21885), .b(n_21171), .o(n_21699) );
no02f80 g760636 ( .a(n_19780), .b(n_19755), .o(n_19886) );
ao12f80 g765948 ( .a(n_14431), .b(n_15090), .c(n_14430), .o(n_15128) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_20_ ( .ck(newNet_2191), .d(n_1127), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_20_) );
in01f80 g768974 ( .a(n_11772), .o(n_11773) );
na02f80 g753228 ( .a(n_27207), .b(FE_OCP_RBN2853_n_26169), .o(n_27303) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_11_ ( .ck(newNet_2124), .d(n_5748), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_) );
in01f80 FE_OCP_RBC3463_n_7886 ( .a(n_7886), .o(FE_OCP_RBN3463_n_7886) );
no02f80 g736980 ( .a(n_43242), .b(n_43298), .o(n_43356) );
in01f80 g744356 ( .a(n_46224), .o(n_36824) );
no02f80 g779728 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n_1620) );
oa22f80 g749561 ( .a(n_30424), .b(n_30147), .c(n_30425), .d(n_30148), .o(n_30492) );
na02f80 g738379 ( .a(n_41768), .b(n_41564), .o(n_41815) );
na02f80 g756244 ( .a(n_24734), .b(n_24733), .o(n_24735) );
no02f80 g774006 ( .a(n_6907), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_4_), .o(n_6930) );
no02f80 g752159 ( .a(n_28593), .b(n_28055), .o(n_28693) );
in01f80 g751365 ( .a(n_28582), .o(n_28583) );
in01f80 fopt783178 ( .a(n_21164), .o(n_44718) );
na02f80 g768314 ( .a(n_12618), .b(n_12617), .o(n_12638) );
no02f80 g749937 ( .a(n_29893), .b(n_29892), .o(n_29926) );
in01f80 g766840 ( .a(n_13631), .o(n_13632) );
in01f80 g772017 ( .a(n_9692), .o(n_9775) );
ms00f80 cos_out_reg_19_ ( .ck(newNet_3728), .d(n_43844), .o(cos_out_19) );
no02f80 g766879 ( .a(n_14216), .b(FE_OCP_RBN2506_n_13896), .o(n_14491) );
in01f80 FE_OCP_RBC2879_n_15553 ( .a(n_15553), .o(FE_OCP_RBN2879_n_15553) );
in01f80 g764456 ( .a(n_16416), .o(n_16417) );
in01f80 FE_OCP_RBC3222_n_22068 ( .a(FE_OCP_RBN3221_n_22068), .o(FE_OCP_RBN3222_n_22068) );
na02f80 g776360 ( .a(n_4546), .b(n_4625), .o(n_4595) );
no02f80 g755528 ( .a(n_24474), .b(n_24230), .o(n_24581) );
in01f80 newInst_789 ( .a(newNet_788), .o(newNet_789) );
in01f80 g777008 ( .a(n_4006), .o(n_4007) );
na02f80 g769919 ( .a(n_10919), .b(n_44464), .o(n_11000) );
in01f80 newInst_3471 ( .a(newNet_2392), .o(newNet_3471) );
ao22s80 FE_RC_1651_0 ( .a(n_25725), .b(n_26265), .c(n_25724), .d(n_26266), .o(n_26398) );
no02f80 g772569 ( .a(n_8324), .b(n_7927), .o(n_8431) );
in01f80 g760666 ( .a(n_19728), .o(n_19748) );
oa12f80 g755830 ( .a(n_25188), .b(n_25220), .c(n_25124), .o(n_25288) );
in01f80 g774721 ( .a(n_6500), .o(n_6490) );
in01f80 g752353 ( .a(n_27934), .o(n_27935) );
in01f80 g739590 ( .a(n_40643), .o(n_40644) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_15_ ( .ck(newNet_2873), .d(n_11252), .o(delay_add_ln22_unr8_stage4_stallmux_q_15_) );
na02f80 g742254 ( .a(n_44887), .b(n_38268), .o(n_38348) );
no02f80 g740816 ( .a(n_39437), .b(n_39164), .o(n_39532) );
in01f80 g775727 ( .a(n_5658), .o(n_5657) );
in01f80 FE_OCP_RBC3380_n_1732 ( .a(n_1732), .o(FE_OCP_RBN3380_n_1732) );
na02f80 g742395 ( .a(n_37758), .b(n_37777), .o(n_37806) );
ao12f80 g746631 ( .a(n_33990), .b(n_34359), .c(n_33971), .o(n_34420) );
in01f80 newInst_1482 ( .a(newNet_1481), .o(newNet_1482) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_9_ ( .ck(newNet_137), .d(n_46368), .o(delay_xor_ln22_unr9_stage4_stallmux_q_9_) );
in01f80 g756851 ( .a(n_23418), .o(n_23419) );
no02f80 g774188 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_17_), .o(n_7099) );
in01f80 g773799 ( .a(n_7258), .o(n_7241) );
no02f80 g752807 ( .a(n_28259), .b(n_28213), .o(n_28498) );
in01f80 g757766 ( .a(n_22631), .o(n_22611) );
no02f80 FE_RC_1863_0 ( .a(FE_RN_571_0), .b(FE_RN_572_0), .o(n_14201) );
no02f80 g748891 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .o(n_32459) );
in01f80 g775359 ( .a(n_5609), .o(n_5648) );
no02f80 FE_RC_2257_0 ( .a(FE_RN_832_0), .b(FE_RN_833_0), .o(FE_RN_834_0) );
na02f80 g768692 ( .a(n_12183), .b(n_12248), .o(n_12285) );
in01f80 g755649 ( .a(n_24450), .o(n_24469) );
no02f80 g769866 ( .a(n_11085), .b(n_11027), .o(n_11086) );
na02f80 g749544 ( .a(n_30494), .b(n_30493), .o(n_30495) );
in01f80 FE_OCP_RBC2347_n_29448 ( .a(n_29448), .o(FE_OCP_RBN2347_n_29448) );
no02f80 g745409 ( .a(FE_OCP_RBN2986_n_35539), .b(n_35631), .o(n_35634) );
oa12f80 g778193 ( .a(n_2693), .b(n_2692), .c(n_2691), .o(n_4142) );
in01f80 g747432 ( .a(n_32659), .o(n_32660) );
na02f80 g749199 ( .a(FE_OCP_RBN3672_n_30820), .b(n_27131), .o(n_30874) );
in01f80 g758095 ( .a(n_22048), .o(n_22079) );
na02f80 g778961 ( .a(n_2148), .b(n_2120), .o(n_2121) );
no02f80 g773443 ( .a(n_7584), .b(n_6784), .o(n_8846) );
no02f80 g757991 ( .a(n_22127), .b(n_21367), .o(n_22201) );
in01f80 g766043 ( .a(n_15823), .o(n_15085) );
na02f80 g742555 ( .a(n_38298), .b(n_37411), .o(n_37511) );
in01f80 FE_OCP_RBC2752_n_15461 ( .a(n_15461), .o(FE_OCP_RBN2752_n_15461) );
na02f80 g758896 ( .a(n_21435), .b(n_21434), .o(n_21544) );
in01f80 FE_OCPC1462_n_23759 ( .a(FE_OCPN1461_n_23759), .o(FE_OCPN1462_n_23759) );
oa12f80 g747050 ( .a(n_32884), .b(n_32931), .c(n_32846), .o(n_32994) );
in01f80 g752992 ( .a(n_27400), .o(n_27401) );
in01f80 newInst_1427 ( .a(newNet_1426), .o(newNet_1427) );
no02f80 g761141 ( .a(n_19062), .b(n_18392), .o(n_19087) );
in01f80 g739773 ( .a(n_40434), .o(n_40435) );
no02f80 g750454 ( .a(n_29503), .b(FE_OCP_RBN2310_n_29298), .o(n_29552) );
in01f80 g753243 ( .a(n_27214), .o(n_27215) );
in01f80 g774101 ( .a(n_6774), .o(n_6725) );
in01f80 FE_OCP_RBC2768_n_9745 ( .a(n_9745), .o(FE_OCP_RBN2768_n_9745) );
in01f80 newInst_2267 ( .a(newNet_1365), .o(newNet_2267) );
in01f80 g738865 ( .a(n_41296), .o(n_41297) );
in01f80 newInst_2875 ( .a(newNet_2874), .o(newNet_2875) );
na02f80 g760110 ( .a(n_20387), .b(n_19238), .o(n_20436) );
na02f80 g765381 ( .a(FE_OCP_RBN3620_n_15135), .b(n_14056), .o(n_15410) );
in01f80 g744363 ( .a(n_46220), .o(n_36818) );
oa12f80 g761791 ( .a(n_18217), .b(n_18379), .c(n_18377), .o(n_18412) );
oa12f80 g771811 ( .a(n_8963), .b(n_8962), .c(n_8961), .o(n_9065) );
ao22s80 FE_RC_252_0 ( .a(n_19497), .b(FE_OCPN1426_n_18099), .c(n_19645), .d(n_19453), .o(n_19580) );
na02f80 g750548 ( .a(n_30441), .b(n_29910), .o(n_30480) );
no02f80 g769185 ( .a(n_12077), .b(n_12078), .o(n_12119) );
no02f80 g757397 ( .a(n_46964), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_2_), .o(n_23122) );
na02f80 g737025 ( .a(n_43030), .b(n_42780), .o(n_43186) );
no02f80 g776580 ( .a(n_4353), .b(n_4147), .o(n_4448) );
no02f80 g737462 ( .a(n_42639), .b(n_42629), .o(n_42638) );
in01f80 g756187 ( .a(n_24222), .o(n_24245) );
no02f80 g773877 ( .a(n_6997), .b(n_6873), .o(n_7028) );
no02f80 g755437 ( .a(n_24688), .b(FE_OCPN1512_n_22280), .o(n_24759) );
in01f80 newInst_2032 ( .a(newNet_2031), .o(newNet_2032) );
na02f80 g739056 ( .a(n_41090), .b(n_41089), .o(n_41091) );
in01f80 g766297 ( .a(n_14283), .o(n_14254) );
in01f80 g738778 ( .a(n_41382), .o(n_41435) );
na02f80 g754859 ( .a(n_25649), .b(n_25694), .o(n_25724) );
na02f80 g745533 ( .a(FE_OCP_RBN2262_n_33691), .b(n_34509), .o(n_34510) );
oa22f80 g762938 ( .a(n_17678), .b(n_17638), .c(n_17621), .d(n_17637), .o(n_19053) );
oa22f80 g784342 ( .a(FE_OCP_RBN3075_FE_OFN807_n_46195), .b(n_5408), .c(FE_OFN775_n_46137), .d(n_5350), .o(n_46148) );
in01f80 g741478 ( .a(n_38761), .o(n_38762) );
na02f80 g774918 ( .a(n_6144), .b(n_6040), .o(n_6178) );
in01f80 g745103 ( .a(n_34728), .o(n_34727) );
in01f80 g754899 ( .a(n_25301), .o(n_25329) );
in01f80 g763820 ( .a(n_17356), .o(n_17357) );
in01f80 g776246 ( .a(n_4851), .o(n_4911) );
na02f80 g775055 ( .a(n_5979), .b(n_6038), .o(n_6090) );
in01f80 FE_OCP_DRV_C3162_n_21419 ( .a(FE_OCP_DRV_N3161_n_21419), .o(FE_OCP_DRV_N3162_n_21419) );
oa22f80 g748025 ( .a(n_31777), .b(n_31919), .c(n_31748), .d(n_31920), .o(n_31996) );
in01f80 FE_OCP_RBC2440_n_8402 ( .a(FE_OCP_RBN2438_n_8402), .o(FE_OCP_RBN2440_n_8402) );
in01f80 g769066 ( .a(n_11656), .o(n_11716) );
in01f80 FE_OCPC1781_FE_OCP_RBN1701_n_19353 ( .a(FE_OCP_RBN1701_n_19353), .o(FE_OCPN1781_FE_OCP_RBN1701_n_19353) );
no02f80 g771075 ( .a(n_9705), .b(n_8334), .o(n_9928) );
na02f80 g771604 ( .a(n_44055), .b(n_9285), .o(n_9395) );
na02f80 g778579 ( .a(n_2416), .b(n_3317), .o(n_2485) );
na02f80 g748874 ( .a(FE_OCPN1229_n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_14_), .o(n_32420) );
no02f80 g769638 ( .a(n_11205), .b(n_11171), .o(n_11275) );
na02f80 g772331 ( .a(n_8660), .b(n_8561), .o(n_8661) );
no02f80 g739947 ( .a(n_40228), .b(n_40118), .o(n_40229) );
in01f80 g751523 ( .a(n_28847), .o(n_28848) );
na02f80 g770299 ( .a(n_10591), .b(n_10617), .o(n_10709) );
no02f80 g760959 ( .a(n_19225), .b(n_18462), .o(n_19255) );
in01f80 g739971 ( .a(n_40398), .o(n_40367) );
in01f80 FE_OCPC1397_n_21973 ( .a(n_21973), .o(FE_OCPN1397_n_21973) );
in01f80 g752573 ( .a(n_27653), .o(n_27635) );
in01f80 g763152 ( .a(n_17504), .o(n_17505) );
in01f80 FE_OCP_RBC2295_n_2438 ( .a(FE_OCP_RBN2291_n_2438), .o(FE_OCP_RBN2295_n_2438) );
no03m80 g748130 ( .a(n_32796), .b(n_32783), .c(n_32486), .o(n_32865) );
na02f80 g764915 ( .a(n_15440), .b(n_15437), .o(n_15586) );
in01f80 FE_OCP_DRV_C3147_n_33225 ( .a(n_33225), .o(FE_OCP_DRV_N3147_n_33225) );
na02f80 g743816 ( .a(n_37217), .b(n_46231), .o(n_37218) );
oa12f80 g739163 ( .a(n_45155), .b(n_40939), .c(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n_40940) );
in01f80 g744706 ( .a(n_35211), .o(n_35256) );
in01f80 g763652 ( .a(n_18404), .o(n_16931) );
in01f80 newInst_3007 ( .a(newNet_3006), .o(newNet_3007) );
in01f80 g765642 ( .a(n_15041), .o(n_15042) );
oa12f80 g745507 ( .a(n_34943), .b(n_35496), .c(n_34941), .o(n_35543) );
in01f80 g750960 ( .a(n_28965), .o(n_28966) );
na02f80 FE_RC_4032_0 ( .a(FE_RN_1751_0), .b(n_26263), .o(n_26376) );
na02f80 g755450 ( .a(n_24661), .b(n_24698), .o(n_24762) );
na02f80 g767916 ( .a(n_12923), .b(n_12856), .o(n_12924) );
in01f80 FE_OCP_RBC3207_n_44365 ( .a(FE_OCP_RBN3210_n_44365), .o(FE_OCP_RBN3207_n_44365) );
in01f80 g764680 ( .a(n_15987), .o(n_15988) );
in01f80 g752524 ( .a(n_27701), .o(n_27702) );
in01f80 g737473 ( .a(n_43130), .o(n_42666) );
in01f80 g739335 ( .a(n_40693), .o(n_40694) );
na02f80 g779779 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .o(n_1423) );
in01f80 FE_OFC361_n_9391 ( .a(FE_OFN360_n_9391), .o(FE_OFN361_n_9391) );
na02f80 g753872 ( .a(n_26218), .b(n_26253), .o(n_26331) );
na02f80 FE_RC_467_0 ( .a(FE_RN_135_0), .b(FE_RN_136_0), .o(FE_RN_137_0) );
in01f80 g771998 ( .a(n_9772), .o(n_9648) );
in01f80 FE_OCP_RBC2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
ao12f80 g738119 ( .a(n_41885), .b(n_42030), .c(n_41791), .o(n_42043) );
ao12f80 g740841 ( .a(n_38905), .b(n_39399), .c(n_38990), .o(n_39462) );
na02f80 g753884 ( .a(n_27032), .b(n_26887), .o(n_27065) );
in01f80 g759736 ( .a(n_20321), .o(n_20349) );
in01f80 g771031 ( .a(n_10040), .o(n_10041) );
in01f80 newInst_834 ( .a(newNet_127), .o(newNet_834) );
in01f80 g738898 ( .a(n_41310), .o(n_41300) );
no02f80 FE_RC_4234_0 ( .a(n_26003), .b(FE_RN_1859_0), .o(n_26049) );
oa22f80 FE_RC_159_0 ( .a(n_20673), .b(n_20946), .c(n_20672), .d(n_20945), .o(n_21087) );
ao12f80 g749747 ( .a(n_31408), .b(n_31311), .c(n_31372), .o(n_31573) );
in01f80 FE_OCPC3171_n_34222 ( .a(n_34222), .o(FE_OCPN3171_n_34222) );
in01f80 g742192 ( .a(n_38276), .o(n_38277) );
na02f80 g751436 ( .a(n_28762), .b(n_28786), .o(n_28787) );
in01f80 newInst_261 ( .a(newNet_260), .o(newNet_261) );
no02f80 g759040 ( .a(n_21422), .b(n_21277), .o(n_21535) );
no02f80 g748238 ( .a(FE_OCPN880_n_31944), .b(n_30554), .o(n_32098) );
in01f80 newInst_1347 ( .a(newNet_1346), .o(newNet_1347) );
in01f80 g745395 ( .a(n_36050), .o(n_36119) );
in01f80 FE_OCP_RBC3117_n_22710 ( .a(n_22710), .o(FE_OCP_RBN3117_n_22710) );
in01f80 FE_OCPC1042_n_3673 ( .a(FE_OCPN1041_n_3673), .o(FE_OCPN1042_n_3673) );
oa12f80 g737846 ( .a(n_42197), .b(n_42178), .c(n_42196), .o(n_42203) );
in01f80 g763495 ( .a(n_16986), .o(n_17023) );
in01f80 newInst_657 ( .a(newNet_656), .o(newNet_657) );
na02f80 g745972 ( .a(n_33924), .b(n_33963), .o(n_34015) );
na02f80 g763684 ( .a(n_16755), .b(n_16728), .o(n_16787) );
na02f80 FE_RC_4213_0 ( .a(n_19976), .b(n_19804), .o(n_20023) );
in01f80 FE_RC_1322_0 ( .a(n_9909), .o(FE_RN_390_0) );
in01f80 FE_RC_2909_0 ( .a(n_13221), .o(FE_RN_1264_0) );
ao12f80 g774385 ( .a(n_6850), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_), .o(n_7481) );
oa12f80 g779812 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_20_), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n_1714) );
na02f80 g781051 ( .a(cos_out_5), .b(FE_OFN2_n_43918), .o(n_341) );
in01f80 g769792 ( .a(n_11252), .o(n_11220) );
in01f80 g771752 ( .a(n_10239), .o(n_10240) );
in01f80 g745403 ( .a(n_35932), .o(n_35880) );
na02f80 g775609 ( .a(n_5497), .b(n_5504), .o(n_5632) );
in01f80 FE_OCP_RBC1191_n_14911 ( .a(FE_OCP_RBN1189_n_14911), .o(FE_OCP_RBN1191_n_14911) );
ao12f80 g767297 ( .a(n_13550), .b(n_13549), .c(n_13548), .o(n_15342) );
in01f80 g776766 ( .a(n_3993), .o(n_4017) );
ao12f80 g741789 ( .a(n_38332), .b(n_38397), .c(n_38281), .o(n_38427) );
no02f80 FE_RC_1932_0 ( .a(FE_RN_613_0), .b(n_18821), .o(FE_RN_614_0) );
no02f80 g755493 ( .a(n_24780), .b(n_24779), .o(n_24781) );
ao12f80 g765254 ( .a(n_15577), .b(n_15576), .c(n_15575), .o(n_16175) );
in01f80 g738992 ( .a(n_41154), .o(n_41159) );
in01f80 g741911 ( .a(n_38432), .o(n_39181) );
ao12f80 g781222 ( .a(n_110), .b(n_128), .c(n_46055), .o(n_129) );
na02f80 g745176 ( .a(n_34818), .b(n_34782), .o(n_35554) );
no02f80 g766494 ( .a(n_14531), .b(n_14530), .o(n_14532) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_3_ ( .ck(newNet_3197), .d(n_35481), .o(delay_add_ln22_unr23_stage9_stallmux_q_3_) );
ao12f80 g750622 ( .a(FE_RN_1513_0), .b(n_29272), .c(n_29160), .o(n_29407) );
na02f80 g772400 ( .a(n_8525), .b(FE_OCP_RBN3465_n_7886), .o(n_8603) );
ao12f80 g747967 ( .a(n_31848), .b(n_32060), .c(n_32139), .o(n_32186) );
ao12f80 g760472 ( .a(n_20514), .b(n_20513), .c(n_20512), .o(n_21371) );
na02f80 g761265 ( .a(n_19934), .b(n_19905), .o(n_19935) );
na02f80 g776807 ( .a(n_4168), .b(n_2583), .o(n_4275) );
na02f80 g777630 ( .a(n_3334), .b(n_3200), .o(n_3416) );
no02f80 g768788 ( .a(n_12095), .b(n_12094), .o(n_12096) );
in01f80 g758844 ( .a(n_21552), .o(n_21553) );
no02f80 g776420 ( .a(n_4343), .b(n_4093), .o(n_4403) );
no02f80 g742451 ( .a(n_37648), .b(n_37666), .o(n_37742) );
in01f80 FE_OCP_RBC3541_n_34487 ( .a(n_34487), .o(FE_OCP_RBN3541_n_34487) );
ao22s80 g761808 ( .a(FE_OCP_RBN1155_n_18375), .b(n_16968), .c(FE_OCP_RBN1157_n_18375), .d(n_18483), .o(n_18642) );
in01f80 newInst_3306 ( .a(newNet_3305), .o(newNet_3306) );
na02f80 g775498 ( .a(n_5716), .b(n_5665), .o(n_5666) );
no02f80 g753449 ( .a(n_26960), .b(n_26876), .o(n_26983) );
na02f80 g776856 ( .a(n_3968), .b(FE_OCP_RBN2486_n_3498), .o(n_4155) );
no02f80 g762822 ( .a(n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .o(n_17758) );
no02f80 g750507 ( .a(n_29481), .b(n_29400), .o(n_29483) );
na02f80 g771018 ( .a(n_9989), .b(n_9988), .o(n_10027) );
in01f80 g779384 ( .a(n_1541), .o(n_1589) );
na02f80 g750651 ( .a(n_29437), .b(n_29436), .o(n_29438) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_1_ ( .ck(newNet_1520), .d(n_31226), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_1_) );
in01f80 newInst_2176 ( .a(newNet_2115), .o(newNet_2176) );
in01f80 newInst_3410 ( .a(newNet_3409), .o(newNet_3410) );
oa12f80 g784664 ( .a(n_6224), .b(n_6178), .c(n_6119), .o(n_46994) );
no02f80 g776975 ( .a(n_3774), .b(n_3846), .o(n_3948) );
oa12f80 g749009 ( .a(n_31124), .b(n_31123), .c(n_31122), .o(n_31176) );
na02f80 g741242 ( .a(n_38847), .b(n_38509), .o(n_39060) );
in01f80 newInst_103 ( .a(newNet_102), .o(newNet_103) );
oa12f80 g767233 ( .a(n_13252), .b(n_13696), .c(n_13249), .o(n_13770) );
na02f80 FE_RC_2407_0 ( .a(n_6540), .b(n_6569), .o(FE_RN_948_0) );
no02f80 g769968 ( .a(n_10883), .b(n_10859), .o(n_10896) );
no02f80 g771864 ( .a(n_9432), .b(n_9547), .o(n_10217) );
ao12f80 g769190 ( .a(FE_OCP_RBN1927_cordic_combinational_sub_ln23_0_unr12_z_0__), .b(FE_OCP_RBN1991_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .c(n_45224), .o(n_11537) );
in01f80 g770630 ( .a(n_10422), .o(n_10527) );
no02f80 g770612 ( .a(FE_OCP_RBN2830_n_10198), .b(FE_OCP_RBN3594_n_44561), .o(n_10267) );
na02f80 g736362 ( .a(n_43789), .b(n_43291), .o(n_43811) );
no02f80 g765186 ( .a(n_15079), .b(FE_OCPN1007_n_13962), .o(n_15123) );
na02f80 g740937 ( .a(n_39254), .b(n_39253), .o(n_39255) );
na02f80 g763062 ( .a(n_17620), .b(delay_add_ln22_unr11_stage5_stallmux_q_5_), .o(n_17715) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_24_ ( .ck(newNet_3136), .d(n_40549), .o(delay_add_ln22_unr27_stage10_stallmux_q_24_) );
no02f80 FE_RC_2782_0 ( .a(FE_RN_1187_0), .b(FE_OCPN1426_n_18099), .o(n_19784) );
ao22s80 g750026 ( .a(n_29869), .b(n_29083), .c(n_29896), .d(n_29113), .o(n_30447) );
na02f80 g748804 ( .a(n_32450), .b(n_32318), .o(n_32451) );
in01f80 g762326 ( .a(n_18198), .o(n_18199) );
na02f80 g739317 ( .a(n_40673), .b(n_40735), .o(n_40799) );
in01f80 g737850 ( .a(n_42693), .o(n_42694) );
in01f80 g776541 ( .a(n_4378), .o(n_4379) );
oa22f80 FE_RC_975_0 ( .a(n_32243), .b(n_31796), .c(n_32225), .d(n_31797), .o(n_32339) );
ao12f80 g750578 ( .a(n_29515), .b(n_29514), .c(n_29513), .o(n_30917) );
na02f80 g763607 ( .a(n_16809), .b(n_16761), .o(n_16833) );
in01f80 newInst_1212 ( .a(newNet_1211), .o(newNet_1212) );
ao22s80 g769311 ( .a(n_12164), .b(FE_OCPN1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .c(n_11707), .d(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_), .o(n_12356) );
na02f80 g756494 ( .a(n_23762), .b(n_23761), .o(n_23788) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_15_ ( .ck(newNet_3069), .d(n_1188), .o(delay_add_ln22_unr2_stage2_stallmux_q_15_) );
in01f80 g775204 ( .a(n_5962), .o(n_5963) );
ao12f80 g741222 ( .a(n_38903), .b(FE_OCP_RBN2550_n_44944), .c(n_38953), .o(n_39322) );
in01f80 newInst_2314 ( .a(newNet_2313), .o(newNet_2314) );
oa22f80 g784545 ( .a(n_11494), .b(FE_OFN801_n_46285), .c(n_11463), .d(FE_OCP_RBN3044_n_46337), .o(n_46366) );
na02f80 g736816 ( .a(FE_OCP_RBN3096_n_43489), .b(n_43553), .o(n_43621) );
in01f80 newInst_889 ( .a(newNet_888), .o(newNet_889) );
no02f80 g737054 ( .a(n_43171), .b(n_43170), .o(n_43202) );
no02f80 g756795 ( .a(n_23460), .b(n_23097), .o(n_23440) );
no02f80 g776741 ( .a(n_4110), .b(n_4164), .o(n_4340) );
na02f80 g762271 ( .a(n_18622), .b(n_18614), .o(n_18845) );
in01f80 FE_OCP_RBC2419_n_19601 ( .a(n_19601), .o(FE_OCP_RBN2419_n_19601) );
na02f80 g781338 ( .a(n_51), .b(n_46055), .o(n_91) );
in01f80 g776645 ( .a(n_4492), .o(n_4493) );
no02f80 FE_RC_1660_0 ( .a(n_37709), .b(n_37559), .o(FE_RN_462_0) );
na02f80 g771284 ( .a(FE_OCP_RBN2660_n_9292), .b(FE_OCP_RBN3555_n_44575), .o(n_9371) );
in01f80 FE_OCP_RBC2266_n_2430 ( .a(n_2430), .o(FE_OCP_RBN2266_n_2430) );
na02f80 g749261 ( .a(n_30792), .b(n_27130), .o(n_30845) );
no02f80 FE_RC_2733_0 ( .a(FE_RN_1156_0), .b(FE_RN_1157_0), .o(FE_RN_1158_0) );
oa12f80 g746525 ( .a(n_34417), .b(n_34475), .c(n_35542), .o(n_34529) );
ao22s80 FE_RC_3460_0 ( .a(n_31014), .b(FE_RN_729_0), .c(n_30937), .d(FE_RN_730_0), .o(n_31165) );
in01f80 FE_OCP_RBC3214_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3214_n_44365) );
in01f80 newInst_2775 ( .a(newNet_2774), .o(newNet_2775) );
na04m80 FE_RC_1524_0 ( .a(n_44962), .b(FE_OCPN1236_n_32791), .c(n_32721), .d(n_32790), .o(n_32795) );
in01f80 g747459 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .o(n_32613) );
no02f80 g742250 ( .a(n_44887), .b(n_37334), .o(n_38254) );
na02f80 g777809 ( .a(n_4336), .b(n_2759), .o(n_3257) );
no02f80 g770886 ( .a(FE_OCP_RBN2770_n_9892), .b(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .o(n_9967) );
in01f80 fopt782910 ( .a(n_32169), .o(n_44358) );
in01f80 g743591 ( .a(n_36529), .o(n_36530) );
oa12f80 g754832 ( .a(n_25254), .b(n_25923), .c(n_25189), .o(n_25952) );
in01f80 g766301 ( .a(n_14439), .o(n_14821) );
na02f80 g764785 ( .a(n_15730), .b(n_15695), .o(n_15795) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_14_ ( .ck(newNet_2019), .d(n_11212), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_) );
no02f80 g740175 ( .a(FE_OCP_RBN3056_n_39913), .b(n_39947), .o(n_40116) );
na02f80 FE_RC_1951_0 ( .a(n_24438), .b(n_25786), .o(FE_RN_627_0) );
no02f80 g758088 ( .a(FE_OCPN3166_n_44267), .b(FE_OCP_RBN1371_n_20763), .o(n_22345) );
no02f80 g760050 ( .a(n_20577), .b(FE_OCPN1261_n_20242), .o(n_20631) );
in01f80 g760797 ( .a(n_19637), .o(n_19621) );
no02f80 g776904 ( .a(n_3955), .b(FE_OCP_RBN3575_n_4528), .o(n_3901) );
in01f80 g784794 ( .a(n_47334), .o(n_47335) );
in01f80 g744749 ( .a(n_35121), .o(n_35348) );
na02f80 g766363 ( .a(n_14163), .b(n_13322), .o(n_14194) );
in01f80 g740428 ( .a(n_39829), .o(n_39830) );
in01f80 FE_OCP_RBC1141_n_25816 ( .a(n_25816), .o(FE_OCP_RBN1141_n_25816) );
oa12f80 g783828 ( .a(n_45841), .b(n_39596), .c(n_39607), .o(n_45514) );
in01f80 g764015 ( .a(n_19418), .o(n_18119) );
in01f80 g777033 ( .a(n_3814), .o(n_3845) );
in01f80 newInst_449 ( .a(newNet_448), .o(newNet_449) );
na02f80 g738594 ( .a(n_41445), .b(n_41444), .o(n_41446) );
in01f80 g767726 ( .a(n_13206), .o(n_13207) );
in01f80 g770602 ( .a(n_10411), .o(n_10394) );
no02f80 FE_RC_2890_0 ( .a(FE_RN_1251_0), .b(n_24870), .o(n_24918) );
in01f80 g754171 ( .a(n_26048), .o(n_26110) );
na02f80 g761331 ( .a(n_19709), .b(n_19652), .o(n_19764) );
in01f80 g748789 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_2_), .o(n_32654) );
na02f80 g777059 ( .a(n_3720), .b(n_3029), .o(n_3753) );
in01f80 newInst_3461 ( .a(newNet_3460), .o(newNet_3461) );
in01f80 FE_OCPC991_n_22249 ( .a(FE_OCPN990_n_22249), .o(FE_OCPN991_n_22249) );
in01f80 g776695 ( .a(n_4220), .o(n_4221) );
in01f80 g764122 ( .a(n_16928), .o(n_16929) );
in01f80 FE_RC_676_0 ( .a(n_17582), .o(FE_RN_217_0) );
in01f80 g757876 ( .a(n_22392), .o(n_22355) );
na02f80 g767968 ( .a(n_13248), .b(n_13161), .o(n_13274) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_10_ ( .ck(newNet_470), .d(n_27780), .o(delay_xor_ln22_unr18_stage7_stallmux_q_10_) );
in01f80 g739381 ( .a(n_40892), .o(n_40840) );
no02f80 g751880 ( .a(n_28859), .b(n_29200), .o(n_28926) );
na02f80 g741735 ( .a(n_38476), .b(n_38497), .o(n_38545) );
in01f80 newInst_1052 ( .a(newNet_458), .o(newNet_1052) );
in01f80 g739122 ( .a(n_41060), .o(n_41046) );
ms00f80 mux_while_ln12_psv_q_reg_3_ ( .ck(newNet_116), .d(n_181), .o(mux_while_ln12_psv_q_3_) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_31_ ( .ck(newNet_2252), .d(n_40579), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_31_) );
in01f80 newInst_2809 ( .a(newNet_2808), .o(newNet_2809) );
in01f80 g737688 ( .a(n_42395), .o(n_42396) );
na02f80 g738265 ( .a(n_41894), .b(n_41893), .o(n_41895) );
no02f80 g770187 ( .a(n_10784), .b(FE_OCP_RBN2677_n_9247), .o(n_10871) );
in01f80 newInst_2384 ( .a(newNet_2383), .o(newNet_2384) );
na02f80 g770933 ( .a(n_9806), .b(n_9624), .o(n_9853) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_23_ ( .ck(newNet_3614), .d(n_17630), .o(delay_add_ln22_unr11_stage5_stallmux_q_23_) );
no02f80 g781198 ( .a(n_168), .b(n_264), .o(n_173) );
ao12f80 g779481 ( .a(n_1945), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_20_), .o(n_1996) );
in01f80 FE_RC_3206_0 ( .a(n_1102), .o(FE_RN_1425_0) );
na02f80 g740745 ( .a(n_39412), .b(n_39444), .o(n_39969) );
in01f80 g776813 ( .a(n_4075), .o(n_4213) );
na02f80 g764153 ( .a(n_16499), .b(n_46421), .o(n_16518) );
in01f80 g750288 ( .a(n_29753), .o(n_29754) );
oa12f80 g763516 ( .a(n_17541), .b(n_17424), .c(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17542) );
na02f80 g772721 ( .a(FE_OCP_RBN3498_n_8187), .b(n_7743), .o(n_8217) );
na03f80 g747394 ( .a(n_33579), .b(n_33533), .c(n_33417), .o(n_33863) );
in01f80 g769628 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_), .o(n_12672) );
na02f80 g776706 ( .a(n_4186), .b(n_4116), .o(n_4245) );
no02f80 g763609 ( .a(n_16791), .b(FE_OCP_RBN2761_n_15200), .o(n_16808) );
in01f80 FE_OCP_RBC3553_n_44575 ( .a(FE_OCP_RBN3546_n_44575), .o(FE_OCP_RBN3553_n_44575) );
in01f80 FE_OCP_DRV_C1558_n_19590 ( .a(FE_OCP_DRV_N1557_n_19590), .o(FE_OCP_DRV_N1558_n_19590) );
in01f80 g769393 ( .a(n_11473), .o(n_11474) );
in01f80 g736652 ( .a(n_43565), .o(n_43525) );
in01f80 newInst_25 ( .a(newNet_24), .o(newNet_25) );
no02f80 g775898 ( .a(n_5011), .b(n_4902), .o(n_5121) );
no02f80 g778435 ( .a(n_2479), .b(n_2378), .o(n_2480) );
na02f80 g773754 ( .a(n_7232), .b(n_7219), .o(n_7272) );
na02f80 g756574 ( .a(n_23581), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_17_), .o(n_23583) );
in01f80 g764994 ( .a(n_15468), .o(n_15469) );
in01f80 g757595 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_25_), .o(n_22858) );
in01f80 g776085 ( .a(FE_OCP_RBN2820_n_4872), .o(n_4900) );
no02f80 g762018 ( .a(n_18462), .b(n_18461), .o(n_18463) );
na02f80 g770413 ( .a(n_10483), .b(n_44490), .o(n_10535) );
in01f80 g766945 ( .a(n_13869), .o(n_13870) );
oa12f80 g778358 ( .a(n_2447), .b(n_2446), .c(n_2445), .o(n_2531) );
no02f80 g775336 ( .a(n_5700), .b(n_4875), .o(n_5808) );
no02f80 g747870 ( .a(n_33172), .b(n_33171), .o(n_33173) );
ao12f80 g756357 ( .a(n_24416), .b(n_24415), .c(n_24414), .o(n_25090) );
no02f80 g748106 ( .a(n_32809), .b(n_32421), .o(n_32843) );
oa12f80 g776827 ( .a(n_3568), .b(n_3630), .c(n_3535), .o(n_3786) );
in01f80 g744784 ( .a(n_35177), .o(n_35227) );
no02f80 g772850 ( .a(n_7976), .b(n_7975), .o(n_7977) );
oa12f80 g753845 ( .a(n_26508), .b(n_27035), .c(n_26549), .o(n_27079) );
in01f80 g770721 ( .a(n_10456), .o(n_10457) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_3_ ( .ck(newNet_1288), .d(n_738), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_) );
in01f80 newInst_3590 ( .a(newNet_3589), .o(newNet_3590) );
in01f80 FE_OCP_RBC3002_n_10805 ( .a(n_10805), .o(FE_OCP_RBN3002_n_10805) );
na02f80 g736707 ( .a(n_43269), .b(FE_OCPN912_n_43022), .o(n_43365) );
no02f80 FE_RC_3818_0 ( .a(FE_RN_1664_0), .b(FE_RN_1665_0), .o(FE_RN_1666_0) );
no02f80 g773232 ( .a(n_7669), .b(n_7737), .o(n_7738) );
na02f80 g772919 ( .a(n_7749), .b(n_7366), .o(n_7791) );
in01f80 g748209 ( .a(n_32120), .o(n_32121) );
no02f80 FE_RC_1842_0 ( .a(n_35751), .b(n_35667), .o(FE_RN_558_0) );
oa22f80 FE_RC_246_0 ( .a(n_13626), .b(n_13607), .c(n_13617), .d(n_13625), .o(n_13683) );
in01f80 g768522 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_17_), .o(n_12360) );
in01f80 g766348 ( .a(n_14197), .o(n_14198) );
in01f80 g780573 ( .a(n_1015), .o(n_1016) );
in01f80 g751180 ( .a(n_30028), .o(n_30090) );
oa12f80 g741954 ( .a(n_37988), .b(n_44036), .c(n_37987), .o(n_38060) );
oa12f80 g773483 ( .a(n_6944), .b(n_7525), .c(n_6756), .o(n_7538) );
in01f80 g761587 ( .a(n_20231), .o(n_20252) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_30_ ( .ck(newNet_2528), .d(n_27783), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_) );
na02f80 g775200 ( .a(n_5895), .b(n_5621), .o(n_5914) );
no02f80 g743514 ( .a(n_37673), .b(n_37672), .o(n_37674) );
no02f80 g739991 ( .a(n_40120), .b(n_40081), .o(n_40156) );
in01f80 g743162 ( .a(n_37029), .o(n_36982) );
in01f80 g749971 ( .a(n_30220), .o(n_30221) );
no02f80 g766822 ( .a(n_14343), .b(n_14426), .o(n_14429) );
na02f80 g780291 ( .a(n_833), .b(n_881), .o(n_970) );
na02f80 g762141 ( .a(n_18817), .b(n_18816), .o(n_18932) );
no02f80 g772606 ( .a(n_8392), .b(n_8293), .o(n_8421) );
in01f80 g740123 ( .a(n_40318), .o(n_40319) );
na02f80 g745388 ( .a(FE_OCP_RBN2987_n_35539), .b(n_36019), .o(n_36121) );
in01f80 g739358 ( .a(n_40908), .o(n_40842) );
na02f80 g757658 ( .a(FE_OCP_RBN1194_n_22542), .b(n_22231), .o(n_22584) );
na02f80 g764401 ( .a(n_16655), .b(n_16674), .o(n_16721) );
in01f80 g737190 ( .a(n_43388), .o(n_43005) );
in01f80 FE_RC_1353_0 ( .a(n_30403), .o(FE_RN_402_0) );
in01f80 newInst_3254 ( .a(newNet_201), .o(newNet_3254) );
no02f80 g748084 ( .a(n_31907), .b(n_31953), .o(n_31971) );
in01f80 g768907 ( .a(n_12747), .o(n_11943) );
na02f80 g779388 ( .a(n_1782), .b(n_1746), .o(n_1840) );
na02f80 g760364 ( .a(n_20169), .b(n_20123), .o(n_20192) );
in01f80 g762374 ( .a(n_18737), .o(n_18611) );
in01f80 g745292 ( .a(n_35935), .o(n_35936) );
oa22f80 g763212 ( .a(n_46974), .b(n_17336), .c(n_17003), .d(n_16338), .o(n_17144) );
in01f80 FE_OCPC1490_n_30823 ( .a(FE_OCPN1489_n_30823), .o(FE_OCPN1490_n_30823) );
na02f80 g770501 ( .a(n_10411), .b(n_44464), .o(n_10503) );
in01f80 newInst_1902 ( .a(newNet_1721), .o(newNet_1902) );
na02f80 g764420 ( .a(n_16169), .b(n_14420), .o(n_16170) );
oa12f80 g741976 ( .a(n_37919), .b(n_37918), .c(n_37917), .o(n_38791) );
oa12f80 g757918 ( .a(n_22012), .b(n_22106), .c(n_21982), .o(n_22168) );
in01f80 newInst_2836 ( .a(newNet_2835), .o(newNet_2836) );
in01f80 g772537 ( .a(n_8386), .o(n_8387) );
in01f80 newInst_904 ( .a(newNet_582), .o(newNet_904) );
in01f80 newInst_2348 ( .a(newNet_736), .o(newNet_2348) );
in01f80 g766105 ( .a(n_14607), .o(n_14608) );
no02f80 g762685 ( .a(FE_OCP_RBN2140_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_11_), .o(n_17851) );
in01f80 g769617 ( .a(n_11327), .o(n_11328) );
ao12f80 g738757 ( .a(FE_OCPN1013_n_41478), .b(n_41526), .c(n_41123), .o(n_41692) );
no02f80 g755829 ( .a(n_25087), .b(n_25032), .o(n_25142) );
na02f80 g780582 ( .a(n_923), .b(n_633), .o(n_1052) );
ao22s80 g780250 ( .a(n_980), .b(n_1099), .c(n_979), .d(n_1098), .o(n_1106) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_19_ ( .ck(newNet_1322), .d(n_1241), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_) );
ao12f80 g750409 ( .a(n_29525), .b(n_29570), .c(n_29606), .o(n_29666) );
in01f80 g771718 ( .a(n_8842), .o(n_8865) );
no02f80 g769004 ( .a(n_11844), .b(n_11691), .o(n_11829) );
no02f80 g779574 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_21_), .o(n_1971) );
na02f80 g737036 ( .a(n_43032), .b(n_43031), .o(n_43048) );
no02f80 g777909 ( .a(n_3183), .b(n_3122), .o(n_3196) );
na02f80 g775512 ( .a(n_5419), .b(n_5443), .o(n_5505) );
in01f80 g746514 ( .a(n_34812), .o(n_34865) );
ao22s80 g779499 ( .a(n_1370), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(n_1358), .d(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .o(n_1448) );
ao22s80 g780394 ( .a(n_847), .b(n_1098), .c(n_815), .d(n_1099), .o(n_875) );
no02f80 g773596 ( .a(n_45865), .b(n_6943), .o(n_7434) );
in01f80 FE_OCP_RBC2416_n_8293 ( .a(n_8293), .o(FE_OCP_RBN2416_n_8293) );
oa12f80 g775743 ( .a(n_5052), .b(n_5367), .c(n_4980), .o(n_5455) );
in01f80 g762185 ( .a(n_18193), .o(n_18217) );
in01f80 g753231 ( .a(n_27336), .o(n_27337) );
no02f80 g767935 ( .a(n_12741), .b(n_12740), .o(n_12742) );
ao22s80 g779520 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(n_1371), .c(FE_OCP_RBN3242_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .d(delay_xor_ln22_unr3_stage2_stallmux_q_0_), .o(n_1941) );
in01f80 g776500 ( .a(n_4544), .o(n_4688) );
oa12f80 g765226 ( .a(n_15719), .b(n_15787), .c(n_15786), .o(n_15836) );
na02f80 g756279 ( .a(n_24079), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24121) );
no02f80 g774481 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_21_), .o(n_6863) );
in01f80 g763874 ( .a(n_17526), .o(n_17527) );
na02f80 g771526 ( .a(n_9396), .b(n_9388), .o(n_9484) );
na02f80 g740978 ( .a(n_39253), .b(n_39233), .o(n_39280) );
in01f80 g751395 ( .a(n_29388), .o(n_29358) );
in01f80 g751705 ( .a(n_28387), .o(n_28388) );
in01f80 newInst_120 ( .a(newNet_119), .o(newNet_120) );
in01f80 g746199 ( .a(n_33675), .o(n_33691) );
in01f80 fopt783916 ( .a(n_7594), .o(n_45616) );
ms00f80 sin_out_reg_30_ ( .ck(newNet_31), .d(n_43919), .o(sin_out_30) );
oa12f80 g759212 ( .a(n_21892), .b(n_21891), .c(n_21890), .o(n_21933) );
no02f80 g762005 ( .a(n_18227), .b(n_18204), .o(n_18302) );
na02f80 g769972 ( .a(n_10886), .b(n_10894), .o(n_10965) );
in01f80 g779763 ( .a(n_1619), .o(n_1584) );
no02f80 g759761 ( .a(n_21407), .b(n_21378), .o(n_21408) );
in01f80 g768835 ( .a(n_12019), .o(n_12020) );
no02f80 g748233 ( .a(FE_OCP_RBN3734_n_31819), .b(n_31770), .o(n_32103) );
ao12f80 g750152 ( .a(n_30096), .b(n_30923), .c(n_30431), .o(n_30973) );
na02f80 g744809 ( .a(n_36464), .b(n_35941), .o(n_36479) );
in01f80 newInst_1444 ( .a(newNet_1443), .o(newNet_1444) );
in01f80 newInst_2156 ( .a(newNet_2155), .o(newNet_2156) );
no02f80 g771262 ( .a(n_9313), .b(n_8232), .o(n_9552) );
no02f80 g740681 ( .a(n_39551), .b(n_45840), .o(n_39569) );
in01f80 g747351 ( .a(n_32638), .o(n_32616) );
in01f80 g753097 ( .a(n_27398), .o(n_27399) );
oa12f80 g754986 ( .a(n_25801), .b(n_25800), .c(n_25799), .o(n_26544) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_1_ ( .ck(newNet_1408), .d(n_35726), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_) );
in01f80 g746280 ( .a(n_33549), .o(n_33568) );
in01f80 g762301 ( .a(n_18161), .o(n_18162) );
in01f80 FE_OCP_RBC2522_n_8951 ( .a(n_8951), .o(FE_OCP_RBN2522_n_8951) );
in01f80 g775572 ( .a(n_5849), .o(n_5850) );
in01f80 g759955 ( .a(n_20271), .o(n_20272) );
na02f80 FE_RC_2362_0 ( .a(FE_RN_911_0), .b(FE_RN_913_0), .o(n_19339) );
ao12f80 g740949 ( .a(n_38865), .b(n_38934), .c(n_38897), .o(n_39088) );
na03f80 FE_RC_660_0 ( .a(n_37754), .b(n_37755), .c(n_37756), .o(n_37780) );
na02f80 g773771 ( .a(n_7203), .b(n_7040), .o(n_7232) );
in01f80 g751745 ( .a(n_29078), .o(n_29132) );
no02f80 g776313 ( .a(n_4552), .b(n_3951), .o(n_4616) );
in01f80 g775451 ( .a(n_5540), .o(n_5541) );
ao12f80 g768801 ( .a(n_12147), .b(n_45685), .c(delay_xor_ln21_unr9_stage4_stallmux_q_13_), .o(n_12477) );
in01f80 g743807 ( .a(n_36324), .o(n_36073) );
na02f80 g756197 ( .a(n_24742), .b(n_24090), .o(n_24791) );
na02f80 g747184 ( .a(n_32827), .b(delay_add_ln22_unr20_stage8_stallmux_q_5_), .o(n_32867) );
no02f80 g770359 ( .a(n_10567), .b(n_10586), .o(n_10597) );
in01f80 g776982 ( .a(n_3966), .o(n_3967) );
no02f80 g754687 ( .a(n_26231), .b(n_26310), .o(n_26385) );
oa12f80 g746105 ( .a(n_33822), .b(n_33868), .c(n_33821), .o(n_33940) );
in01f80 g777993 ( .a(n_3154), .o(n_3199) );
in01f80 g776949 ( .a(n_3630), .o(n_3656) );
in01f80 FE_OCP_RBC2280_n_24199 ( .a(n_24199), .o(FE_OCP_RBN2280_n_24199) );
na02f80 g750880 ( .a(n_28979), .b(n_28598), .o(n_29039) );
na02f80 g750303 ( .a(n_29674), .b(n_29589), .o(n_29736) );
na02f80 g764179 ( .a(n_16529), .b(n_16406), .o(n_16596) );
in01f80 FE_OCP_RBC3681_n_26171 ( .a(n_26171), .o(FE_OCP_RBN3681_n_26171) );
in01f80 g781354 ( .a(beta_10), .o(n_38) );
no02f80 g763570 ( .a(n_16717), .b(n_16764), .o(n_16836) );
ao12f80 g746452 ( .a(n_33401), .b(n_33453), .c(n_33036), .o(n_33456) );
na02f80 g738555 ( .a(n_41500), .b(n_41483), .o(n_41573) );
in01f80 g742768 ( .a(n_37350), .o(n_37337) );
in01f80 FE_OCP_RBC2277_n_24173 ( .a(n_24173), .o(FE_OCP_RBN2277_n_24173) );
no02f80 g771402 ( .a(n_9563), .b(n_9687), .o(n_9564) );
no02f80 g742917 ( .a(n_37071), .b(n_37070), .o(n_37428) );
ao12f80 g752751 ( .a(n_27548), .b(FE_OCPN964_n_27287), .c(n_27510), .o(n_27561) );
no02f80 g776052 ( .a(n_5224), .b(n_5146), .o(n_5225) );
in01f80 newInst_1623 ( .a(newNet_1622), .o(newNet_1623) );
in01f80 g767740 ( .a(n_13130), .o(n_13131) );
in01f80 g738965 ( .a(n_41213), .o(n_41214) );
in01f80 g749091 ( .a(n_30961), .o(n_30962) );
no02f80 g761556 ( .a(n_18939), .b(n_17644), .o(n_19022) );
no02f80 g777752 ( .a(n_3316), .b(n_3298), .o(n_4228) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_3_ ( .ck(newNet_3283), .d(n_31110), .o(delay_add_ln22_unr20_stage8_stallmux_q_3_) );
in01f80 g748343 ( .a(n_31831), .o(n_31832) );
na02f80 g765324 ( .a(FE_OCP_RBN2433_n_14018), .b(n_15135), .o(n_15302) );
no02f80 g741690 ( .a(n_38530), .b(n_38778), .o(n_38551) );
in01f80 fopt783662 ( .a(n_27782), .o(n_45309) );
no02f80 g761459 ( .a(n_19609), .b(n_19608), .o(n_19651) );
no02f80 g774062 ( .a(n_6777), .b(n_6790), .o(n_6907) );
na02f80 g771195 ( .a(n_9489), .b(FE_OCP_RBN3588_n_9408), .o(n_9572) );
ao22s80 FE_RC_2623_0 ( .a(n_14417), .b(n_14514), .c(FE_OCPN1055_n_14098), .d(n_14418), .o(n_14585) );
na02f80 g743122 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .o(n_37042) );
in01f80 newInst_1933 ( .a(newNet_1932), .o(newNet_1933) );
no02f80 g764691 ( .a(n_15772), .b(n_15771), .o(n_15773) );
in01f80 g764845 ( .a(FE_OCP_RBN2779_n_15595), .o(n_15651) );
in01f80 g759651 ( .a(n_20641), .o(n_20642) );
in01f80 g744086 ( .a(n_35650), .o(n_35621) );
in01f80 g743565 ( .a(n_37613), .o(n_37614) );
in01f80 newInst_3249 ( .a(newNet_1216), .o(newNet_3249) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_5_ ( .ck(newNet_149), .d(n_46370), .o(delay_xor_ln22_unr9_stage4_stallmux_q_5_) );
in01f80 newInst_2864 ( .a(newNet_2863), .o(newNet_2864) );
na02f80 g771194 ( .a(n_9495), .b(n_9351), .o(n_9553) );
in01f80 g759959 ( .a(n_20501), .o(n_20502) );
in01f80 fopt782977 ( .a(n_24992), .o(n_44445) );
in01f80 FE_RC_3582_0 ( .a(n_14224), .o(FE_RN_1561_0) );
na02f80 g763604 ( .a(n_16731), .b(n_16736), .o(n_16763) );
in01f80 g743840 ( .a(n_37168), .o(n_37169) );
in01f80 newInst_1472 ( .a(newNet_843), .o(newNet_1472) );
in01f80 newInst_785 ( .a(newNet_784), .o(newNet_785) );
in01f80 g762184 ( .a(n_18217), .o(n_18200) );
in01f80 g780588 ( .a(n_677), .o(n_706) );
no02f80 g773620 ( .a(n_7345), .b(n_7344), .o(n_7349) );
no02f80 g742064 ( .a(n_37973), .b(n_37974), .o(n_38008) );
in01f80 g763227 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_18_), .o(n_17050) );
ao12f80 g755303 ( .a(n_24788), .b(n_24787), .c(n_24660), .o(n_24898) );
no02f80 g775115 ( .a(n_5734), .b(n_5760), .o(n_5893) );
in01f80 g780374 ( .a(n_903), .o(n_922) );
in01f80 newInst_667 ( .a(newNet_666), .o(newNet_667) );
na02f80 g742956 ( .a(n_37174), .b(n_37084), .o(n_37203) );
in01f80 newInst_1368 ( .a(newNet_1367), .o(newNet_1368) );
no02f80 g762143 ( .a(n_18814), .b(n_18577), .o(n_18815) );
in01f80 g753140 ( .a(n_27459), .o(n_27460) );
no02f80 g746618 ( .a(n_34473), .b(n_34472), .o(n_34496) );
no02f80 g767358 ( .a(n_13480), .b(n_13548), .o(n_13481) );
na02f80 g738375 ( .a(n_41630), .b(FE_OCP_RBN2312_n_41420), .o(n_41753) );
in01f80 newInst_2067 ( .a(newNet_2066), .o(newNet_2067) );
in01f80 FE_OCP_RBC3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
no02f80 g742809 ( .a(n_37233), .b(n_37083), .o(n_37258) );
in01f80 g749727 ( .a(n_31537), .o(n_31538) );
ao12f80 g755631 ( .a(n_23850), .b(n_24463), .c(FE_OCPN1476_n_23708), .o(n_24562) );
na02f80 g742741 ( .a(n_37353), .b(n_37366), .o(n_37395) );
ao12f80 g740771 ( .a(n_39313), .b(n_39314), .c(n_39010), .o(n_39414) );
no02f80 g748134 ( .a(n_32769), .b(n_32796), .o(n_32824) );
no03m80 g766083 ( .a(n_14947), .b(n_14948), .c(n_14338), .o(n_15030) );
in01f80 FE_OCP_RBC2681_n_15048 ( .a(n_15048), .o(FE_OCP_RBN2681_n_15048) );
oa12f80 g751419 ( .a(n_28284), .b(n_28428), .c(n_28252), .o(n_28478) );
na02f80 g763572 ( .a(n_16933), .b(n_16898), .o(n_17128) );
in01f80 newInst_2979 ( .a(newNet_2978), .o(newNet_2979) );
ms00f80 sin_out_reg_24_ ( .ck(newNet_48), .d(n_43910), .o(sin_out_24) );
no02f80 g770576 ( .a(n_10106), .b(n_10105), .o(n_10197) );
no02f80 g778680 ( .a(n_2365), .b(n_2363), .o(n_2449) );
in01f80 g771781 ( .a(n_9177), .o(n_9178) );
in01f80 FE_RC_1798_0 ( .a(n_46955), .o(FE_RN_531_0) );
in01f80 g779641 ( .a(n_1499), .o(n_1500) );
in01f80 g752349 ( .a(n_27827), .o(n_27828) );
no02f80 g765830 ( .a(n_14932), .b(FE_OCP_RBN2503_n_13896), .o(n_15017) );
oa12f80 g752982 ( .a(n_26877), .b(n_27028), .c(n_26822), .o(n_27075) );
in01f80 g762028 ( .a(n_18335), .o(n_18336) );
in01f80 g764745 ( .a(n_15808), .o(n_15853) );
no02f80 g739346 ( .a(n_45147), .b(delay_add_ln22_unr27_stage10_stallmux_q_14_), .o(n_40704) );
no02f80 g742194 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37871), .o(n_38276) );
ao12f80 g737290 ( .a(n_42420), .b(n_42864), .c(n_42463), .o(n_42912) );
na02f80 g757981 ( .a(n_22079), .b(n_22047), .o(n_22167) );
no02f80 g775002 ( .a(n_6132), .b(n_6131), .o(n_6153) );
no02f80 g752942 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n_27876) );
oa12f80 g764768 ( .a(n_15891), .b(n_15890), .c(n_15889), .o(n_15979) );
na02f80 g750084 ( .a(n_30896), .b(n_30234), .o(n_30969) );
oa22f80 FE_RC_2975_0 ( .a(FE_OFN751_n_45003), .b(FE_OCP_RBN1363_n_20412), .c(n_45065), .d(n_20412), .o(n_20542) );
in01f80 g768759 ( .a(n_12144), .o(n_12112) );
in01f80 newInst_1474 ( .a(newNet_1473), .o(newNet_1474) );
in01f80 FE_OCP_RBC3379_n_7073 ( .a(n_7073), .o(FE_OCP_RBN3379_n_7073) );
in01f80 g766747 ( .a(n_13879), .o(n_13880) );
no02f80 g769557 ( .a(n_11328), .b(n_11280), .o(n_11355) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_1_ ( .ck(newNet_1232), .d(n_4031), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_) );
no02f80 g741995 ( .a(n_38333), .b(n_38313), .o(n_38402) );
in01f80 g775901 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_6_), .o(n_5268) );
na02f80 g776099 ( .a(FE_OCP_RBN2862_n_5024), .b(n_4441), .o(n_5102) );
no02f80 g750406 ( .a(n_29605), .b(n_29580), .o(n_29657) );
na02f80 g746972 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_24_), .o(n_32959) );
no02f80 g776924 ( .a(n_47015), .b(n_3788), .o(n_3893) );
in01f80 g775533 ( .a(n_5572), .o(n_5596) );
in01f80 g739354 ( .a(n_40814), .o(n_40815) );
na02f80 g752928 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_28212) );
in01f80 FE_OCP_RBC2692_FE_OCPN843_n_3912 ( .a(FE_OCPN843_n_3912), .o(FE_OCP_RBN2692_FE_OCPN843_n_3912) );
in01f80 g771192 ( .a(n_9573), .o(n_9574) );
no02f80 g757654 ( .a(n_22675), .b(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n_22676) );
na02f80 g739884 ( .a(n_40200), .b(n_39862), .o(n_40234) );
oa22f80 g738863 ( .a(n_41253), .b(n_40906), .c(n_41252), .d(n_40907), .o(n_41563) );
no02f80 g764565 ( .a(n_16007), .b(n_14452), .o(n_16009) );
no02f80 g765989 ( .a(n_14617), .b(n_14635), .o(n_14721) );
in01f80 g774657 ( .a(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_7217) );
in01f80 g771732 ( .a(n_10484), .o(n_8937) );
oa22f80 FE_RC_1686_0 ( .a(n_17881), .b(FE_OCPN968_n_19342), .c(n_19418), .d(n_19372), .o(n_19450) );
na02f80 g743128 ( .a(n_36914), .b(n_36934), .o(n_37211) );
in01f80 g770264 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .o(n_10812) );
na02f80 FE_RC_361_0 ( .a(n_17332), .b(FE_RN_107_0), .o(n_17457) );
no02f80 g759757 ( .a(n_21378), .b(n_21377), .o(n_22052) );
in01f80 g766474 ( .a(n_14149), .o(n_14169) );
no02f80 g744076 ( .a(n_44222), .b(n_34932), .o(n_36148) );
na02f80 g763453 ( .a(n_17115), .b(n_17167), .o(n_17315) );
in01f80 g774223 ( .a(n_6731), .o(n_6732) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_11_ ( .ck(newNet_1651), .d(n_27094), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_11_) );
na03f80 g764203 ( .a(n_16379), .b(n_16371), .c(n_16329), .o(n_16469) );
oa22f80 FE_RC_2366_0 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .b(n_1742), .c(n_1686), .d(n_1787), .o(FE_RN_917_0) );
no02f80 g751837 ( .a(n_28074), .b(n_28045), .o(n_28127) );
in01f80 g775442 ( .a(n_5785), .o(n_5786) );
oa22f80 g770720 ( .a(FE_OCP_RBN3652_n_10100), .b(n_8865), .c(FE_OCP_RBN3654_n_10100), .d(n_8908), .o(n_10305) );
na02f80 g748807 ( .a(n_32491), .b(n_32490), .o(n_33118) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_20_ ( .ck(newNet_1230), .d(n_5922), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_) );
no02f80 g779180 ( .a(FE_OCP_RBN2176_n_1864), .b(n_1668), .o(n_1916) );
in01f80 g744781 ( .a(n_35123), .o(n_35084) );
na02f80 g762371 ( .a(FE_OFN750_n_45003), .b(n_18572), .o(n_18841) );
oa12f80 g768402 ( .a(n_12414), .b(n_12381), .c(FE_OCPN1002_n_45660), .o(n_12734) );
na02f80 g749938 ( .a(n_29985), .b(FE_OCP_RBN1906_n_29080), .o(n_29961) );
in01f80 FE_OCPC3765_FE_OCP_RBN2222_n_13010 ( .a(FE_OCPN3764_FE_OCP_RBN2222_n_13010), .o(FE_OCPN3765_FE_OCP_RBN2222_n_13010) );
na02f80 g768011 ( .a(n_12633), .b(n_12649), .o(n_12681) );
oa12f80 g748995 ( .a(n_30877), .b(n_30942), .c(n_31003), .o(n_31053) );
no02f80 g776691 ( .a(FE_OCP_RBN2584_n_3858), .b(n_3857), .o(n_3916) );
in01f80 fopt782963 ( .a(n_44426), .o(n_44425) );
in01f80 g768036 ( .a(n_13075), .o(n_13076) );
in01f80 g738106 ( .a(n_42100), .o(n_42112) );
no02f80 g747172 ( .a(n_32851), .b(n_32652), .o(n_32852) );
no03m80 FE_RC_2805_0 ( .a(n_25272), .b(n_25359), .c(FE_RN_1200_0), .o(n_25458) );
na02f80 g754328 ( .a(n_25812), .b(n_25538), .o(n_25854) );
in01f80 newInst_1973 ( .a(newNet_1972), .o(newNet_1973) );
na02f80 g752660 ( .a(n_27404), .b(n_27139), .o(n_27476) );
no02f80 g758308 ( .a(FE_OCPN991_n_22249), .b(n_21278), .o(n_22461) );
oa22f80 FE_RC_3782_0 ( .a(n_17031), .b(n_17513), .c(n_17071), .d(n_17492), .o(n_17685) );
oa12f80 g758001 ( .a(n_22725), .b(n_22759), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n_22848) );
no02f80 g770206 ( .a(n_10620), .b(n_10574), .o(n_10711) );
in01f80 g752841 ( .a(n_28023), .o(n_28024) );
no02f80 g776160 ( .a(n_4743), .b(n_4609), .o(n_4772) );
na02f80 g769695 ( .a(n_11242), .b(n_11156), .o(n_11273) );
ao12f80 g771039 ( .a(n_9366), .b(n_9496), .c(n_9213), .o(n_9625) );
in01f80 g747568 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_24_), .o(n_32283) );
oa12f80 g758639 ( .a(n_21825), .b(n_22430), .c(n_21772), .o(n_22523) );
no02f80 g763109 ( .a(n_45450), .b(delay_xor_ln22_unr12_stage5_stallmux_q_7_), .o(n_17547) );
in01f80 newInst_2887 ( .a(newNet_2886), .o(newNet_2887) );
na02f80 g760578 ( .a(n_19881), .b(n_19941), .o(n_19999) );
no02f80 g755160 ( .a(n_25201), .b(n_24201), .o(n_25295) );
no02f80 g756015 ( .a(n_25139), .b(n_25138), .o(n_25191) );
oa22f80 g779358 ( .a(n_1578), .b(FE_OCPN3753_n_1448), .c(n_1577), .d(n_1449), .o(n_1660) );
no02f80 g741152 ( .a(FE_OCP_RBN2689_n_38870), .b(n_39181), .o(n_39203) );
na02f80 g750151 ( .a(n_30895), .b(n_30255), .o(n_30924) );
na02f80 g769186 ( .a(n_11976), .b(n_11897), .o(n_11898) );
na02f80 g773595 ( .a(n_7363), .b(n_7197), .o(n_7405) );
na02f80 g767913 ( .a(n_12920), .b(n_13621), .o(n_13038) );
in01f80 g742753 ( .a(n_37317), .o(n_37379) );
in01f80 g745974 ( .a(n_35277), .o(n_35278) );
ao22s80 FE_RC_1500_0 ( .a(n_20279), .b(n_20376), .c(n_20280), .d(n_20344), .o(n_20504) );
in01f80 g770938 ( .a(n_10013), .o(n_9964) );
no02f80 g761442 ( .a(n_19611), .b(n_19610), .o(n_19612) );
in01f80 g754823 ( .a(n_25401), .o(n_25362) );
na02f80 g750338 ( .a(n_29749), .b(n_29550), .o(n_29750) );
in01f80 g773724 ( .a(n_7237), .o(n_7238) );
na02f80 FE_RC_3659_0 ( .a(FE_RN_1606_0), .b(n_21658), .o(FE_RN_1605_0) );
oa22f80 FE_RC_1250_0 ( .a(n_28824), .b(n_29343), .c(n_29344), .d(n_28825), .o(n_29485) );
in01f80 FE_OCPC1750_n_27223 ( .a(FE_OCPN1749_n_27223), .o(FE_OCPN1750_n_27223) );
no02f80 g755035 ( .a(n_25127), .b(n_25126), .o(n_25431) );
na02f80 g740976 ( .a(n_39139), .b(n_39141), .o(n_39142) );
in01f80 g749495 ( .a(n_30510), .o(n_30511) );
ao12f80 g751425 ( .a(n_28460), .b(n_28631), .c(n_28630), .o(n_28649) );
in01f80 g753520 ( .a(n_27537), .o(n_27538) );
in01f80 g741742 ( .a(n_38498), .o(n_38953) );
no02f80 g754167 ( .a(n_26136), .b(n_26075), .o(n_26137) );
na02f80 g769177 ( .a(n_11546), .b(n_11634), .o(n_11635) );
no02f80 g751742 ( .a(n_29246), .b(n_29245), .o(n_29247) );
no02f80 g754094 ( .a(n_26098), .b(n_23317), .o(n_26121) );
na02f80 g777062 ( .a(n_5328), .b(n_5387), .o(n_6250) );
no02f80 g744140 ( .a(n_35690), .b(n_35567), .o(n_35689) );
na02f80 g758373 ( .a(FE_OCP_RBN1847_n_22068), .b(n_20691), .o(n_22185) );
no02f80 g744465 ( .a(n_35459), .b(n_35430), .o(n_35488) );
ao12f80 g736283 ( .a(n_43422), .b(n_43885), .c(n_43520), .o(n_43894) );
in01f80 g750254 ( .a(n_29831), .o(n_29841) );
na02f80 g765214 ( .a(n_16342), .b(n_16341), .o(n_16343) );
no02f80 g768302 ( .a(n_12535), .b(n_12051), .o(n_12573) );
in01f80 newInst_530 ( .a(newNet_529), .o(newNet_530) );
na02f80 g771584 ( .a(n_9026), .b(n_9006), .o(n_9115) );
no02f80 g756479 ( .a(n_23765), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n_23766) );
in01f80 newInst_883 ( .a(newNet_882), .o(newNet_883) );
in01f80 g778068 ( .a(n_3101), .o(n_3043) );
na02f80 g740165 ( .a(n_39816), .b(n_39917), .o(n_39950) );
ao12f80 g739052 ( .a(n_41129), .b(n_41128), .c(n_41127), .o(n_41173) );
in01f80 g768426 ( .a(n_12475), .o(n_12476) );
no02f80 g748140 ( .a(n_31931), .b(n_31902), .o(n_31948) );
no02f80 g757930 ( .a(n_22049), .b(n_21921), .o(n_22088) );
no03m80 FE_RC_3679_0 ( .a(n_33380), .b(n_33160), .c(n_33159), .o(FE_RN_885_0) );
in01f80 FE_OCP_RBC2825_n_15231 ( .a(n_15231), .o(FE_OCP_RBN2825_n_15231) );
ao22s80 g774096 ( .a(n_6679), .b(n_6613), .c(n_6734), .d(n_6612), .o(n_6804) );
ao12f80 g784144 ( .a(n_45894), .b(n_37825), .c(n_37790), .o(n_45895) );
in01f80 g766453 ( .a(n_14228), .o(n_14266) );
no02f80 g745844 ( .a(n_44102), .b(n_34003), .o(n_34283) );
in01f80 newInst_1686 ( .a(newNet_1260), .o(newNet_1686) );
na02f80 g742911 ( .a(n_36959), .b(n_37074), .o(n_37120) );
in01f80 FE_RC_2021_0 ( .a(FE_RN_671_0), .o(n_20422) );
no02f80 g736783 ( .a(n_43316), .b(n_42980), .o(n_43317) );
in01f80 newInst_23 ( .a(newNet_22), .o(newNet_23) );
in01f80 FE_RC_307_0 ( .a(n_21535), .o(FE_RN_91_0) );
na02f80 g775925 ( .a(n_5157), .b(n_5156), .o(n_5158) );
in01f80 g751353 ( .a(n_28805), .o(n_28806) );
in01f80 g758684 ( .a(n_21961), .o(n_21982) );
ao12f80 g760075 ( .a(n_21021), .b(n_21050), .c(n_21020), .o(n_21720) );
no02f80 g744978 ( .a(n_34994), .b(n_34993), .o(n_34995) );
oa22f80 FE_RC_3345_0 ( .a(n_26493), .b(n_26849), .c(n_26494), .d(n_26848), .o(n_27010) );
in01f80 g779701 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_6_), .o(n_1363) );
in01f80 FE_OCP_RBC3081_n_16977 ( .a(FE_OCP_RBN3080_n_16977), .o(FE_OCP_RBN3081_n_16977) );
na02f80 g749207 ( .a(n_30805), .b(n_30768), .o(n_30914) );
in01f80 g736859 ( .a(n_43615), .o(n_43616) );
no02f80 g755463 ( .a(n_24801), .b(n_24782), .o(n_24894) );
no02f80 g761149 ( .a(n_19058), .b(n_18975), .o(n_19147) );
in01f80 g768191 ( .a(FE_OCP_RBN2250_n_13017), .o(n_13418) );
in01f80 g771349 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_9777) );
in01f80 g745080 ( .a(FE_OCPN1422_n_35611), .o(n_34899) );
ms00f80 state_cordic_reg_1_ ( .ck(newNet_3699), .d(rst), .o(state_cordic_1_) );
in01f80 g780149 ( .a(n_1169), .o(n_1158) );
in01f80 g746825 ( .a(n_33019), .o(n_33020) );
in01f80 fopt783534 ( .a(n_45144), .o(n_45147) );
ao12f80 g751264 ( .a(n_29250), .b(n_29722), .c(n_29203), .o(n_29802) );
no02f80 g758123 ( .a(n_44267), .b(n_21413), .o(n_22198) );
no02f80 g759627 ( .a(n_20548), .b(n_20615), .o(n_20690) );
na02f80 g767372 ( .a(n_13620), .b(n_13602), .o(n_13603) );
na02f80 g743571 ( .a(n_36471), .b(n_36488), .o(n_36549) );
na02f80 g775423 ( .a(n_5824), .b(n_5886), .o(n_5899) );
in01f80 g738286 ( .a(n_42212), .o(n_41910) );
oa22f80 FE_RC_3805_0 ( .a(n_20620), .b(n_20499), .c(n_20465), .d(n_20653), .o(n_20804) );
oa12f80 g739834 ( .a(n_40064), .b(n_40432), .c(n_39931), .o(n_40448) );
in01f80 FE_OCP_RBC1143_n_29292 ( .a(n_29292), .o(FE_OCP_RBN1143_n_29292) );
no02f80 g759205 ( .a(n_21837), .b(n_21836), .o(n_21909) );
in01f80 g744930 ( .a(n_35049), .o(n_35050) );
oa12f80 FE_RC_4260_0 ( .a(FE_RN_1876_0), .b(n_22801), .c(n_22596), .o(n_22629) );
ao12f80 g742362 ( .a(n_37767), .b(n_37799), .c(n_37818), .o(n_37863) );
na02f80 g746127 ( .a(n_33803), .b(n_33826), .o(n_33874) );
na02f80 g779785 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_1_), .o(n_1395) );
in01f80 FE_OCP_RBC3138_n_40568 ( .a(n_40568), .o(FE_OCP_RBN3138_n_40568) );
na02f80 g747259 ( .a(n_33748), .b(n_33495), .o(n_33764) );
na02f80 g779380 ( .a(n_1533), .b(n_1529), .o(n_1530) );
no02f80 g779771 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_), .o(n_1470) );
in01f80 fopt783231 ( .a(n_44775), .o(n_44776) );
in01f80 g779396 ( .a(n_1571), .o(n_1572) );
no02f80 g748725 ( .a(n_31062), .b(n_31063), .o(n_31142) );
na02f80 g743427 ( .a(n_36651), .b(n_36750), .o(n_36652) );
no02f80 FE_RC_3016_0 ( .a(delay_sub_ln23_0_unr22_stage8_stallmux_q), .b(FE_RN_1322_0), .o(FE_RN_1323_0) );
no02f80 g737509 ( .a(n_42475), .b(n_42631), .o(n_42649) );
no02f80 g758250 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_14_), .o(n_22918) );
na02f80 g780403 ( .a(n_784), .b(n_7), .o(n_785) );
no02f80 g771268 ( .a(n_9255), .b(n_9113), .o(n_9314) );
in01f80 g756353 ( .a(n_23892), .o(n_23893) );
in01f80 newInst_881 ( .a(newNet_80), .o(newNet_881) );
in01f80 g751560 ( .a(n_28533), .o(n_28492) );
na02f80 g745072 ( .a(n_34728), .b(n_34282), .o(n_34755) );
no02f80 g773879 ( .a(n_7044), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_9_), .o(n_7068) );
in01f80 g760078 ( .a(n_20578), .o(n_20579) );
in01f80 g770281 ( .a(n_10834), .o(n_10835) );
ao12f80 g756337 ( .a(n_24456), .b(n_24455), .c(n_24454), .o(n_24541) );
oa22f80 FE_RC_3377_0 ( .a(n_20194), .b(n_20047), .c(n_20046), .d(n_20174), .o(n_20273) );
in01f80 newInst_1496 ( .a(newNet_1495), .o(newNet_1496) );
na02f80 g778771 ( .a(n_2297), .b(delay_add_ln22_unr2_stage2_stallmux_q_21_), .o(n_2386) );
no02f80 g753112 ( .a(n_27141), .b(n_27170), .o(n_27226) );
in01f80 g779929 ( .a(FE_OCP_RBN3242_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1852) );
in01f80 g774761 ( .a(n_6356), .o(n_6357) );
in01f80 newInst_2338 ( .a(newNet_2337), .o(newNet_2338) );
na02f80 g765994 ( .a(n_14666), .b(n_14694), .o(n_14768) );
na02f80 g778722 ( .a(n_2365), .b(n_2898), .o(n_2436) );
in01f80 newInst_398 ( .a(newNet_397), .o(newNet_398) );
no02f80 g781254 ( .a(n_69), .b(n_152), .o(n_251) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_24_ ( .ck(newNet_1727), .d(n_22545), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_) );
in01f80 g776851 ( .a(n_3830), .o(n_3831) );
na02f80 g771813 ( .a(n_8800), .b(n_8610), .o(n_8839) );
no02f80 g759433 ( .a(n_20932), .b(n_20713), .o(n_20997) );
in01f80 g747669 ( .a(n_33297), .o(n_34070) );
in01f80 g775820 ( .a(n_5071), .o(n_5072) );
na02f80 g772408 ( .a(n_8420), .b(n_8540), .o(n_8627) );
in01f80 newInst_2778 ( .a(newNet_2777), .o(newNet_2778) );
in01f80 g745352 ( .a(n_36155), .o(n_36156) );
no02f80 g745890 ( .a(n_34040), .b(n_34014), .o(n_34097) );
no02f80 FE_RC_3112_0 ( .a(FE_RN_1377_0), .b(n_32086), .o(n_31880) );
in01f80 g742570 ( .a(n_37556), .o(n_37574) );
in01f80 g775552 ( .a(n_5456), .o(n_5457) );
in01f80 g747588 ( .a(n_32364), .o(n_32365) );
no02f80 g762341 ( .a(FE_OCP_RBN3410_n_45120), .b(n_18422), .o(n_18453) );
no02f80 g776053 ( .a(n_4581), .b(n_4544), .o(n_4729) );
no02f80 g772373 ( .a(n_8441), .b(n_8522), .o(n_8601) );
no02f80 g766758 ( .a(n_14489), .b(n_14528), .o(n_14529) );
oa12f80 g768807 ( .a(n_11687), .b(n_11929), .c(n_11635), .o(n_12065) );
in01f80 newInst_2566 ( .a(newNet_2565), .o(newNet_2566) );
na02f80 g777658 ( .a(n_3511), .b(n_3458), .o(n_3528) );
in01f80 g772539 ( .a(n_8354), .o(n_8376) );
in01f80 g772687 ( .a(n_8101), .o(n_8111) );
in01f80 g746014 ( .a(n_34055), .o(n_34056) );
in01f80 g756559 ( .a(n_23757), .o(n_23758) );
na02f80 g773810 ( .a(n_7117), .b(n_7116), .o(n_7505) );
no02f80 g773003 ( .a(n_8027), .b(n_7954), .o(n_7955) );
no02f80 g742606 ( .a(n_37427), .b(n_37451), .o(n_37559) );
na02f80 g775979 ( .a(n_5134), .b(n_5042), .o(n_5169) );
no02f80 g779545 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .o(n_1878) );
no02f80 g749954 ( .a(n_29895), .b(n_29865), .o(n_30225) );
na02f80 g748439 ( .a(n_31474), .b(FE_OCPN1446_n_31473), .o(n_31521) );
in01f80 newInst_1024 ( .a(newNet_1023), .o(newNet_1024) );
ao12f80 g747690 ( .a(n_32108), .b(n_32238), .c(n_32021), .o(n_32280) );
oa22f80 g739635 ( .a(n_40593), .b(n_40598), .c(n_40584), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_40599) );
oa12f80 g747350 ( .a(n_33579), .b(n_33578), .c(n_33359), .o(n_33630) );
na02f80 g784080 ( .a(n_7654), .b(n_45820), .o(n_45826) );
in01f80 g756421 ( .a(n_23640), .o(n_23694) );
na02f80 g763287 ( .a(n_16911), .b(n_17039), .o(n_17088) );
in01f80 g768397 ( .a(n_12539), .o(n_12540) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_0_ ( .ck(newNet_2328), .d(n_39716), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_0_) );
na02f80 g770894 ( .a(n_9864), .b(FE_OCPN1255_n_8499), .o(n_10016) );
in01f80 newInst_1085 ( .a(newNet_1084), .o(newNet_1085) );
na02f80 g744993 ( .a(n_34928), .b(n_34748), .o(n_34990) );
no02f80 g739483 ( .a(FE_OCPN932_n_40736), .b(n_40479), .o(n_40711) );
in01f80 g755991 ( .a(n_24229), .o(n_24230) );
in01f80 FE_OCPC1783_n_26801 ( .a(n_26801), .o(FE_OCPN1783_n_26801) );
in01f80 g737244 ( .a(n_46937), .o(n_43179) );
in01f80 g767492 ( .a(n_13097), .o(n_13151) );
no02f80 g773741 ( .a(n_7246), .b(n_7099), .o(n_7287) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_8_ ( .ck(newNet_769), .d(n_1315), .o(delay_xor_ln21_unr3_stage2_stallmux_q_8_) );
in01f80 g739905 ( .a(n_40339), .o(n_40340) );
no02f80 g759218 ( .a(FE_OCP_RBN1726_n_20924), .b(n_20943), .o(n_20982) );
na02f80 g753486 ( .a(n_26788), .b(n_26764), .o(n_26765) );
no02f80 g756545 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n_23638) );
na02f80 g744521 ( .a(n_35386), .b(n_35410), .o(n_35449) );
in01f80 g767744 ( .a(n_46414), .o(n_13129) );
in01f80 g778741 ( .a(n_2402), .o(n_2378) );
no02f80 FE_RC_1167_0 ( .a(FE_RN_353_0), .b(n_28013), .o(n_28125) );
oa12f80 g753303 ( .a(n_27057), .b(n_27024), .c(n_27073), .o(n_27074) );
in01f80 newInst_2356 ( .a(newNet_2355), .o(newNet_2356) );
na02f80 g760915 ( .a(n_19330), .b(n_19279), .o(n_19388) );
in01f80 g747166 ( .a(n_34547), .o(n_33992) );
no02f80 g780087 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_11_), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_12_), .o(n_1193) );
no02f80 g738584 ( .a(n_41487), .b(n_41458), .o(n_41890) );
na02f80 g766492 ( .a(n_13927), .b(FE_OCP_RBN2246_n_13017), .o(n_13959) );
no02f80 g754215 ( .a(FE_OCP_RBN1202_n_25898), .b(n_23254), .o(n_26004) );
no02f80 g750114 ( .a(FE_OCP_RBN3567_n_29857), .b(FE_OCP_RBN1144_n_29292), .o(n_30116) );
na02f80 g761332 ( .a(n_20082), .b(n_20113), .o(n_20256) );
ms00f80 delay_xor_ln21_unr28_stage10_stallmux_q_reg_0_ ( .ck(newNet_865), .d(n_40591), .o(delay_xor_ln21_unr28_stage10_stallmux_q_0_) );
no02f80 g774346 ( .a(n_6582), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n_6583) );
in01f80 FE_OCP_RBC2451_n_34278 ( .a(n_34278), .o(FE_OCP_RBN2451_n_34278) );
in01f80 FE_OCP_RBC2850_n_46982 ( .a(FE_OCP_RBN2849_n_46982), .o(FE_OCP_RBN2850_n_46982) );
no02f80 g757009 ( .a(n_47337), .b(n_23267), .o(n_23329) );
in01f80 newInst_3317 ( .a(newNet_2405), .o(newNet_3317) );
in01f80 g760359 ( .a(n_20222), .o(n_20223) );
in01f80 g742789 ( .a(n_37384), .o(n_37385) );
oa22f80 g742039 ( .a(FE_OCP_RBN3451_n_37945), .b(FE_OCP_RBN2188_n_37686), .c(FE_OCP_RBN3452_n_37945), .d(FE_OCP_RBN2187_n_37686), .o(n_38258) );
oa12f80 g780014 ( .a(n_977), .b(n_1259), .c(n_925), .o(n_1267) );
no02f80 g745154 ( .a(n_34820), .b(n_34399), .o(n_34749) );
in01f80 FE_OCP_RBC3533_n_13765 ( .a(FE_OCP_RBN3530_n_13765), .o(FE_OCP_RBN3533_n_13765) );
no02f80 g756833 ( .a(n_23936), .b(n_23868), .o(n_23956) );
in01f80 g746495 ( .a(n_33273), .o(n_33291) );
no02f80 g761727 ( .a(n_19401), .b(n_19367), .o(n_19368) );
ao12f80 g767658 ( .a(n_12823), .b(n_13000), .c(n_13013), .o(n_13047) );
in01f80 newInst_2972 ( .a(newNet_2971), .o(newNet_2972) );
na02f80 g759006 ( .a(n_21531), .b(n_21496), .o(n_22039) );
in01f80 g764225 ( .a(n_16526), .o(n_16552) );
na02f80 g769099 ( .a(n_11510), .b(n_11516), .o(n_11596) );
na02f80 g777874 ( .a(n_3221), .b(FE_OCP_RBN2424_n_47023), .o(n_3277) );
ao12f80 g767489 ( .a(n_13292), .b(n_13291), .c(n_13290), .o(n_14977) );
na03f80 FE_RC_3680_0 ( .a(FE_RN_1031_0), .b(n_23109), .c(n_45312), .o(n_23195) );
na02f80 g774915 ( .a(n_6100), .b(n_6000), .o(n_6122) );
na02f80 g779044 ( .a(n_2044), .b(n_1899), .o(n_2106) );
na02f80 g775166 ( .a(n_5994), .b(n_5990), .o(n_5991) );
in01f80 g745373 ( .a(n_35799), .o(n_35888) );
in01f80 g759082 ( .a(n_21959), .o(n_22011) );
oa12f80 g752121 ( .a(n_28668), .b(n_28667), .c(n_28666), .o(n_29067) );
in01f80 FE_OCPC1029_n_28423 ( .a(n_28423), .o(FE_OCPN1029_n_28423) );
na02f80 g745720 ( .a(n_34259), .b(n_44102), .o(n_34307) );
no02f80 g751582 ( .a(n_28817), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(n_28842) );
no02f80 g754386 ( .a(n_25734), .b(n_25706), .o(n_25816) );
ao12f80 g767837 ( .a(n_12725), .b(FE_OCPN3757_n_13889), .c(n_12724), .o(n_12795) );
no02f80 g775725 ( .a(n_5462), .b(FE_OCP_RBN2702_n_4041), .o(n_5577) );
in01f80 g740070 ( .a(n_40139), .o(n_40140) );
no02f80 g755430 ( .a(n_24656), .b(n_24386), .o(n_24700) );
na02f80 g773104 ( .a(n_7880), .b(n_7923), .o(n_7924) );
in01f80 newInst_3048 ( .a(newNet_3047), .o(newNet_3048) );
no02f80 g760863 ( .a(n_19365), .b(n_18786), .o(n_19393) );
in01f80 g737376 ( .a(n_42813), .o(n_42814) );
no02f80 g751052 ( .a(n_30088), .b(n_30063), .o(n_30064) );
ao12f80 g760162 ( .a(n_20052), .b(n_20953), .c(n_19959), .o(n_21102) );
in01f80 FE_OCPC1052_n_31674 ( .a(FE_OCPN1051_n_31674), .o(FE_OCPN1052_n_31674) );
in01f80 FE_RC_1281_0 ( .a(n_2333), .o(FE_RN_378_0) );
in01f80 g776829 ( .a(n_3737), .o(n_3738) );
no02f80 g747311 ( .a(n_33628), .b(n_33627), .o(n_45753) );
na02f80 g761434 ( .a(n_18829), .b(n_18370), .o(n_18876) );
no02f80 g763040 ( .a(n_17415), .b(n_17405), .o(n_17510) );
no02f80 g758262 ( .a(FE_OCP_RBN2050_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_11_), .o(n_22692) );
in01f80 newInst_896 ( .a(newNet_5), .o(newNet_896) );
na02f80 g759979 ( .a(n_20469), .b(n_20374), .o(n_20470) );
no02f80 g771859 ( .a(n_9954), .b(n_10039), .o(n_10841) );
ao12f80 g743474 ( .a(n_37674), .b(n_37673), .c(n_37672), .o(n_37749) );
ao12f80 g779462 ( .a(n_1972), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_22_), .o(n_2019) );
in01f80 fopt783997 ( .a(n_22564), .o(n_45721) );
na02f80 g747159 ( .a(n_32886), .b(n_32885), .o(n_32887) );
oa22f80 g752698 ( .a(n_27242), .b(n_27214), .c(n_27241), .d(n_27215), .o(n_27364) );
in01f80 g743656 ( .a(n_36378), .o(n_36379) );
in01f80 g761548 ( .a(n_18996), .o(n_18997) );
na02f80 g760555 ( .a(n_19865), .b(n_18230), .o(n_19973) );
na02f80 g751877 ( .a(n_29025), .b(n_29045), .o(n_29046) );
na02f80 g771624 ( .a(n_9355), .b(n_9237), .o(n_9438) );
no02f80 g745406 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35765), .o(n_36079) );
in01f80 g742812 ( .a(n_37277), .o(n_37278) );
in01f80 g766038 ( .a(n_14714), .o(n_14715) );
na02f80 g769067 ( .a(n_11552), .b(n_11580), .o(n_11656) );
na02f80 FE_RC_2876_0 ( .a(FE_RN_1241_0), .b(n_20070), .o(FE_RN_1242_0) );
na02f80 g770228 ( .a(n_10568), .b(n_44463), .o(n_10594) );
oa12f80 g742017 ( .a(n_37947), .b(FE_OCP_RBN3445_n_37945), .c(n_37981), .o(n_38426) );
in01f80 newInst_421 ( .a(newNet_420), .o(newNet_421) );
no02f80 g744543 ( .a(n_35365), .b(FE_OCP_RBN2666_n_35207), .o(n_35370) );
na02f80 g738819 ( .a(n_41313), .b(delay_sub_ln23_0_unr28_stage10_stallmux_q), .o(n_41329) );
oa12f80 g754879 ( .a(n_25008), .b(n_25128), .c(n_25066), .o(n_25247) );
na02f80 g747372 ( .a(n_32401), .b(n_44962), .o(n_32577) );
in01f80 g762921 ( .a(n_17718), .o(n_17719) );
na02f80 g758894 ( .a(n_21360), .b(n_45072), .o(n_21395) );
in01f80 g749087 ( .a(n_31018), .o(n_31048) );
in01f80 FE_OCPC1429_n_23792 ( .a(n_23792), .o(FE_OCPN1429_n_23792) );
in01f80 newInst_2282 ( .a(newNet_1875), .o(newNet_2282) );
oa22f80 FE_RC_1625_0 ( .a(n_32209), .b(n_32236), .c(n_32208), .d(n_32237), .o(n_32281) );
in01f80 g761035 ( .a(n_19344), .o(n_19374) );
na02f80 g780519 ( .a(n_842), .b(n_829), .o(n_843) );
in01f80 FE_RC_2723_0 ( .a(n_8326), .o(FE_RN_1151_0) );
in01f80 FE_OCP_RBC2862_n_5024 ( .a(n_5024), .o(FE_OCP_RBN2862_n_5024) );
no02f80 g760085 ( .a(n_21050), .b(n_21020), .o(n_21021) );
in01f80 FE_RC_3490_0 ( .a(FE_RN_1504_0), .o(FE_RN_1503_0) );
no02f80 g759155 ( .a(n_21275), .b(n_21314), .o(n_21466) );
in01f80 newInst_1757 ( .a(newNet_1189), .o(newNet_1757) );
in01f80 fopt783507 ( .a(n_45002), .o(n_45003) );
in01f80 g760631 ( .a(n_19854), .o(n_19938) );
in01f80 newInst_2790 ( .a(newNet_2789), .o(newNet_2790) );
ao22s80 g778566 ( .a(n_2213), .b(n_1489), .c(n_2212), .d(n_1490), .o(n_2285) );
na02f80 g759460 ( .a(n_20908), .b(n_45032), .o(n_20995) );
na02f80 g775335 ( .a(n_5558), .b(n_5649), .o(n_5677) );
in01f80 g765559 ( .a(n_15127), .o(n_15258) );
no02f80 g769116 ( .a(n_47279), .b(n_11622), .o(n_11801) );
in01f80 g746372 ( .a(n_33604), .o(n_33605) );
na02f80 g759077 ( .a(n_21130), .b(n_20668), .o(n_21165) );
in01f80 g757513 ( .a(n_22778), .o(n_22757) );
no02f80 g775763 ( .a(n_5421), .b(n_5051), .o(n_5532) );
oa22f80 FE_RC_1483_0 ( .a(n_32287), .b(FE_OCP_RBN3142_n_32395), .c(n_28336), .d(n_32395), .o(n_32515) );
na02f80 g741724 ( .a(n_46417), .b(n_38199), .o(n_38546) );
oa12f80 g745029 ( .a(n_34506), .b(n_34786), .c(n_34535), .o(n_34876) );
na02f80 g770128 ( .a(n_10730), .b(FE_OCPN955_n_44460), .o(n_10792) );
in01f80 g742610 ( .a(n_37527), .o(n_37551) );
no02f80 g754498 ( .a(n_26313), .b(n_26193), .o(n_26938) );
in01f80 g780732 ( .a(n_808), .o(n_610) );
in01f80 FE_RC_1092_0 ( .a(n_17894), .o(FE_RN_321_0) );
in01f80 g759168 ( .a(n_21016), .o(n_21017) );
in01f80 g771689 ( .a(n_9201), .o(n_9130) );
in01f80 newInst_3612 ( .a(newNet_3611), .o(newNet_3612) );
in01f80 g749807 ( .a(n_31623), .o(n_31624) );
na02f80 FE_RC_399_0 ( .a(FE_RN_117_0), .b(FE_OCP_RBN2799_n_15434), .o(FE_RN_119_0) );
no02f80 g775819 ( .a(n_5276), .b(n_5231), .o(n_5317) );
na02f80 g743678 ( .a(n_36327), .b(n_35587), .o(n_36351) );
na02f80 g754042 ( .a(n_26101), .b(n_26089), .o(n_26221) );
no02f80 g769259 ( .a(n_11439), .b(n_10613), .o(n_11436) );
no02f80 g778227 ( .a(n_2674), .b(FE_OCP_RBN3487_n_2438), .o(n_2675) );
na02f80 g748645 ( .a(n_32645), .b(n_32448), .o(n_32646) );
no02f80 FE_RC_2566_0 ( .a(FE_RN_1053_0), .b(n_34632), .o(n_34661) );
ao12f80 g738994 ( .a(n_40791), .b(n_41114), .c(n_40829), .o(n_41169) );
no02f80 g764303 ( .a(n_16328), .b(n_14588), .o(n_16376) );
ao12f80 g767577 ( .a(n_13179), .b(n_13178), .c(n_13177), .o(n_13288) );
no02f80 g742252 ( .a(n_37843), .b(n_37881), .o(n_37987) );
na02f80 g767701 ( .a(n_13243), .b(n_13192), .o(n_13766) );
in01f80 g779218 ( .a(n_2255), .o(n_1871) );
in01f80 newInst_1488 ( .a(newNet_1487), .o(newNet_1488) );
in01f80 g748083 ( .a(n_31971), .o(n_31994) );
no02f80 g777850 ( .a(n_3273), .b(n_47022), .o(n_3330) );
na02f80 FE_RC_2146_0 ( .a(n_15219), .b(FE_RN_755_0), .o(FE_RN_756_0) );
in01f80 g742824 ( .a(n_37392), .o(n_37309) );
in01f80 newInst_2444 ( .a(newNet_2279), .o(newNet_2444) );
ao12f80 g781114 ( .a(n_230), .b(n_229), .c(n_228), .o(n_241) );
ao12f80 g761376 ( .a(n_19612), .b(n_19611), .c(n_19610), .o(n_19712) );
no02f80 g746266 ( .a(n_33530), .b(n_33081), .o(n_33570) );
in01f80 fopt783475 ( .a(n_45080), .o(n_45081) );
in01f80 g739978 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_4_), .o(n_40084) );
in01f80 newInst_1387 ( .a(newNet_751), .o(newNet_1387) );
ao12f80 g767997 ( .a(n_12680), .b(n_12679), .c(n_12678), .o(n_13116) );
ao12f80 g784432 ( .a(n_46218), .b(n_46204), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n_46244) );
no02f80 FE_RC_3543_0 ( .a(n_17732), .b(n_18713), .o(FE_RN_1535_0) );
no02f80 g781093 ( .a(n_247), .b(n_246), .o(n_248) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_5_ ( .ck(newNet_1002), .d(n_17004), .o(delay_xor_ln21_unr12_stage5_stallmux_q_5_) );
in01f80 FE_OCP_RBC2765_n_25895 ( .a(n_25895), .o(FE_OCP_RBN2765_n_25895) );
na02f80 g777125 ( .a(n_3828), .b(n_47023), .o(n_3873) );
no02f80 g778624 ( .a(FE_OCPN871_n_2737), .b(n_2719), .o(n_2768) );
in01f80 FE_OCP_RBC2927_n_39614 ( .a(n_39614), .o(FE_OCP_RBN2927_n_39614) );
in01f80 newInst_651 ( .a(newNet_301), .o(newNet_651) );
oa12f80 g752313 ( .a(n_28436), .b(n_28435), .c(n_28434), .o(n_28942) );
oa12f80 g779377 ( .a(n_1530), .b(n_1533), .c(n_1529), .o(n_1593) );
in01f80 newInst_128 ( .a(newNet_56), .o(newNet_128) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_25_ ( .ck(newNet_1098), .d(n_11286), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_) );
in01f80 g760174 ( .a(n_20336), .o(n_20367) );
oa22f80 FE_RC_1208_0 ( .a(FE_OCP_RBN2382_n_3502), .b(n_3055), .c(FE_OCP_RBN2380_n_3502), .d(n_3054), .o(n_3066) );
in01f80 g739553 ( .a(n_41309), .o(n_40657) );
in01f80 g759942 ( .a(n_21600), .o(n_21560) );
ao12f80 g766985 ( .a(n_13792), .b(n_13791), .c(n_13790), .o(n_13877) );
in01f80 g775221 ( .a(n_46997), .o(n_6004) );
in01f80 FE_OCP_RBC3093_n_11475 ( .a(FE_OCP_RBN3091_n_11475), .o(FE_OCP_RBN3093_n_11475) );
no02f80 g769276 ( .a(n_11627), .b(FE_OCP_RBN2887_n_10570), .o(n_11620) );
ao12f80 g746764 ( .a(n_33108), .b(n_33305), .c(n_32355), .o(n_33269) );
in01f80 FE_OCP_RBC2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2048_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01f80 FE_RC_3115_0 ( .a(n_31103), .o(FE_RN_1380_0) );
no02f80 g738735 ( .a(n_41483), .b(n_41211), .o(n_41531) );
in01f80 FE_OCP_RBC1182_n_19726 ( .a(n_19726), .o(FE_OCP_RBN1182_n_19726) );
in01f80 FE_OCP_RBC1922_cordic_combinational_sub_ln23_0_unr12_z_0__ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN1922_cordic_combinational_sub_ln23_0_unr12_z_0__) );
no02f80 g738313 ( .a(n_41737), .b(n_41736), .o(n_41738) );
in01f80 g749396 ( .a(n_30697), .o(n_30696) );
na02f80 g747332 ( .a(FE_OCP_RBN2102_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_8_), .o(n_32690) );
na02f80 g757333 ( .a(n_22970), .b(n_22937), .o(n_23002) );
na02f80 g768317 ( .a(n_12522), .b(n_12503), .o(n_12547) );
in01f80 g770919 ( .a(n_9809), .o(n_9810) );
in01f80 g774923 ( .a(n_6270), .o(n_6281) );
in01f80 g754257 ( .a(n_25982), .o(n_26055) );
in01f80 g755599 ( .a(n_25172), .o(n_25468) );
in01f80 g756702 ( .a(n_23563), .o(n_23551) );
na02f80 g771954 ( .a(FE_OFN754_n_44461), .b(n_9367), .o(n_9480) );
oa22f80 FE_RC_483_0 ( .a(n_23718), .b(n_24018), .c(n_23685), .d(n_24019), .o(n_24079) );
in01f80 FE_OCP_RBC1150_n_17239 ( .a(n_17239), .o(FE_OCP_RBN1150_n_17239) );
in01f80 FE_RC_3519_0 ( .a(n_22998), .o(FE_RN_1520_0) );
no02f80 g777833 ( .a(n_3230), .b(n_3205), .o(n_3498) );
ao12f80 g774260 ( .a(n_6583), .b(n_6582), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_1_), .o(n_7630) );
no02f80 g744123 ( .a(n_36030), .b(n_36000), .o(n_36065) );
in01f80 g743141 ( .a(n_37085), .o(n_37171) );
oa22f80 FE_RC_3456_0 ( .a(n_45010), .b(n_20622), .c(n_45012), .d(n_20621), .o(n_20771) );
in01f80 FE_OCP_RBC2464_n_4336 ( .a(n_4336), .o(FE_OCP_RBN2464_n_4336) );
no02f80 g745023 ( .a(n_34769), .b(n_34362), .o(n_34831) );
na02f80 g771286 ( .a(n_9688), .b(n_9687), .o(n_9689) );
no02f80 g762785 ( .a(n_17942), .b(delay_add_ln22_unr11_stage5_stallmux_q_10_), .o(n_17964) );
in01f80 FE_OCP_RBC3051_n_16596 ( .a(n_16596), .o(FE_OCP_RBN3051_n_16596) );
in01f80 g752110 ( .a(n_28782), .o(n_28781) );
in01f80 newInst_2758 ( .a(newNet_2757), .o(newNet_2758) );
na02f80 g741103 ( .a(n_39150), .b(n_39179), .o(n_39247) );
in01f80 g775082 ( .a(n_6019), .o(n_6020) );
no02f80 g762359 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18494), .o(n_18583) );
in01f80 newInst_2253 ( .a(newNet_586), .o(newNet_2253) );
na02f80 g779018 ( .a(n_2058), .b(n_1892), .o(n_2103) );
no02f80 g759411 ( .a(n_21036), .b(n_21035), .o(n_21062) );
oa22f80 FE_RC_3733_0 ( .a(n_15076), .b(n_15164), .c(n_15075), .d(n_15163), .o(n_15319) );
ao22s80 FE_RC_95_0 ( .a(n_18874), .b(n_18408), .c(n_18873), .d(n_18407), .o(n_18986) );
in01f80 g777000 ( .a(n_4143), .o(n_4144) );
in01f80 g770347 ( .a(n_10740), .o(n_10681) );
in01f80 newInst_77 ( .a(newNet_76), .o(newNet_77) );
in01f80 FE_OCPC1473_n_24624 ( .a(n_24624), .o(FE_OCPN1473_n_24624) );
na02f80 g748923 ( .a(n_46107), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_16_), .o(n_32485) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_31_ ( .ck(newNet_1963), .d(n_12162), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_31_) );
in01f80 FE_OCP_RBC2720_n_9494 ( .a(n_9494), .o(FE_OCP_RBN2720_n_9494) );
oa12f80 g758955 ( .a(n_21391), .b(n_21470), .c(n_21280), .o(n_21428) );
na02f80 g764929 ( .a(n_15753), .b(n_15752), .o(n_15754) );
no02f80 g780555 ( .a(FE_OCPN852_n_694), .b(n_521), .o(n_845) );
in01f80 g761460 ( .a(n_19830), .o(n_19763) );
na02f80 g746461 ( .a(n_33291), .b(n_33276), .o(n_33277) );
no02f80 FE_RC_683_0 ( .a(FE_RN_221_0), .b(n_32697), .o(n_32722) );
in01f80 FE_OCP_RBC2740_n_20565 ( .a(n_20565), .o(FE_OCP_RBN2740_n_20565) );
in01f80 FE_OCPC1858_n_22207 ( .a(FE_OCPN1857_n_22207), .o(FE_OCPN1858_n_22207) );
in01f80 FE_OCPC1020_n_23078 ( .a(FE_OCPN1018_n_23078), .o(FE_OCPN1020_n_23078) );
na02f80 g763197 ( .a(n_17280), .b(n_17398), .o(n_17434) );
no02f80 g777320 ( .a(n_3705), .b(n_3323), .o(n_3741) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_25_ ( .ck(newNet_3217), .d(n_36549), .o(delay_add_ln22_unr23_stage9_stallmux_q_25_) );
oa12f80 g773987 ( .a(n_6975), .b(n_6974), .c(n_6973), .o(n_7819) );
na02f80 g771055 ( .a(n_9359), .b(n_8232), .o(n_9579) );
oa12f80 g744110 ( .a(n_35552), .b(n_35551), .c(n_35556), .o(n_35592) );
no02f80 g740445 ( .a(n_39719), .b(n_39645), .o(n_39721) );
in01f80 FE_RC_3574_0 ( .a(n_35831), .o(FE_RN_1554_0) );
no02f80 g751721 ( .a(n_28331), .b(n_28346), .o(n_28422) );
in01f80 g736510 ( .a(n_43712), .o(n_43713) );
in01f80 g737429 ( .a(n_42780), .o(n_42750) );
no02f80 g753647 ( .a(n_26766), .b(n_26584), .o(n_26762) );
na02f80 g775406 ( .a(n_5680), .b(n_5712), .o(n_5767) );
no02f80 g756779 ( .a(n_24171), .b(n_24170), .o(n_24172) );
na02f80 g778200 ( .a(n_2799), .b(FE_OCPN3759_n_2346), .o(n_2800) );
in01f80 g767390 ( .a(n_13390), .o(n_13362) );
in01f80 FE_OCP_RBC2301_n_7817 ( .a(FE_OCP_RBN2300_n_7817), .o(FE_OCP_RBN2301_n_7817) );
in01f80 newInst_2947 ( .a(newNet_2946), .o(newNet_2947) );
na02f80 g744080 ( .a(n_44222), .b(n_35003), .o(n_36191) );
in01f80 g737686 ( .a(n_42397), .o(n_42444) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_16_ ( .ck(newNet_966), .d(n_22957), .o(delay_xor_ln21_unr15_stage6_stallmux_q_16_) );
na02f80 g768064 ( .a(n_12709), .b(n_12692), .o(n_12860) );
in01f80 FE_OCP_RBC3669_n_46982 ( .a(n_46982), .o(FE_OCP_RBN3669_n_46982) );
in01f80 g746420 ( .a(n_34123), .o(n_33500) );
ao12f80 g748102 ( .a(n_32805), .b(n_32804), .c(n_32803), .o(n_33437) );
in01f80 g753513 ( .a(n_26872), .o(n_26871) );
oa22f80 g743663 ( .a(n_36393), .b(n_35866), .c(n_36392), .d(n_35865), .o(n_36439) );
ao12f80 g738928 ( .a(n_40961), .b(n_41221), .c(n_40841), .o(n_41304) );
no02f80 g764789 ( .a(n_15755), .b(n_13879), .o(n_15938) );
na02f80 g746218 ( .a(n_35087), .b(n_34581), .o(n_35045) );
in01f80 newInst_406 ( .a(newNet_405), .o(newNet_406) );
in01f80 newInst_75 ( .a(newNet_74), .o(newNet_75) );
na02f80 g765081 ( .a(n_15200), .b(n_14215), .o(n_15240) );
na02f80 g748170 ( .a(n_31851), .b(n_32119), .o(n_32210) );
in01f80 newInst_1704 ( .a(newNet_1703), .o(newNet_1704) );
in01f80 g750352 ( .a(n_31210), .o(n_30718) );
na02f80 g781049 ( .a(sin_out_30), .b(FE_OFN4_n_43918), .o(n_294) );
in01f80 g736763 ( .a(n_43321), .o(n_43322) );
no02f80 g765886 ( .a(n_15245), .b(n_15244), .o(n_15246) );
in01f80 g750458 ( .a(n_29550), .o(n_29551) );
in01f80 g779651 ( .a(n_1771), .o(n_1772) );
na02f80 g772922 ( .a(n_8091), .b(n_7802), .o(n_7907) );
no02f80 g744745 ( .a(n_35169), .b(n_35171), .o(n_35226) );
in01f80 g754156 ( .a(n_26293), .o(n_26051) );
na02f80 g751048 ( .a(n_29854), .b(n_29853), .o(n_29879) );
oa12f80 g756790 ( .a(n_24059), .b(n_24151), .c(n_24150), .o(n_24152) );
na02f80 g739865 ( .a(n_40402), .b(n_40151), .o(n_40417) );
na02f80 g736818 ( .a(n_43133), .b(n_43217), .o(n_43263) );
na02f80 g746980 ( .a(n_33013), .b(n_33052), .o(n_33236) );
oa12f80 g737859 ( .a(n_42360), .b(n_42547), .c(n_42304), .o(n_42618) );
oa12f80 g764721 ( .a(n_15604), .b(n_15739), .c(n_15487), .o(n_15802) );
na02f80 g775312 ( .a(n_5805), .b(n_5606), .o(n_5834) );
na02f80 g775834 ( .a(n_5493), .b(n_47015), .o(n_5584) );
in01f80 g749973 ( .a(n_30259), .o(n_30260) );
no02f80 g744137 ( .a(n_35616), .b(n_35690), .o(n_35737) );
in01f80 newInst_968 ( .a(newNet_620), .o(newNet_968) );
ms00f80 sin_out_reg_7_ ( .ck(newNet_13), .d(n_43707), .o(sin_out_7) );
no02f80 g771143 ( .a(n_9509), .b(FE_OCPN1253_n_8348), .o(n_9578) );
oa12f80 g742946 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37111), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n_37112) );
no02f80 g771424 ( .a(n_9044), .b(n_9012), .o(n_9095) );
in01f80 newInst_3604 ( .a(newNet_3603), .o(newNet_3604) );
oa22f80 g758663 ( .a(n_22426), .b(n_21627), .c(n_22395), .d(n_21628), .o(n_22521) );
in01f80 g777327 ( .a(n_3768), .o(n_3769) );
in01f80 fopt783317 ( .a(FE_OCP_RBN2241_n_44881), .o(n_44887) );
na02f80 g745760 ( .a(n_34183), .b(n_34182), .o(n_34198) );
oa12f80 g737207 ( .a(n_42417), .b(n_42927), .c(n_42279), .o(n_42973) );
no02f80 g779591 ( .a(n_1410), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(n_1466) );
oa12f80 g759823 ( .a(n_21139), .b(n_21138), .c(n_21137), .o(n_21750) );
no02f80 g740638 ( .a(n_39571), .b(n_39557), .o(n_40028) );
na02f80 g754517 ( .a(n_26931), .b(n_26930), .o(n_26932) );
na02f80 g737479 ( .a(n_42552), .b(n_42314), .o(n_42567) );
oa22f80 FE_RC_1163_0 ( .a(n_12819), .b(n_13343), .c(n_12820), .d(n_13344), .o(n_13489) );
no02f80 g741006 ( .a(n_39063), .b(n_38962), .o(n_39109) );
in01f80 newInst_469 ( .a(newNet_143), .o(newNet_469) );
ao12f80 g779439 ( .a(n_1544), .b(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_9_), .o(n_1563) );
no02f80 g755291 ( .a(n_24861), .b(n_24887), .o(n_24924) );
in01f80 newInst_1545 ( .a(newNet_1544), .o(newNet_1545) );
na02f80 g775154 ( .a(n_5978), .b(n_6023), .o(n_6105) );
na02f80 g750802 ( .a(n_29097), .b(n_29065), .o(n_29163) );
na02f80 g765417 ( .a(n_15402), .b(n_15448), .o(n_15567) );
no02f80 g757838 ( .a(n_22983), .b(n_22694), .o(n_23009) );
na02f80 g771337 ( .a(n_9205), .b(n_9202), .o(n_9354) );
no02f80 g760715 ( .a(n_19606), .b(n_19642), .o(n_19752) );
oa22f80 FE_RC_36_0 ( .a(n_5556), .b(n_5674), .c(n_5557), .d(n_5675), .o(n_5813) );
in01f80 g745118 ( .a(n_34751), .o(n_34752) );
na02f80 FE_RC_3525_0 ( .a(n_27227), .b(n_27175), .o(FE_RN_1524_0) );
na02f80 g739420 ( .a(n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_30_), .o(n_40917) );
oa12f80 g747624 ( .a(n_33374), .b(n_33356), .c(n_33392), .o(n_33481) );
no02f80 g740042 ( .a(n_39983), .b(n_39982), .o(n_40018) );
no02f80 g739339 ( .a(n_40816), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_13_), .o(n_40817) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_31_ ( .ck(newNet_3285), .d(n_32310), .o(delay_add_ln22_unr20_stage8_stallmux_q_31_) );
no02f80 g760410 ( .a(n_20739), .b(n_20054), .o(n_20740) );
in01f80 newInst_1178 ( .a(newNet_1177), .o(newNet_1178) );
na02f80 g768451 ( .a(n_12398), .b(n_12354), .o(n_12596) );
in01f80 g741696 ( .a(n_38521), .o(n_38522) );
na02f80 g766214 ( .a(n_14204), .b(n_14251), .o(n_14380) );
ao12f80 g737324 ( .a(n_42300), .b(n_42812), .c(n_42327), .o(n_42844) );
ao12f80 g746846 ( .a(n_32948), .b(FE_OCP_RBN2169_n_32892), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .o(n_33262) );
in01f80 g736391 ( .a(n_43848), .o(n_43849) );
ao22s80 FE_RC_1246_0 ( .a(n_33569), .b(n_33183), .c(n_33182), .d(n_33568), .o(n_33697) );
na02f80 g784593 ( .a(FE_OCP_RBN3452_n_37945), .b(n_37567), .o(n_46416) );
in01f80 g777348 ( .a(n_5069), .o(n_5147) );
na02f80 g744100 ( .a(n_35735), .b(n_44174), .o(n_35822) );
ao22s80 FE_RC_228_0 ( .a(n_12827), .b(n_12593), .c(FE_OCP_RBN1132_n_12827), .d(n_12592), .o(n_13005) );
no02f80 g754804 ( .a(n_25401), .b(n_25358), .o(n_25402) );
no02f80 g768042 ( .a(n_12739), .b(n_12738), .o(n_12782) );
in01f80 newInst_147 ( .a(newNet_58), .o(newNet_147) );
na02f80 g766906 ( .a(n_13615), .b(n_13628), .o(n_13743) );
oa12f80 g753787 ( .a(n_26340), .b(n_26359), .c(n_26368), .o(n_26444) );
na02f80 g745255 ( .a(n_35656), .b(FE_OFN221_n_35655), .o(n_35657) );
na02f80 g738759 ( .a(n_41456), .b(n_41125), .o(n_41479) );
in01f80 g775787 ( .a(n_5128), .o(n_5129) );
in01f80 g773561 ( .a(n_7460), .o(n_7461) );
in01f80 g760689 ( .a(n_19724), .o(n_19744) );
in01f80 newInst_3356 ( .a(newNet_354), .o(newNet_3356) );
no02f80 g750684 ( .a(n_29236), .b(n_28788), .o(n_29353) );
na02f80 g754524 ( .a(n_26607), .b(FE_OCP_RBN2959_n_26231), .o(n_26687) );
na02f80 g758787 ( .a(n_21556), .b(n_21430), .o(n_21621) );
no02f80 g742862 ( .a(n_37445), .b(n_37164), .o(n_37270) );
in01f80 g737080 ( .a(n_43199), .o(n_43276) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_12_ ( .ck(newNet_754), .d(n_46167), .o(delay_xor_ln21_unr6_stage3_stallmux_q_12_) );
in01f80 newInst_2231 ( .a(newNet_1783), .o(newNet_2231) );
in01f80 FE_OCPUNCOC1803_n_18111 ( .a(n_18111), .o(FE_OCPUNCON1803_n_18111) );
in01f80 g774152 ( .a(n_7123), .o(n_7124) );
in01f80 g763713 ( .a(n_16690), .o(n_16736) );
in01f80 g766398 ( .a(n_14359), .o(n_14358) );
in01f80 FE_RC_1160_0 ( .a(n_41612), .o(FE_RN_349_0) );
in01f80 g767676 ( .a(n_13375), .o(n_13376) );
oa12f80 g771021 ( .a(n_9593), .b(n_9703), .c(n_9542), .o(n_9890) );
no02f80 g748688 ( .a(n_31163), .b(n_31141), .o(n_31166) );
na02f80 g753992 ( .a(n_26131), .b(n_26159), .o(n_26297) );
na02f80 g744403 ( .a(n_35471), .b(n_35468), .o(n_35532) );
in01f80 g776357 ( .a(n_4496), .o(n_4497) );
in01f80 g768913 ( .a(n_11927), .o(n_11833) );
in01f80 g775049 ( .a(n_6082), .o(n_6098) );
in01f80 FE_OCPC1506_n_17680 ( .a(FE_OCPN1505_n_17680), .o(FE_OCPN1506_n_17680) );
ao22s80 g736431 ( .a(n_43740), .b(n_43582), .c(n_43739), .d(n_43581), .o(n_43784) );
na02f80 g737008 ( .a(FE_OCP_RBN3067_n_43230), .b(n_43007), .o(n_43523) );
in01f80 newInst_2695 ( .a(newNet_829), .o(newNet_2695) );
in01f80 g777110 ( .a(n_3959), .o(n_3960) );
in01f80 g776364 ( .a(n_4727), .o(n_4728) );
no02f80 g775959 ( .a(n_5181), .b(n_4549), .o(n_5218) );
no02f80 g754441 ( .a(n_25726), .b(n_25512), .o(n_25753) );
na02f80 g754552 ( .a(n_26864), .b(n_26417), .o(n_26418) );
na02f80 g760226 ( .a(n_20249), .b(FE_OCP_RBN1352_n_19148), .o(n_20288) );
in01f80 g758990 ( .a(n_21644), .o(n_21575) );
in01f80 newInst_1679 ( .a(newNet_1678), .o(newNet_1679) );
in01f80 newInst_3139 ( .a(newNet_3138), .o(newNet_3139) );
na02f80 g745278 ( .a(n_36120), .b(n_36049), .o(n_36221) );
in01f80 newInst_359 ( .a(newNet_358), .o(newNet_359) );
no03m80 FE_RC_2512_0 ( .a(FE_RN_1022_0), .b(n_17929), .c(n_17998), .o(n_18021) );
in01f80 g775102 ( .a(n_6021), .o(n_6022) );
na02f80 g780052 ( .a(n_1238), .b(n_927), .o(n_1240) );
in01f80 g746062 ( .a(FE_OCP_DRV_N1578_n_33904), .o(n_33905) );
na02f80 g778195 ( .a(n_2699), .b(n_2698), .o(n_2700) );
no02f80 g770738 ( .a(n_11253), .b(FE_RN_1433_0), .o(n_10098) );
na02f80 FE_RC_2186_0 ( .a(FE_RN_781_0), .b(n_22750), .o(FE_RN_782_0) );
na02f80 g770760 ( .a(FE_OCP_RBN3652_n_10100), .b(n_9173), .o(n_10376) );
in01f80 g775090 ( .a(n_6009), .o(n_6010) );
oa12f80 g738257 ( .a(n_41871), .b(n_41870), .c(n_41869), .o(n_41949) );
in01f80 newInst_1900 ( .a(newNet_1713), .o(newNet_1900) );
no02f80 g755085 ( .a(n_25043), .b(n_24751), .o(n_25106) );
in01f80 g780655 ( .a(n_890), .o(n_923) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_18_ ( .ck(newNet_2005), .d(n_46986), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_18_) );
in01f80 g744292 ( .a(n_35856), .o(n_35974) );
no02f80 g762033 ( .a(FE_OCPN1776_n_18263), .b(n_18311), .o(n_18333) );
in01f80 newInst_3229 ( .a(newNet_3228), .o(newNet_3229) );
na02f80 g777352 ( .a(n_4675), .b(n_5168), .o(n_5287) );
in01f80 g776241 ( .a(n_4962), .o(n_4963) );
ao22s80 FE_RC_1348_0 ( .a(n_43012), .b(FE_OCP_RBN3033_n_43000), .c(delay_sub_ln23_0_unr30_stage10_stallmux_q), .d(n_43000), .o(n_43026) );
in01f80 g761635 ( .a(n_18971), .o(n_19127) );
na02f80 g781074 ( .a(sin_out_23), .b(FE_OFN3_n_43918), .o(n_289) );
na02f80 g769895 ( .a(n_10938), .b(n_10912), .o(n_11052) );
in01f80 g739751 ( .a(n_40528), .o(n_40529) );
oa22f80 g745643 ( .a(n_35451), .b(n_34962), .c(n_35452), .d(n_34963), .o(n_35525) );
in01f80 newInst_2821 ( .a(newNet_2820), .o(newNet_2821) );
oa12f80 g746443 ( .a(n_35018), .b(n_35017), .c(n_35016), .o(n_36111) );
in01f80 g748214 ( .a(n_32768), .o(n_32769) );
in01f80 g753964 ( .a(n_26251), .o(n_26252) );
na02f80 g744614 ( .a(n_35325), .b(n_33905), .o(n_35375) );
oa12f80 g736522 ( .a(n_43477), .b(n_43661), .c(n_43275), .o(n_43722) );
na02f80 g776224 ( .a(n_4830), .b(n_4516), .o(n_4876) );
no02f80 g745414 ( .a(FE_OCP_RBN2986_n_35539), .b(n_35633), .o(n_36055) );
na02f80 g754910 ( .a(n_25481), .b(n_24794), .o(n_25626) );
oa22f80 g771516 ( .a(n_9042), .b(n_9030), .c(FE_OCP_RBN2650_n_9042), .d(FE_OCP_RBN2651_n_9030), .o(n_9247) );
in01f80 FE_RC_2979_0 ( .a(n_29451), .o(FE_RN_1301_0) );
in01f80 g770249 ( .a(n_10891), .o(n_10979) );
na02f80 g740896 ( .a(n_39146), .b(n_39060), .o(n_39168) );
in01f80 g740633 ( .a(n_39633), .o(n_39634) );
no02f80 g761017 ( .a(n_19204), .b(n_18032), .o(n_19252) );
na02f80 g769122 ( .a(n_11621), .b(n_11557), .o(n_11745) );
in01f80 g745887 ( .a(n_34094), .o(n_34139) );
oa12f80 g778013 ( .a(n_2986), .b(n_3008), .c(n_2985), .o(n_4298) );
na02f80 g740962 ( .a(n_39086), .b(n_38879), .o(n_39110) );
ao12f80 g774196 ( .a(n_7097), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .o(n_7154) );
in01f80 g780314 ( .a(n_991), .o(n_992) );
na02f80 g774145 ( .a(n_6818), .b(n_6844), .o(n_6866) );
in01f80 g772464 ( .a(n_8413), .o(n_8414) );
in01f80 g779872 ( .a(n_1285), .o(n_1286) );
na02f80 g741029 ( .a(n_39010), .b(n_39009), .o(n_39011) );
in01f80 g738707 ( .a(n_41577), .o(n_41487) );
in01f80 g751259 ( .a(n_29800), .o(n_29818) );
no02f80 g773438 ( .a(n_7533), .b(n_6704), .o(n_7603) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_15_ ( .ck(newNet_1422), .d(n_36542), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_) );
in01f80 FE_OCP_RBC3729_n_43230 ( .a(FE_OCP_RBN3068_n_43230), .o(FE_OCP_RBN3729_n_43230) );
oa22f80 FE_RC_2730_0 ( .a(n_27827), .b(n_27831), .c(n_27828), .d(n_27832), .o(n_27939) );
in01f80 g746450 ( .a(n_33346), .o(n_33347) );
in01f80 FE_RC_1134_0 ( .a(n_2746), .o(FE_RN_342_0) );
no02f80 g777175 ( .a(n_4675), .b(n_5166), .o(n_5191) );
in01f80 newInst_3579 ( .a(newNet_3578), .o(newNet_3579) );
in01f80 newInst_226 ( .a(newNet_173), .o(newNet_226) );
na02f80 g747832 ( .a(n_33392), .b(n_33554), .o(n_33600) );
in01f80 newInst_1167 ( .a(newNet_1067), .o(newNet_1167) );
na02f80 g756721 ( .a(n_23539), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_14_), .o(n_23635) );
na02f80 g749210 ( .a(n_30683), .b(n_30713), .o(n_30862) );
in01f80 newInst_232 ( .a(newNet_231), .o(newNet_232) );
in01f80 g741239 ( .a(n_38880), .o(n_38881) );
in01f80 FE_RC_2026_0 ( .a(n_23271), .o(FE_RN_674_0) );
no02f80 g773498 ( .a(n_7462), .b(n_7292), .o(n_7490) );
na02f80 g744747 ( .a(n_36495), .b(n_35936), .o(n_36555) );
in01f80 FE_RC_4212_0 ( .a(n_19976), .o(n_19970) );
oa12f80 g738356 ( .a(n_41519), .b(n_41518), .c(n_41517), .o(n_42188) );
na02f80 g737540 ( .a(n_42290), .b(n_42262), .o(n_42291) );
in01f80 FE_RC_68_0 ( .a(n_17661), .o(FE_RN_18_0) );
no02f80 g777363 ( .a(n_3637), .b(n_3663), .o(n_3665) );
in01f80 newInst_830 ( .a(newNet_829), .o(newNet_830) );
ao12f80 g762889 ( .a(n_17655), .b(n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_8_), .o(n_17726) );
in01f80 newInst_1820 ( .a(newNet_1819), .o(newNet_1820) );
na02f80 g738519 ( .a(n_41582), .b(n_41695), .o(n_41748) );
in01f80 g746191 ( .a(n_33895), .o(n_33896) );
oa22f80 g748028 ( .a(n_44346), .b(n_32530), .c(n_44347), .d(n_32531), .o(n_33336) );
oa22f80 FE_RC_3030_0 ( .a(delay_sub_ln23_0_unr23_stage8_stallmux_q), .b(n_36709), .c(n_36654), .d(n_36750), .o(n_36722) );
in01f80 g759352 ( .a(n_21147), .o(n_21175) );
in01f80 newInst_1160 ( .a(newNet_1159), .o(newNet_1160) );
no02f80 g772697 ( .a(n_8267), .b(n_8258), .o(n_8364) );
in01f80 g770270 ( .a(n_10772), .o(n_10773) );
in01f80 newInst_1169 ( .a(newNet_1168), .o(newNet_1169) );
na02f80 g781141 ( .a(n_205), .b(n_207), .o(n_214) );
ao22s80 g743721 ( .a(n_37329), .b(n_46245), .c(n_37328), .d(n_36849), .o(n_37473) );
no02f80 FE_RC_1636_0 ( .a(FE_RN_453_0), .b(FE_RN_454_0), .o(FE_RN_455_0) );
oa22f80 FE_RC_2680_0 ( .a(n_2973), .b(n_4132), .c(n_2974), .d(n_4184), .o(n_4396) );
in01f80 g737186 ( .a(n_42998), .o(n_43009) );
na02f80 g758304 ( .a(n_22288), .b(n_20978), .o(n_22404) );
in01f80 g738213 ( .a(n_41962), .o(n_41974) );
no02f80 FE_RC_1913_0 ( .a(n_18950), .b(FE_RN_601_0), .o(n_19058) );
no02f80 g755095 ( .a(n_25268), .b(n_25204), .o(n_25460) );
oa12f80 g742950 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(n_37110), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n_37271) );
in01f80 newInst_3165 ( .a(newNet_3164), .o(newNet_3165) );
no03m80 g743395 ( .a(n_37750), .b(n_37785), .c(n_37749), .o(n_37825) );
oa12f80 g760592 ( .a(n_19502), .b(n_19728), .c(n_19552), .o(n_19818) );
in01f80 newInst_2475 ( .a(newNet_2474), .o(newNet_2475) );
no02f80 g768071 ( .a(n_12709), .b(n_12692), .o(n_12748) );
no02f80 g779327 ( .a(n_1708), .b(n_1707), .o(n_1709) );
no02f80 g766379 ( .a(FE_OCP_RBN2455_n_14157), .b(n_14274), .o(n_14276) );
in01f80 g737942 ( .a(n_42343), .o(n_42344) );
na02f80 g739438 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_18_), .o(n_40766) );
in01f80 g750323 ( .a(n_29689), .o(n_29690) );
no02f80 g775144 ( .a(n_6015), .b(n_5850), .o(n_6036) );
in01f80 g755069 ( .a(n_25477), .o(n_25478) );
in01f80 g752275 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .o(n_27806) );
in01f80 newInst_1272 ( .a(newNet_1271), .o(newNet_1272) );
oa12f80 g773574 ( .a(n_7421), .b(n_7420), .c(n_7419), .o(n_7468) );
in01f80 g738182 ( .a(n_42011), .o(n_42012) );
na02f80 g746557 ( .a(n_35041), .b(n_34549), .o(n_35086) );
in01f80 newInst_1077 ( .a(newNet_1040), .o(newNet_1077) );
no02f80 g772493 ( .a(n_8462), .b(FE_OCP_RBN3466_n_7886), .o(n_8463) );
in01f80 newInst_2797 ( .a(newNet_2796), .o(newNet_2797) );
ao22s80 g780350 ( .a(n_1122), .b(n_789), .c(n_1208), .d(n_856), .o(n_899) );
in01f80 g748847 ( .a(n_31056), .o(n_31057) );
in01f80 g777016 ( .a(n_3853), .o(n_3854) );
ao12f80 g773044 ( .a(n_7730), .b(n_7763), .c(n_7828), .o(n_7818) );
no02f80 g755982 ( .a(n_24184), .b(n_23769), .o(n_24251) );
in01f80 newInst_727 ( .a(newNet_174), .o(newNet_727) );
oa12f80 g737536 ( .a(n_42268), .b(n_42265), .c(FE_OCPN936_n_42192), .o(n_42532) );
na02f80 g745183 ( .a(n_36230), .b(n_35604), .o(n_36056) );
oa12f80 g758731 ( .a(FE_OCP_RBN2952_n_21489), .b(n_21805), .c(n_21490), .o(n_21895) );
ao12f80 g746760 ( .a(n_33108), .b(n_33107), .c(n_32222), .o(n_33109) );
na02f80 g768554 ( .a(n_12327), .b(FE_OCPN1002_n_45660), .o(n_12371) );
in01f80 FE_OCPC1782_FE_OCP_RBN1701_n_19353 ( .a(FE_OCPN1781_FE_OCP_RBN1701_n_19353), .o(FE_OCPN1782_FE_OCP_RBN1701_n_19353) );
no02f80 g780910 ( .a(n_377), .b(n_398), .o(n_404) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_22_ ( .ck(newNet_1225), .d(n_6042), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_22_) );
ao12f80 g766848 ( .a(n_13741), .b(n_13740), .c(n_13739), .o(n_15686) );
in01f80 newInst_2686 ( .a(newNet_316), .o(newNet_2686) );
oa12f80 g757612 ( .a(n_22633), .b(n_22632), .c(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_), .o(n_24097) );
in01f80 g736341 ( .a(n_43831), .o(n_43832) );
in01f80 FE_RC_3865_0 ( .a(FE_RN_1689_0), .o(n_22496) );
na02f80 FE_RC_2511_0 ( .a(FE_RN_1020_0), .b(FE_RN_1021_0), .o(FE_RN_1022_0) );
in01f80 g769237 ( .a(n_12429), .o(n_12430) );
ao12f80 g779644 ( .a(n_1431), .b(n_1452), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_28_), .o(n_1487) );
no02f80 g771404 ( .a(n_9167), .b(n_8905), .o(n_9293) );
oa22f80 g749477 ( .a(n_31886), .b(n_31564), .c(n_31885), .d(n_31565), .o(n_31960) );
no02f80 g753950 ( .a(n_26190), .b(n_23447), .o(n_26219) );
no02f80 g736625 ( .a(n_43193), .b(n_43067), .o(n_43238) );
in01f80 g750751 ( .a(n_29368), .o(n_29369) );
na02f80 g774306 ( .a(n_6938), .b(n_6879), .o(n_6976) );
in01f80 g739370 ( .a(n_40949), .o(n_40950) );
ao22s80 g762630 ( .a(n_17914), .b(n_17916), .c(n_17998), .d(n_17915), .o(n_18049) );
no02f80 g748152 ( .a(n_31902), .b(FE_OCP_RBN1213_n_31847), .o(n_31988) );
in01f80 g747120 ( .a(n_32788), .o(n_32789) );
in01f80 g779260 ( .a(n_1820), .o(n_1821) );
in01f80 g762055 ( .a(n_18248), .o(n_18203) );
na02f80 g766326 ( .a(n_14133), .b(n_14117), .o(n_14245) );
na02f80 FE_RC_43_0 ( .a(FE_RN_9_0), .b(FE_RN_10_0), .o(FE_RN_11_0) );
no02f80 FE_RC_3819_0 ( .a(FE_RN_1238_0), .b(FE_RN_1666_0), .o(n_24684) );
na02f80 g741832 ( .a(n_38366), .b(n_38365), .o(n_38367) );
in01f80 g765161 ( .a(n_15276), .o(n_15308) );
in01f80 newInst_1242 ( .a(newNet_1241), .o(newNet_1242) );
in01f80 fopt783796 ( .a(n_45474), .o(n_45475) );
na02f80 g778149 ( .a(n_2932), .b(n_2743), .o(n_2987) );
no02f80 g775719 ( .a(n_5221), .b(n_4182), .o(n_5256) );
oa12f80 g753292 ( .a(n_27627), .b(n_27657), .c(n_26896), .o(n_27677) );
na02f80 g771226 ( .a(n_9448), .b(FE_OCP_RBN2554_n_44576), .o(n_9593) );
no02f80 g773939 ( .a(n_6994), .b(n_7000), .o(n_6995) );
no02f80 g758218 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .o(n_22850) );
in01f80 newInst_2111 ( .a(newNet_2110), .o(newNet_2111) );
no02f80 g751515 ( .a(n_29177), .b(n_28906), .o(n_29175) );
in01f80 g763899 ( .a(n_17421), .o(n_17100) );
no02f80 g757818 ( .a(FE_OCP_RBN1920_n_22476), .b(n_22554), .o(n_22555) );
in01f80 g738528 ( .a(n_41580), .o(n_41581) );
oa12f80 g777942 ( .a(n_2265), .b(n_3092), .c(n_2244), .o(n_3147) );
no02f80 g742635 ( .a(n_37525), .b(n_37524), .o(n_37526) );
na02f80 FE_RC_652_0 ( .a(FE_RN_207_0), .b(FE_RN_208_0), .o(FE_RN_209_0) );
ao12f80 g754473 ( .a(n_25292), .b(n_25544), .c(n_25206), .o(n_25600) );
in01f80 g771112 ( .a(n_9724), .o(n_9796) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_23_ ( .ck(newNet_1224), .d(n_6159), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_) );
in01f80 g773676 ( .a(n_7365), .o(n_7366) );
no02f80 g743867 ( .a(n_36011), .b(n_36100), .o(n_36102) );
na02f80 FE_RC_3050_0 ( .a(FE_RN_1334_0), .b(FE_RN_1335_0), .o(FE_RN_1336_0) );
in01f80 newInst_3026 ( .a(newNet_3025), .o(newNet_3026) );
ao12f80 g757104 ( .a(n_23378), .b(n_44068), .c(delay_xor_ln22_unr15_stage6_stallmux_q_12_), .o(n_23178) );
oa12f80 g743903 ( .a(n_35484), .b(n_35538), .c(n_35502), .o(n_35627) );
no02f80 g766051 ( .a(n_14608), .b(n_14506), .o(n_14663) );
na02f80 g764687 ( .a(n_15895), .b(n_15736), .o(n_15943) );
in01f80 newInst_2665 ( .a(newNet_1184), .o(newNet_2665) );
oa22f80 FE_RC_2205_0 ( .a(n_27526), .b(n_27675), .c(n_27525), .d(n_27697), .o(n_27785) );
in01f80 g737227 ( .a(n_43002), .o(n_42982) );
in01f80 newInst_1582 ( .a(newNet_452), .o(newNet_1582) );
in01f80 g781317 ( .a(n_56), .o(n_106) );
na02f80 g776781 ( .a(n_3994), .b(n_3788), .o(n_4105) );
in01f80 g745878 ( .a(n_34067), .o(n_34068) );
na02f80 g739175 ( .a(n_40894), .b(n_40855), .o(n_40942) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_18_ ( .ck(newNet_1528), .d(n_32247), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_18_) );
in01f80 g767712 ( .a(n_13363), .o(n_13364) );
in01f80 g763784 ( .a(n_46976), .o(n_16774) );
na02f80 FE_RC_2851_0 ( .a(FE_RN_1227_0), .b(n_19770), .o(n_19854) );
no02f80 g779531 ( .a(n_1445), .b(n_1470), .o(n_1746) );
ao12f80 g779472 ( .a(n_1882), .b(n_1852), .c(delay_xor_ln21_unr3_stage2_stallmux_q_18_), .o(n_1931) );
in01f80 g739465 ( .a(n_41077), .o(n_41078) );
in01f80 newInst_3147 ( .a(newNet_2059), .o(newNet_3147) );
no02f80 g777818 ( .a(n_3292), .b(n_3271), .o(n_3375) );
in01f80 g751075 ( .a(n_30124), .o(n_30125) );
no02f80 g743037 ( .a(n_37098), .b(n_37097), .o(n_37482) );
ao12f80 g763031 ( .a(n_17504), .b(n_17635), .c(n_17580), .o(n_17717) );
na02f80 g765928 ( .a(n_14726), .b(n_45519), .o(n_14818) );
in01f80 newInst_3728 ( .a(newNet_3138), .o(newNet_3728) );
no02f80 g752197 ( .a(n_28009), .b(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n_27973) );
no02f80 g750500 ( .a(n_29507), .b(FE_OCPN1464_n_29630), .o(n_29508) );
in01f80 FE_OCP_RBC3564_n_29857 ( .a(n_29857), .o(FE_OCP_RBN3564_n_29857) );
no02f80 g764920 ( .a(n_15357), .b(FE_OCPN1257_n_13831), .o(n_15358) );
in01f80 newInst_1910 ( .a(newNet_1909), .o(newNet_1910) );
na02f80 g753268 ( .a(n_27287), .b(n_25980), .o(n_27329) );
oa12f80 g773693 ( .a(n_7357), .b(n_8174), .c(n_7364), .o(n_9331) );
ao22s80 g781178 ( .a(n_174), .b(n_124), .c(n_171), .d(n_123), .o(n_368) );
no02f80 g739006 ( .a(n_41192), .b(n_41183), .o(n_41184) );
na02f80 g739605 ( .a(n_40614), .b(n_44610), .o(n_40654) );
na02f80 g745215 ( .a(n_36125), .b(n_35995), .o(n_36228) );
na02f80 g770813 ( .a(n_10051), .b(n_10107), .o(n_10176) );
na03f80 g784624 ( .a(n_36385), .b(n_35795), .c(n_35717), .o(n_46953) );
no02f80 g774520 ( .a(FE_OCPN895_n_6521), .b(n_6473), .o(n_6828) );
na02f80 g749864 ( .a(FE_OCP_RBN3011_n_31117), .b(n_31210), .o(n_31571) );
in01f80 g759197 ( .a(n_21346), .o(n_22156) );
in01f80 g737852 ( .a(n_42691), .o(n_42692) );
na02f80 g752031 ( .a(n_28042), .b(n_28003), .o(n_28101) );
in01f80 g761573 ( .a(n_20086), .o(n_20231) );
in01f80 FE_OCP_RBC1193_n_22542 ( .a(n_22542), .o(FE_OCP_RBN1193_n_22542) );
in01f80 newInst_2070 ( .a(newNet_2069), .o(newNet_2070) );
in01f80 g736595 ( .a(n_43417), .o(n_43446) );
in01f80 newInst_3253 ( .a(newNet_3252), .o(newNet_3253) );
no02f80 g778081 ( .a(n_2892), .b(n_2925), .o(n_4587) );
ao12f80 g772757 ( .a(n_7368), .b(n_7905), .c(n_7403), .o(n_7986) );
in01f80 g752541 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_17_), .o(n_27712) );
oa12f80 g765914 ( .a(n_14870), .b(n_14898), .c(n_14869), .o(n_14972) );
no02f80 g773469 ( .a(n_7516), .b(n_7515), .o(n_7551) );
oa12f80 g752207 ( .a(n_28005), .b(FE_OCP_RBN2126_n_44734), .c(delay_xor_ln21_unr18_stage7_stallmux_q_13_), .o(n_28033) );
in01f80 newInst_1596 ( .a(newNet_1595), .o(newNet_1596) );
no02f80 g773977 ( .a(n_7217), .b(delay_xor_ln22_unr6_stage3_stallmux_q_23_), .o(n_7257) );
na02f80 g737017 ( .a(n_43230), .b(n_42666), .o(n_43492) );
ao12f80 g748837 ( .a(n_32445), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_), .o(n_33124) );
in01f80 g758765 ( .a(n_22247), .o(n_22248) );
in01f80 newInst_773 ( .a(newNet_772), .o(newNet_773) );
in01f80 g741230 ( .a(n_39176), .o(n_39177) );
no02f80 g779637 ( .a(n_1409), .b(n_1484), .o(n_2013) );
in01f80 FE_OCP_RBC1148_n_27966 ( .a(n_27966), .o(FE_OCP_RBN1148_n_27966) );
in01f80 g751464 ( .a(n_28849), .o(n_28850) );
in01f80 newInst_2552 ( .a(newNet_2551), .o(newNet_2552) );
ao22s80 FE_RC_330_0 ( .a(n_44364), .b(n_22462), .c(n_22464), .d(n_22705), .o(n_22790) );
in01f80 g774935 ( .a(n_6209), .o(n_6210) );
in01f80 FE_OCP_RBC3001_n_42959 ( .a(n_42959), .o(FE_OCP_RBN3001_n_42959) );
na02f80 g749322 ( .a(n_30817), .b(n_30791), .o(n_30865) );
in01f80 newInst_2535 ( .a(newNet_2534), .o(newNet_2535) );
no02f80 g738358 ( .a(n_41455), .b(n_41410), .o(n_41476) );
ao12f80 FE_RC_2817_0 ( .a(FE_RN_1206_0), .b(n_34423), .c(n_34908), .o(n_35005) );
in01f80 newInst_3265 ( .a(newNet_1062), .o(newNet_3265) );
na02f80 g772615 ( .a(n_8283), .b(n_7859), .o(n_8337) );
in01f80 g742481 ( .a(n_37649), .o(n_38047) );
in01f80 newInst_2629 ( .a(newNet_2628), .o(newNet_2629) );
in01f80 FE_OCP_RBC1923_cordic_combinational_sub_ln23_0_unr12_z_0__ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN1923_cordic_combinational_sub_ln23_0_unr12_z_0__) );
na02f80 g757011 ( .a(n_23305), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_8_), .o(n_23373) );
in01f80 g749646 ( .a(n_30180), .o(n_30250) );
in01f80 g739211 ( .a(n_40743), .o(n_40744) );
in01f80 newInst_2255 ( .a(newNet_2254), .o(newNet_2255) );
na02f80 g774815 ( .a(n_6312), .b(n_6171), .o(n_6360) );
na02f80 g739180 ( .a(n_40801), .b(n_40799), .o(n_40800) );
in01f80 FE_OCP_RBC2395_n_8288 ( .a(FE_OCP_RBN2394_n_8288), .o(FE_OCP_RBN2395_n_8288) );
ao12f80 g759258 ( .a(n_21374), .b(n_21755), .c(n_21835), .o(n_21836) );
no02f80 FE_RC_2070_0 ( .a(n_24924), .b(FE_RN_704_0), .o(FE_RN_705_0) );
na02f80 g762929 ( .a(n_17987), .b(n_17986), .o(n_17988) );
na02f80 g763177 ( .a(n_17047), .b(n_17091), .o(n_17250) );
in01f80 FE_OCP_RBC2387_n_13860 ( .a(n_13860), .o(FE_OCP_RBN2387_n_13860) );
na02f80 FE_RC_2433_0 ( .a(FE_RN_967_0), .b(FE_RN_968_0), .o(FE_RN_969_0) );
no02f80 g763735 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_), .o(n_17605) );
na02f80 g772993 ( .a(n_7777), .b(n_7746), .o(n_7875) );
na02f80 g751187 ( .a(n_29800), .b(n_28928), .o(n_29854) );
in01f80 g736861 ( .a(n_43613), .o(n_43614) );
no02f80 g755457 ( .a(n_24802), .b(n_24696), .o(n_24823) );
in01f80 newInst_455 ( .a(newNet_454), .o(newNet_455) );
na02f80 g778695 ( .a(n_2438), .b(FE_OFN813_n_2540), .o(n_2571) );
na02f80 g776373 ( .a(n_4646), .b(n_3645), .o(n_4750) );
na02f80 g749028 ( .a(n_30960), .b(n_27131), .o(n_31007) );
no02f80 g767291 ( .a(n_13680), .b(n_13679), .o(n_13681) );
na02f80 g740447 ( .a(n_39719), .b(n_39687), .o(n_39720) );
na02f80 g756373 ( .a(n_24301), .b(n_24300), .o(n_24302) );
in01f80 FE_RC_1957_0 ( .a(n_14321), .o(FE_RN_630_0) );
no02f80 g772955 ( .a(n_8550), .b(n_7995), .o(n_8105) );
na02f80 g742590 ( .a(n_37572), .b(n_37571), .o(n_37573) );
na02f80 g741658 ( .a(n_38540), .b(n_38240), .o(n_38575) );
in01f80 FE_OCP_RBC2390_n_19434 ( .a(n_19434), .o(FE_OCP_RBN2390_n_19434) );
ao12f80 g757272 ( .a(n_23022), .b(n_44068), .c(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .o(n_23045) );
oa12f80 g736301 ( .a(n_292), .b(n_43868), .c(FE_OFN1_n_43918), .o(n_43897) );
oa22f80 g736912 ( .a(n_43230), .b(n_42936), .c(FE_OCP_RBN3729_n_43230), .d(n_46940), .o(n_43630) );
oa22f80 FE_RC_2835_0 ( .a(n_15671), .b(n_15818), .c(n_15672), .d(n_15819), .o(n_16011) );
in01f80 g752568 ( .a(n_27691), .o(n_27659) );
in01f80 g764992 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_3_), .o(n_17496) );
ms00f80 delay_sub_ln23_0_unr1_stage2_stallmux_q_reg_0_ ( .ck(newNet_1665), .d(n_50), .o(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_) );
in01f80 FE_OCP_RBC2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
ao12f80 g754961 ( .a(n_25153), .b(n_25152), .c(n_25151), .o(n_26820) );
in01f80 newInst_820 ( .a(newNet_819), .o(newNet_820) );
in01f80 FE_OCPC1744_n_24962 ( .a(FE_OCPN1743_n_24962), .o(FE_OCPN1744_n_24962) );
in01f80 newInst_3736 ( .a(newNet_3735), .o(newNet_3736) );
na02f80 g760947 ( .a(n_19357), .b(n_19332), .o(n_19453) );
in01f80 newInst_1788 ( .a(newNet_1601), .o(newNet_1788) );
in01f80 g745039 ( .a(n_34924), .o(n_34925) );
no02f80 g750699 ( .a(n_29392), .b(n_29391), .o(n_29465) );
in01f80 newInst_2198 ( .a(newNet_2197), .o(newNet_2198) );
na02f80 g776017 ( .a(n_5061), .b(n_5009), .o(n_5036) );
na02f80 g740214 ( .a(n_39893), .b(n_39942), .o(n_39943) );
in01f80 g777594 ( .a(n_3817), .o(n_3819) );
in01f80 g765711 ( .a(FE_OFN767_n_15670), .o(n_17753) );
in01f80 g761059 ( .a(n_21454), .o(n_20179) );
no02f80 g747955 ( .a(n_33072), .b(n_32561), .o(n_33087) );
no02f80 g756296 ( .a(n_24068), .b(n_24067), .o(n_24069) );
na02f80 g745833 ( .a(n_44102), .b(n_33750), .o(n_34258) );
no02f80 g763202 ( .a(FE_OCP_RBN3689_n_16146), .b(n_17195), .o(n_17248) );
na02f80 g780839 ( .a(n_461), .b(n_444), .o(n_462) );
in01f80 g737491 ( .a(n_42564), .o(n_42565) );
no02f80 g763429 ( .a(n_16839), .b(n_15651), .o(n_16882) );
in01f80 g766254 ( .a(n_14462), .o(n_14463) );
no02f80 g763246 ( .a(n_17006), .b(n_16998), .o(n_17249) );
na02f80 g784703 ( .a(n_47177), .b(FE_RN_968_0), .o(n_47179) );
na02f80 g754241 ( .a(n_25939), .b(n_25881), .o(n_25964) );
no02f80 g760791 ( .a(n_19480), .b(n_18705), .o(n_19539) );
no02f80 g738060 ( .a(n_42089), .b(n_41903), .o(n_42110) );
na02f80 g760437 ( .a(n_20655), .b(n_20013), .o(n_20739) );
na02f80 g766553 ( .a(n_14115), .b(n_14140), .o(n_14172) );
oa22f80 g753744 ( .a(n_27080), .b(n_26893), .c(n_27079), .d(n_26892), .o(n_27134) );
no02f80 g757455 ( .a(FE_OCP_RBN3823_n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_4_), .o(n_22869) );
na02f80 g757287 ( .a(n_23188), .b(n_23128), .o(n_23206) );
na02f80 g777656 ( .a(n_3568), .b(n_3536), .o(n_3623) );
na02f80 g772673 ( .a(n_8299), .b(n_8270), .o(n_8390) );
na02f80 g746543 ( .a(n_34499), .b(n_34498), .o(n_34525) );
oa12f80 g766561 ( .a(n_46415), .b(n_13866), .c(n_13138), .o(n_13928) );
in01f80 g757684 ( .a(n_22790), .o(n_22857) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_7_ ( .ck(newNet_207), .d(n_46143), .o(delay_xor_ln22_unr6_stage3_stallmux_q_7_) );
oa22f80 FE_RC_4111_0 ( .a(n_32122), .b(n_32360), .c(n_44213), .d(n_32123), .o(n_32516) );
na02f80 g767275 ( .a(n_13489), .b(n_12914), .o(n_13530) );
ao12f80 g780420 ( .a(n_884), .b(n_820), .c(n_799), .o(n_885) );
in01f80 g777285 ( .a(n_5091), .o(n_4884) );
oa22f80 g773692 ( .a(n_7321), .b(n_6730), .c(n_8135), .d(n_7286), .o(n_9391) );
in01f80 g749787 ( .a(n_31315), .o(n_31316) );
in01f80 FE_OFC762_n_15670 ( .a(n_15670), .o(FE_OFN762_n_15670) );
in01f80 g740845 ( .a(n_39293), .o(n_39314) );
no02f80 g745998 ( .a(n_33977), .b(n_33975), .o(n_34011) );
in01f80 FE_OCP_RBC2688_n_38870 ( .a(FE_OCP_RBN3625_n_38870), .o(FE_OCP_RBN2688_n_38870) );
in01f80 g741136 ( .a(n_39423), .o(n_39424) );
in01f80 g744513 ( .a(n_35423), .o(n_35424) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_10_ ( .ck(newNet_275), .d(n_46158), .o(delay_xor_ln22_unr6_stage3_stallmux_q_10_) );
na02f80 FE_RC_3634_0 ( .a(n_31795), .b(n_30350), .o(FE_RN_1593_0) );
na02f80 g781001 ( .a(n_279), .b(n_278), .o(n_280) );
oa12f80 g779194 ( .a(n_1851), .b(n_1862), .c(n_1850), .o(n_1915) );
na02f80 g750099 ( .a(n_29857), .b(n_29031), .o(n_29985) );
no02f80 g764910 ( .a(n_15552), .b(n_14452), .o(n_15554) );
na02f80 g750977 ( .a(n_29947), .b(FE_OCP_RBN2561_n_29819), .o(n_30039) );
in01f80 FE_OCP_DRV_C1592_n_34327 ( .a(FE_OCP_DRV_N1591_n_34327), .o(FE_OCP_DRV_N1592_n_34327) );
in01f80 g765394 ( .a(n_15369), .o(n_15370) );
in01f80 FE_RC_4065_0 ( .a(n_26564), .o(FE_RN_1769_0) );
na02f80 g766936 ( .a(n_14258), .b(n_14386), .o(n_14992) );
ao22s80 g736504 ( .a(n_43710), .b(n_43261), .c(n_43709), .d(n_43262), .o(n_43737) );
na02f80 FE_RC_2565_0 ( .a(n_34242), .b(n_34241), .o(FE_RN_1053_0) );
oa12f80 g755912 ( .a(n_25163), .b(n_25160), .c(n_25133), .o(n_25772) );
na02f80 g758914 ( .a(n_21291), .b(n_21328), .o(n_21475) );
oa22f80 g758703 ( .a(n_22242), .b(n_21857), .c(n_22243), .d(n_21858), .o(n_22362) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_8_ ( .ck(newNet_391), .d(n_32571), .o(delay_xor_ln22_unr21_stage8_stallmux_q_8_) );
in01f80 newInst_1554 ( .a(newNet_1553), .o(newNet_1554) );
na02f80 g766650 ( .a(FE_OCP_RBN2387_n_13860), .b(n_13916), .o(n_13917) );
in01f80 g738553 ( .a(n_41541), .o(n_41574) );
in01f80 newInst_1181 ( .a(newNet_201), .o(newNet_1181) );
in01f80 FE_OCP_RBC3802_n_44721 ( .a(n_44721), .o(FE_OCP_RBN3802_n_44721) );
na02f80 g768556 ( .a(n_12235), .b(n_11867), .o(n_12298) );
na02f80 g774502 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .o(n_6591) );
in01f80 g738891 ( .a(n_41302), .o(n_41319) );
no02f80 g744516 ( .a(n_35399), .b(n_35304), .o(n_35412) );
in01f80 g759727 ( .a(n_20477), .o(n_20478) );
no02f80 g741864 ( .a(n_38286), .b(n_38166), .o(n_38386) );
in01f80 g740513 ( .a(n_39756), .o(n_39757) );
in01f80 g781083 ( .a(n_259), .o(n_272) );
in01f80 newInst_1714 ( .a(newNet_344), .o(newNet_1714) );
no02f80 g779551 ( .a(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .o(n_1503) );
in01f80 g773403 ( .a(n_7569), .o(n_7577) );
no02f80 g744066 ( .a(n_44222), .b(n_35905), .o(n_35984) );
in01f80 g766860 ( .a(n_13659), .o(n_13673) );
na02f80 g765969 ( .a(n_15090), .b(n_14385), .o(n_15088) );
oa12f80 g748989 ( .a(n_31458), .b(n_32295), .c(n_31483), .o(n_32314) );
oa12f80 g736252 ( .a(n_294), .b(n_43911), .c(FE_OFN4_n_43918), .o(n_43919) );
in01f80 g760136 ( .a(n_20491), .o(n_20492) );
ao12f80 g766696 ( .a(n_13788), .b(n_13836), .c(n_13634), .o(n_13886) );
in01f80 newInst_2852 ( .a(newNet_2851), .o(newNet_2852) );
ao22s80 g780438 ( .a(FE_OFN795_n_45813), .b(n_923), .c(n_1203), .d(n_890), .o(n_1068) );
na02f80 g742044 ( .a(n_38137), .b(n_46416), .o(n_38201) );
na02f80 g764314 ( .a(n_16398), .b(n_14805), .o(n_16429) );
in01f80 g764609 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_9_), .o(n_17931) );
in01f80 newInst_1719 ( .a(newNet_1718), .o(newNet_1719) );
na02f80 g743197 ( .a(n_36908), .b(n_36884), .o(n_36932) );
in01f80 newInst_1777 ( .a(newNet_1776), .o(newNet_1777) );
na02f80 g750780 ( .a(n_29230), .b(n_29292), .o(n_29293) );
na02f80 g771564 ( .a(n_9076), .b(n_9201), .o(n_9202) );
in01f80 FE_OCP_RBC2714_n_14982 ( .a(n_14982), .o(FE_OCP_RBN2714_n_14982) );
na02f80 g751750 ( .a(n_28307), .b(n_28295), .o(n_28366) );
in01f80 g740772 ( .a(n_39905), .o(n_39562) );
in01f80 g755996 ( .a(n_25570), .o(n_25571) );
in01f80 g772314 ( .a(n_8608), .o(n_8609) );
na02f80 g763798 ( .a(n_16799), .b(delay_add_ln22_unr11_stage5_stallmux_q_0_), .o(n_17226) );
in01f80 newInst_910 ( .a(newNet_198), .o(newNet_910) );
na02f80 g770689 ( .a(n_10353), .b(n_10288), .o(n_10289) );
in01f80 g774535 ( .a(n_6513), .o(n_6514) );
no02f80 g736948 ( .a(FE_OCPN912_n_43022), .b(n_43211), .o(n_43255) );
oa12f80 g762297 ( .a(n_17999), .b(n_18080), .c(n_17952), .o(n_18138) );
ms00f80 delay_sub_ln23_unr25_stage8_stallmux_q_reg_1_ ( .ck(newNet_1047), .d(n_32292), .o(delay_sub_ln23_unr25_stage8_stallmux_q_1_) );
in01f80 g764118 ( .a(n_16962), .o(n_16963) );
na02f80 g753870 ( .a(n_26301), .b(n_26258), .o(n_26332) );
oa22f80 FE_RC_3197_0 ( .a(n_6639), .b(n_6665), .c(n_6640), .d(n_6666), .o(n_6832) );
in01f80 g765092 ( .a(n_15580), .o(n_15490) );
na02f80 g757335 ( .a(n_22968), .b(n_23019), .o(n_23072) );
oa12f80 g762895 ( .a(n_17329), .b(n_17494), .c(n_17325), .o(n_17627) );
no02f80 g748065 ( .a(n_31994), .b(FE_OCP_RBN1214_n_31847), .o(n_32028) );
na02f80 g777089 ( .a(n_3805), .b(FE_OCP_RBN2580_n_3734), .o(n_3958) );
oa22f80 g752369 ( .a(n_28397), .b(n_28277), .c(n_28398), .d(n_28276), .o(n_28901) );
in01f80 FE_RC_836_0 ( .a(n_9271), .o(FE_RN_250_0) );
no02f80 g770008 ( .a(n_10800), .b(n_10793), .o(n_10915) );
in01f80 g776485 ( .a(n_4585), .o(n_4586) );
na02f80 g745970 ( .a(n_33906), .b(n_34590), .o(n_33944) );
in01f80 g757083 ( .a(n_23303), .o(n_23304) );
na02f80 g771830 ( .a(n_9874), .b(n_9873), .o(n_9875) );
na02f80 g750886 ( .a(n_29020), .b(n_28682), .o(n_29034) );
na02f80 g770450 ( .a(n_10497), .b(n_44464), .o(n_10598) );
no02f80 g743406 ( .a(n_36568), .b(n_36586), .o(n_36709) );
in01f80 FE_RC_2175_0 ( .a(n_26202), .o(FE_RN_775_0) );
in01f80 FE_OCP_RBC1372_n_35275 ( .a(n_35275), .o(FE_OCP_RBN1372_n_35275) );
in01f80 g780451 ( .a(n_881), .o(n_803) );
no02f80 g771988 ( .a(n_44592), .b(n_8809), .o(n_8955) );
in01f80 g778993 ( .a(n_2228), .o(n_2229) );
in01f80 g771487 ( .a(n_9485), .o(n_9523) );
no02f80 g749330 ( .a(n_30627), .b(n_30649), .o(n_30733) );
na02f80 g754480 ( .a(n_26352), .b(FE_OCP_RBN2959_n_26231), .o(n_26831) );
na02f80 g773197 ( .a(n_7650), .b(n_7700), .o(n_7739) );
oa12f80 g762907 ( .a(n_18035), .b(n_18034), .c(n_18033), .o(n_18102) );
no02f80 g742140 ( .a(n_38007), .b(n_37570), .o(n_38121) );
no02f80 FE_RC_1284_0 ( .a(FE_RN_380_0), .b(n_3032), .o(n_47022) );
in01f80 FE_RC_2509_0 ( .a(n_17967), .o(FE_RN_1020_0) );
no02f80 g738112 ( .a(n_42057), .b(n_42056), .o(n_42058) );
na02f80 g780549 ( .a(FE_OCPN852_n_694), .b(n_420), .o(n_1111) );
no02f80 g767324 ( .a(n_13390), .b(n_13368), .o(n_13436) );
in01f80 g779078 ( .a(n_2068), .o(n_2069) );
no02f80 g771093 ( .a(n_9514), .b(FE_OCP_RBN2439_n_8402), .o(n_9672) );
ao12f80 g761281 ( .a(n_18473), .b(n_18832), .c(n_47246), .o(n_18955) );
in01f80 FE_OCP_RBC1056_n_18267 ( .a(n_18267), .o(FE_OCP_RBN1056_n_18267) );
na02f80 g751983 ( .a(n_28782), .b(n_27994), .o(n_28840) );
na02f80 g767475 ( .a(n_13145), .b(FE_OCP_RBN1145_n_13098), .o(n_13231) );
in01f80 FE_OFC795_n_45813 ( .a(FE_OFN793_n_45813), .o(FE_OFN795_n_45813) );
no02f80 g779004 ( .a(n_2172), .b(n_1930), .o(n_2186) );
na02f80 g780578 ( .a(n_663), .b(n_546), .o(n_674) );
no02f80 g739270 ( .a(n_44775), .b(n_40817), .o(n_40881) );
no02f80 g752961 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n_28175) );
no02f80 g778484 ( .a(n_2876), .b(n_2741), .o(n_2935) );
in01f80 newInst_1640 ( .a(newNet_1639), .o(newNet_1640) );
in01f80 g743349 ( .a(n_36693), .o(n_36694) );
na02f80 g761258 ( .a(n_19764), .b(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_19765) );
no02f80 g758655 ( .a(n_21769), .b(n_21793), .o(n_21902) );
in01f80 g762003 ( .a(n_18634), .o(n_19478) );
oa12f80 g769100 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(n_11611), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n_11751) );
na03f80 g760977 ( .a(n_18850), .b(n_19275), .c(n_18914), .o(n_19416) );
in01f80 newInst_2343 ( .a(newNet_2342), .o(newNet_2343) );
oa12f80 g749603 ( .a(n_31581), .b(n_31582), .c(n_31580), .o(n_31671) );
in01f80 newInst_1440 ( .a(newNet_1439), .o(newNet_1440) );
no02f80 g746321 ( .a(n_34916), .b(n_34915), .o(n_34917) );
oa22f80 g752513 ( .a(n_27622), .b(n_24350), .c(n_27607), .d(n_27845), .o(n_27652) );
no02f80 g742069 ( .a(n_37973), .b(n_37637), .o(n_38005) );
in01f80 FE_OCPC1441_n_45060 ( .a(n_45060), .o(FE_OCPN1441_n_45060) );
in01f80 g763219 ( .a(n_17282), .o(n_17444) );
na02f80 g772204 ( .a(n_8812), .b(n_8761), .o(n_8857) );
na02f80 g756300 ( .a(n_24609), .b(n_24033), .o(n_24608) );
na02f80 g771368 ( .a(n_9345), .b(n_9243), .o(n_9346) );
no02f80 g758084 ( .a(n_21973), .b(FE_OCP_RBN1911_n_20545), .o(n_22028) );
ao12f80 g747963 ( .a(n_32646), .b(n_33041), .c(n_32555), .o(n_33172) );
in01f80 FE_OCP_RBC3036_n_47269 ( .a(n_47269), .o(FE_OCP_RBN3036_n_47269) );
ao12f80 g761240 ( .a(n_19035), .b(n_18984), .c(n_18980), .o(n_19142) );
no02f80 g771067 ( .a(n_9636), .b(n_9685), .o(n_9745) );
ao22s80 FE_RC_936_0 ( .a(FE_OCPN1508_n_23414), .b(n_26276), .c(FE_OCP_RBN2940_n_26276), .d(n_23466), .o(n_26424) );
na02f80 g774779 ( .a(n_6327), .b(n_6367), .o(n_6456) );
na02f80 g774333 ( .a(n_6667), .b(n_5471), .o(n_6668) );
no02f80 g739102 ( .a(n_41048), .b(n_40939), .o(n_41047) );
na02f80 g759471 ( .a(n_21110), .b(FE_OCP_RBN1729_n_20903), .o(n_21111) );
na02f80 g762368 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18488), .o(n_18612) );
in01f80 newInst_3651 ( .a(newNet_599), .o(newNet_3651) );
in01f80 newInst_3455 ( .a(newNet_3454), .o(newNet_3455) );
in01f80 newInst_580 ( .a(newNet_579), .o(newNet_580) );
ao22s80 FE_RC_3806_0 ( .a(n_25594), .b(n_25940), .c(n_25593), .d(n_25918), .o(n_26020) );
no02f80 g755113 ( .a(n_25173), .b(FE_OCP_RBN1130_n_24179), .o(n_25353) );
in01f80 FE_RC_3605_0 ( .a(FE_OCP_RBN1342_n_19077), .o(FE_RN_1576_0) );
in01f80 g776362 ( .a(n_4714), .o(n_4715) );
in01f80 newInst_2729 ( .a(newNet_2728), .o(newNet_2729) );
in01f80 g763044 ( .a(n_17587), .o(n_17648) );
na02f80 g766076 ( .a(n_14689), .b(n_14685), .o(n_14686) );
in01f80 newInst_2630 ( .a(newNet_2123), .o(newNet_2630) );
no02f80 g752237 ( .a(n_44723), .b(delay_xor_ln21_unr18_stage7_stallmux_q_7_), .o(n_28058) );
in01f80 FE_RC_3672_0 ( .a(FE_OCPN1533_n_29842), .o(FE_RN_1613_0) );
in01f80 FE_OCP_RBC3079_n_16977 ( .a(n_16977), .o(FE_OCP_RBN3079_n_16977) );
no02f80 FE_RC_1355_0 ( .a(FE_RN_402_0), .b(FE_OCP_RBN2846_n_30678), .o(FE_RN_404_0) );
in01f80 g769265 ( .a(n_11500), .o(n_11501) );
in01f80 g744145 ( .a(n_35945), .o(n_35946) );
in01f80 fopt782877 ( .a(n_39290), .o(n_44312) );
no02f80 g744303 ( .a(n_44180), .b(n_35132), .o(n_36059) );
in01f80 g737781 ( .a(n_42408), .o(n_42409) );
na02f80 g779417 ( .a(n_1467), .b(n_1455), .o(n_1495) );
na02f80 g766874 ( .a(n_14008), .b(n_14042), .o(n_14080) );
na02f80 g774483 ( .a(n_6563), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_5_), .o(n_6569) );
in01f80 g746448 ( .a(n_33307), .o(n_33308) );
oa22f80 g753572 ( .a(n_27322), .b(n_26736), .c(n_27321), .d(n_26737), .o(n_27448) );
in01f80 newInst_1442 ( .a(newNet_1441), .o(newNet_1442) );
in01f80 newInst_575 ( .a(newNet_397), .o(newNet_575) );
no02f80 g777770 ( .a(n_3300), .b(n_3231), .o(n_3350) );
na02f80 g749611 ( .a(n_30483), .b(n_30482), .o(n_30484) );
oa22f80 g741533 ( .a(n_38684), .b(n_38778), .c(n_38683), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38729) );
ao12f80 g749752 ( .a(n_29951), .b(n_29961), .c(n_29857), .o(n_30055) );
oa22f80 FE_RC_1670_0 ( .a(delay_sub_ln23_0_unr29_stage10_stallmux_q), .b(n_42128), .c(n_42196), .d(n_42129), .o(n_42156) );
oa22f80 g764131 ( .a(n_16576), .b(n_16594), .c(n_16552), .d(n_16595), .o(n_16699) );
in01f80 g752246 ( .a(n_28002), .o(n_28003) );
oa12f80 g757171 ( .a(n_23185), .b(n_44996), .c(n_23118), .o(n_23616) );
in01f80 newInst_927 ( .a(newNet_926), .o(newNet_927) );
in01f80 g774665 ( .a(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6872) );
no02f80 g751387 ( .a(n_28651), .b(n_28577), .o(n_28681) );
na02f80 g743261 ( .a(n_36828), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .o(n_36931) );
in01f80 g745576 ( .a(n_34320), .o(n_34340) );
in01f80 FE_RC_2321_0 ( .a(FE_RN_883_0), .o(n_45740) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_1_ ( .ck(newNet_1621), .d(n_26997), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_1_) );
na02f80 g770428 ( .a(n_10607), .b(FE_OCP_RBN2568_n_8904), .o(n_10634) );
na02f80 g750174 ( .a(n_29861), .b(FE_OCP_DRV_N1572_n_29860), .o(n_29955) );
ao22s80 g755941 ( .a(n_25160), .b(n_24258), .c(n_25188), .d(n_25002), .o(n_25525) );
in01f80 g756132 ( .a(n_25032), .o(n_25139) );
in01f80 newInst_1232 ( .a(newNet_1231), .o(newNet_1232) );
in01f80 newInst_45 ( .a(newNet_44), .o(newNet_45) );
in01f80 FE_RC_2751_0 ( .a(n_43359), .o(FE_RN_1169_0) );
in01f80 newInst_646 ( .a(newNet_645), .o(newNet_646) );
in01f80 newInst_3487 ( .a(newNet_3486), .o(newNet_3487) );
no02f80 g741291 ( .a(n_44955), .b(n_38907), .o(n_38997) );
na02f80 g778376 ( .a(n_2508), .b(n_2477), .o(n_2478) );
in01f80 FE_RC_1070_0 ( .a(n_11975), .o(FE_RN_316_0) );
na02f80 g750706 ( .a(n_29341), .b(n_29389), .o(n_29437) );
in01f80 g736460 ( .a(n_43764), .o(n_43765) );
in01f80 FE_OCPC3746_n_29439 ( .a(n_29439), .o(FE_OCPN3746_n_29439) );
na02f80 g738883 ( .a(n_41200), .b(n_41049), .o(n_41256) );
na02f80 g743953 ( .a(n_36304), .b(n_35700), .o(n_36320) );
na02f80 g757694 ( .a(n_45203), .b(n_44061), .o(n_22634) );
no02f80 g738977 ( .a(n_41149), .b(n_40914), .o(n_41166) );
no02f80 g778773 ( .a(n_2327), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_), .o(n_2367) );
no02f80 g762227 ( .a(n_18096), .b(n_18024), .o(n_18097) );
na02f80 g769684 ( .a(FE_OCP_RBN3706_n_11146), .b(n_44498), .o(n_11203) );
na02f80 g750180 ( .a(n_29754), .b(n_28657), .o(n_29815) );
na02f80 g737052 ( .a(n_43230), .b(n_43170), .o(n_43484) );
na02f80 g745944 ( .a(n_33969), .b(n_33968), .o(n_34041) );
no02f80 g755677 ( .a(n_24434), .b(n_24412), .o(n_24534) );
in01f80 g775367 ( .a(n_5798), .o(n_5805) );
in01f80 FE_OCP_RBC3308_n_44722 ( .a(FE_OCP_RBN3310_n_44722), .o(FE_OCP_RBN3308_n_44722) );
oa12f80 g754534 ( .a(n_26239), .b(n_26238), .c(n_26237), .o(n_26907) );
no02f80 g736826 ( .a(n_43204), .b(n_43311), .o(n_43344) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_1_ ( .ck(newNet_499), .d(n_22480), .o(n_45204) );
na02f80 g739566 ( .a(n_40609), .b(n_40617), .o(n_40631) );
in01f80 g750535 ( .a(n_29500), .o(n_29546) );
in01f80 g739802 ( .a(n_40423), .o(n_40424) );
na02f80 FE_RC_1560_0 ( .a(FE_RN_443_0), .b(n_2735), .o(n_2821) );
ao12f80 g774217 ( .a(n_6633), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_8_), .o(n_6689) );
na02f80 g776507 ( .a(n_4483), .b(n_4594), .o(n_4780) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_26_ ( .ck(newNet_316), .d(n_1286), .o(delay_xor_ln22_unr3_stage2_stallmux_q_26_) );
oa22f80 g738123 ( .a(n_42016), .b(n_41856), .c(n_42029), .d(n_41857), .o(n_42570) );
na02f80 g749159 ( .a(n_30808), .b(n_30828), .o(n_30908) );
oa22f80 g779168 ( .a(n_1864), .b(n_1689), .c(FE_OCP_RBN2177_n_1864), .d(n_1688), .o(n_1955) );
in01f80 newInst_603 ( .a(newNet_265), .o(newNet_603) );
in01f80 g766889 ( .a(n_14300), .o(n_14301) );
in01f80 FE_RC_4139_0 ( .a(n_45224), .o(FE_RN_1798_0) );
in01f80 g748053 ( .a(n_31708), .o(n_31748) );
no02f80 g741401 ( .a(n_38844), .b(n_38843), .o(n_38845) );
in01f80 FE_RC_2113_0 ( .a(FE_RN_732_0), .o(n_21239) );
in01f80 g773088 ( .a(n_8081), .o(n_8047) );
oa12f80 g754451 ( .a(n_26939), .b(n_26938), .c(n_26937), .o(n_26998) );
ao12f80 g738343 ( .a(n_41735), .b(n_41639), .c(FE_OCP_RBN2316_n_41420), .o(n_41755) );
na02f80 g762393 ( .a(n_45118), .b(n_17785), .o(n_18622) );
in01f80 g751175 ( .a(n_29995), .o(n_29976) );
no02f80 g758617 ( .a(FE_OCPN3178_n_21901), .b(n_21902), .o(n_21921) );
in01f80 g750604 ( .a(n_29383), .o(n_29384) );
ao12f80 g756257 ( .a(n_24674), .b(n_24673), .c(n_24672), .o(n_25130) );
in01f80 FE_RC_3681_0 ( .a(FE_OCPN1017_n_23307), .o(FE_RN_1616_0) );
na02f80 g778107 ( .a(n_2826), .b(n_2938), .o(n_2939) );
no02f80 g736993 ( .a(n_43082), .b(n_43134), .o(n_43266) );
in01f80 newInst_814 ( .a(newNet_813), .o(newNet_814) );
na02f80 g744091 ( .a(n_44256), .b(n_34629), .o(n_35643) );
no02f80 g765530 ( .a(n_15599), .b(n_15718), .o(n_15873) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_21_ ( .ck(newNet_1612), .d(n_27323), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_21_) );
in01f80 newInst_796 ( .a(newNet_235), .o(newNet_796) );
in01f80 g759331 ( .a(n_21149), .o(n_21150) );
na02f80 g773636 ( .a(n_7389), .b(n_7048), .o(n_7390) );
no02f80 g756928 ( .a(n_23900), .b(n_23831), .o(n_24379) );
ao12f80 g751811 ( .a(n_29148), .b(n_29172), .c(n_28919), .o(n_29801) );
no02f80 g741119 ( .a(n_39149), .b(FE_OCP_RBN2603_n_39126), .o(n_39205) );
ao12f80 g738445 ( .a(n_41707), .b(n_41660), .c(n_41310), .o(n_41881) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_10_ ( .ck(newNet_1265), .d(n_5211), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_) );
oa22f80 g784549 ( .a(FE_OFN801_n_46285), .b(n_11212), .c(FE_OCP_RBN3044_n_46337), .d(n_11184), .o(n_46370) );
in01f80 FE_RC_2043_0 ( .a(n_25624), .o(FE_RN_685_0) );
na02f80 g744036 ( .a(FE_OCPN3751_n_44222), .b(n_35703), .o(n_36267) );
in01f80 fopt783405 ( .a(n_45010), .o(n_45008) );
ao12f80 g748948 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_8_), .o(n_32501) );
ao22s80 g780345 ( .a(n_807), .b(n_1203), .c(n_851), .d(FE_OFN795_n_45813), .o(n_918) );
oa22f80 FE_RC_1198_0 ( .a(n_15567), .b(n_15802), .c(n_15568), .d(n_15803), .o(n_16003) );
no02f80 g752128 ( .a(FE_OCPN877_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_9_), .o(n_28014) );
oa22f80 FE_RC_3215_0 ( .a(n_990), .b(n_44636), .c(n_1014), .d(n_1282), .o(n_1285) );
na02f80 g763237 ( .a(n_17243), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_), .o(n_17398) );
oa12f80 g765801 ( .a(n_14646), .b(n_14891), .c(n_14647), .o(n_14912) );
in01f80 FE_OCP_RBC2887_n_10570 ( .a(n_10570), .o(FE_OCP_RBN2887_n_10570) );
na02f80 g764575 ( .a(n_15997), .b(n_16048), .o(n_16113) );
ao12f80 g742722 ( .a(n_37321), .b(n_37320), .c(n_37319), .o(n_37398) );
in01f80 FE_OCP_RBC2134_n_45508 ( .a(n_45508), .o(FE_OCP_RBN2134_n_45508) );
in01f80 g758598 ( .a(n_21965), .o(n_21966) );
ao12f80 g767385 ( .a(n_12695), .b(n_13235), .c(n_12733), .o(n_13336) );
in01f80 FE_RC_1638_0 ( .a(n_23066), .o(FE_RN_456_0) );
na02f80 g769753 ( .a(n_11010), .b(n_11054), .o(n_11146) );
oa12f80 g746021 ( .a(n_34742), .b(n_35191), .c(n_34695), .o(n_35241) );
no02f80 g761121 ( .a(n_19151), .b(n_19175), .o(n_19264) );
na02f80 g741632 ( .a(n_38591), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38624) );
in01f80 g750700 ( .a(n_29413), .o(n_29414) );
in01f80 g763828 ( .a(n_17258), .o(n_17259) );
in01f80 g778241 ( .a(n_2699), .o(n_2645) );
na02f80 g768019 ( .a(n_12616), .b(n_12431), .o(n_12651) );
in01f80 g767312 ( .a(n_13410), .o(n_13411) );
in01f80 FE_RC_2921_0 ( .a(FE_RN_1271_0), .o(n_27620) );
in01f80 newInst_2420 ( .a(newNet_2419), .o(newNet_2420) );
na02f80 g744609 ( .a(n_35349), .b(n_35348), .o(n_35350) );
na03f80 g742461 ( .a(n_37561), .b(n_37563), .c(n_37056), .o(n_37583) );
no02f80 g739013 ( .a(n_41098), .b(n_40830), .o(n_41149) );
na02f80 g749833 ( .a(FE_OCP_RBN3019_n_31117), .b(n_31038), .o(n_31254) );
oa12f80 g757911 ( .a(n_22725), .b(n_22952), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_29_), .o(n_23119) );
na02f80 g737213 ( .a(n_42920), .b(n_42935), .o(n_43298) );
in01f80 g743075 ( .a(n_37086), .o(n_37087) );
ao22s80 FE_RC_4086_0 ( .a(FE_RN_1782_0), .b(FE_RN_1781_0), .c(FE_RN_1786_0), .d(n_17292), .o(n_17417) );
in01f80 g752405 ( .a(n_27804), .o(n_27774) );
ao22s80 FE_RC_251_0 ( .a(n_14441), .b(FE_OCP_RBN3535_n_13765), .c(FE_OCP_RBN3532_n_13765), .d(n_16215), .o(n_14571) );
na02f80 g738028 ( .a(n_42163), .b(n_42162), .o(n_42164) );
na02f80 g749664 ( .a(n_30150), .b(n_29925), .o(n_30248) );
oa12f80 g744586 ( .a(n_36021), .b(n_36598), .c(n_35880), .o(n_36664) );
in01f80 g738401 ( .a(n_41856), .o(n_41857) );
oa22f80 g748203 ( .a(n_31713), .b(n_31700), .c(n_31714), .d(n_31701), .o(n_31806) );
na02f80 g777801 ( .a(n_3285), .b(n_3257), .o(n_3335) );
in01f80 FE_OCP_RBC2675_n_14991 ( .a(FE_OCP_RBN2674_n_14991), .o(FE_OCP_RBN2675_n_14991) );
in01f80 newInst_2452 ( .a(newNet_2451), .o(newNet_2452) );
in01f80 g774835 ( .a(n_6316), .o(n_6317) );
no02f80 g744575 ( .a(n_35351), .b(n_35318), .o(n_35402) );
na02f80 g758978 ( .a(n_21392), .b(n_21322), .o(n_21545) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_4_ ( .ck(newNet_1902), .d(n_36800), .o(delay_sub_ln22_unr24_stage9_stallmux_q_4_) );
no02f80 g776037 ( .a(n_4945), .b(n_4372), .o(n_5144) );
no02f80 g754296 ( .a(n_25828), .b(n_25482), .o(n_25902) );
no03m80 g743355 ( .a(n_37751), .b(n_37826), .c(n_37784), .o(n_37854) );
no02f80 g740600 ( .a(FE_OCP_RBN2894_n_39575), .b(n_45841), .o(n_39606) );
in01f80 g765524 ( .a(n_15967), .o(n_15919) );
ao22s80 g771908 ( .a(n_8700), .b(n_7632), .c(n_45503), .d(n_7631), .o(n_8767) );
in01f80 g767214 ( .a(FE_OCPN1006_n_13962), .o(n_14215) );
in01f80 g764194 ( .a(n_16530), .o(n_16531) );
in01f80 g777098 ( .a(n_3809), .o(n_3810) );
no02f80 g759108 ( .a(n_21387), .b(n_21175), .o(n_21464) );
no02f80 g759671 ( .a(n_20478), .b(n_45101), .o(n_20547) );
na02f80 g745448 ( .a(n_34298), .b(n_34273), .o(n_34274) );
in01f80 g775027 ( .a(n_6118), .o(n_6125) );
in01f80 g746047 ( .a(n_34224), .o(n_34206) );
no02f80 g741625 ( .a(n_38586), .b(n_38778), .o(n_38602) );
no02f80 g744940 ( .a(n_34995), .b(n_34704), .o(n_35048) );
ao12f80 g750315 ( .a(n_30101), .b(n_30688), .c(n_30126), .o(n_30838) );
in01f80 newInst_31 ( .a(newNet_30), .o(newNet_31) );
in01f80 g760024 ( .a(n_21374), .o(n_21406) );
na02f80 g738697 ( .a(n_41491), .b(n_41490), .o(n_41536) );
no02f80 g745067 ( .a(n_34727), .b(n_47254), .o(n_34771) );
na02f80 g764429 ( .a(FE_OCP_RBN2905_n_16197), .b(FE_OCPN3775_n_14730), .o(n_16225) );
in01f80 g757165 ( .a(n_23700), .o(n_23743) );
no02f80 FE_RC_4236_0 ( .a(FE_RN_1860_0), .b(n_26087), .o(FE_RN_696_0) );
no02f80 g742988 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_12_), .o(n_37016) );
in01f80 FE_OCP_RBC3577_n_4528 ( .a(FE_OCP_RBN3575_n_4528), .o(FE_OCP_RBN3577_n_4528) );
ao22s80 FE_RC_3341_0 ( .a(n_30145), .b(n_45629), .c(n_45630), .d(n_30146), .o(n_30428) );
in01f80 FE_OCP_RBC1057_n_18267 ( .a(FE_OCP_RBN1056_n_18267), .o(FE_OCP_RBN1057_n_18267) );
oa22f80 FE_RC_1366_0 ( .a(n_10494), .b(n_10880), .c(n_10495), .d(n_10881), .o(n_11004) );
na02f80 g753846 ( .a(n_27067), .b(n_26610), .o(n_27097) );
na03f80 FE_RC_1301_0 ( .a(n_4070), .b(n_3926), .c(n_4098), .o(n_4173) );
in01f80 g744567 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_20_), .o(n_36744) );
no02f80 g765476 ( .a(n_15041), .b(FE_OCP_RBN3655_n_15097), .o(n_15186) );
in01f80 newInst_1383 ( .a(newNet_1382), .o(newNet_1383) );
in01f80 fopt783183 ( .a(FE_OCP_RBN3308_n_44722), .o(n_44723) );
ao22s80 g780193 ( .a(n_1067), .b(FE_OFN761_n_45813), .c(n_1089), .d(n_1203), .o(n_1143) );
oa22f80 g739705 ( .a(n_40473), .b(n_40283), .c(n_40474), .d(n_40284), .o(n_40507) );
in01f80 g748090 ( .a(n_31668), .o(n_31669) );
in01f80 FE_RC_2261_0 ( .a(n_24605), .o(FE_RN_837_0) );
na02f80 FE_RC_4084_0 ( .a(FE_OCP_RBN2851_n_46982), .b(FE_RN_1783_0), .o(FE_RN_1785_0) );
na02f80 FE_RC_3799_0 ( .a(FE_RN_1660_0), .b(n_20024), .o(FE_RN_1257_0) );
oa12f80 g759678 ( .a(n_21566), .b(n_21449), .c(n_21374), .o(n_21629) );
ao12f80 g774206 ( .a(n_6868), .b(n_6806), .c(delay_xor_ln21_unr6_stage3_stallmux_q_12_), .o(n_6928) );
no02f80 FE_RC_2690_0 ( .a(FE_RN_1126_0), .b(FE_OCP_RBN2564_FE_RN_1125_0), .o(n_9351) );
in01f80 g763321 ( .a(n_17384), .o(n_17385) );
no02f80 g768330 ( .a(n_12486), .b(n_12485), .o(n_12487) );
ao12f80 g776269 ( .a(n_4482), .b(n_4594), .c(n_4827), .o(n_4951) );
in01f80 FE_OCP_RBC2683_n_35213 ( .a(n_35213), .o(FE_OCP_RBN2683_n_35213) );
no02f80 g738262 ( .a(n_41873), .b(n_41872), .o(n_41874) );
in01f80 g736469 ( .a(n_43754), .o(n_43755) );
na02f80 g756767 ( .a(n_23395), .b(n_23427), .o(n_23587) );
ao12f80 g756891 ( .a(n_23311), .b(n_23310), .c(n_23309), .o(n_24613) );
na02f80 g778336 ( .a(n_2554), .b(FE_OCP_RBN2267_n_2430), .o(n_2555) );
ao12f80 g779238 ( .a(n_1590), .b(n_1756), .c(n_1463), .o(n_1859) );
na02f80 g758174 ( .a(n_44277), .b(n_22076), .o(n_22153) );
no02f80 g775658 ( .a(FE_OCP_RBN3688_n_5130), .b(n_4606), .o(n_5190) );
no02f80 g761768 ( .a(n_19232), .b(n_19231), .o(n_19233) );
na02f80 FE_RC_2670_0 ( .a(n_4953), .b(n_3637), .o(FE_RN_1117_0) );
oa22f80 g749344 ( .a(n_31979), .b(n_31369), .c(n_31980), .d(n_31370), .o(n_32064) );
in01f80 newInst_2173 ( .a(newNet_2172), .o(newNet_2173) );
in01f80 g749507 ( .a(n_31599), .o(n_30637) );
in01f80 g776887 ( .a(n_4113), .o(n_4114) );
in01f80 newInst_2782 ( .a(newNet_2781), .o(newNet_2782) );
in01f80 g780336 ( .a(n_897), .o(n_966) );
na02f80 g760672 ( .a(n_19646), .b(n_19669), .o(n_19783) );
oa12f80 g778558 ( .a(n_2497), .b(n_2514), .c(n_2496), .o(n_2628) );
na02f80 g745733 ( .a(n_34303), .b(n_34004), .o(n_34337) );
in01f80 g769648 ( .a(n_11366), .o(n_11367) );
in01f80 g737364 ( .a(n_42829), .o(n_43147) );
in01f80 fopt782834 ( .a(n_33693), .o(n_44259) );
no02f80 g767236 ( .a(n_13701), .b(n_13285), .o(n_13791) );
in01f80 g778447 ( .a(n_2453), .o(n_2502) );
in01f80 newInst_914 ( .a(newNet_609), .o(newNet_914) );
na02f80 g772571 ( .a(n_8296), .b(FE_OCPN890_n_7802), .o(n_8326) );
oa12f80 g768698 ( .a(n_11935), .b(n_44451), .c(n_12003), .o(n_12202) );
in01f80 FE_OCPC1785_n_30134 ( .a(FE_OCP_RBN2572_n_29922), .o(FE_OCPN1785_n_30134) );
in01f80 g757738 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_17_), .o(n_23562) );
no02f80 g781346 ( .a(n_7), .b(beta_27), .o(n_100) );
no02f80 g756443 ( .a(n_23606), .b(n_23660), .o(n_23775) );
na02f80 FE_RC_3667_0 ( .a(n_24848), .b(n_26440), .o(FE_RN_1610_0) );
in01f80 g760103 ( .a(n_20195), .o(n_20215) );
no02f80 g747230 ( .a(n_32627), .b(n_32626), .o(n_32702) );
oa22f80 FE_RC_3308_0 ( .a(n_30274), .b(n_30501), .c(n_30273), .d(n_30512), .o(n_30608) );
ao22s80 g751345 ( .a(n_28611), .b(n_28418), .c(n_28551), .d(n_28417), .o(n_28654) );
in01f80 newInst_930 ( .a(newNet_929), .o(newNet_930) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_8_ ( .ck(newNet_3576), .d(n_15979), .o(delay_add_ln22_unr11_stage5_stallmux_q_8_) );
in01f80 FE_RC_4079_0 ( .a(FE_OCP_RBN2812_n_15433), .o(FE_RN_1779_0) );
in01f80 g762759 ( .a(n_17811), .o(n_17781) );
oa22f80 g751089 ( .a(n_30303), .b(n_30083), .c(n_30156), .d(n_29691), .o(n_30720) );
no02f80 g763911 ( .a(n_17015), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_11_), .o(n_17425) );
in01f80 g740568 ( .a(n_39697), .o(n_39706) );
na02f80 g767692 ( .a(n_12824), .b(n_12900), .o(n_12935) );
in01f80 g776278 ( .a(n_4654), .o(n_4655) );
no02f80 g776658 ( .a(n_3916), .b(n_3834), .o(n_4101) );
oa12f80 g776607 ( .a(n_4500), .b(n_4499), .c(n_4498), .o(n_4600) );
na02f80 g751272 ( .a(n_29747), .b(n_29746), .o(n_29748) );
na02f80 g776046 ( .a(n_4989), .b(FE_OCP_RBN2609_n_3807), .o(n_5134) );
in01f80 g772608 ( .a(n_8261), .o(n_8294) );
na02f80 g749810 ( .a(n_31285), .b(n_31508), .o(n_31621) );
in01f80 g755568 ( .a(n_24684), .o(n_24717) );
na02f80 g758862 ( .a(n_21474), .b(n_21544), .o(n_21579) );
no02f80 g767038 ( .a(FE_OCP_RBN2458_n_13765), .b(n_13875), .o(n_13900) );
in01f80 g766927 ( .a(n_14076), .o(n_14077) );
na02f80 g743423 ( .a(n_36632), .b(n_36750), .o(n_36633) );
in01f80 g769160 ( .a(delay_xor_ln21_unr9_stage4_stallmux_q_1_), .o(n_11561) );
no02f80 g779573 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_11_), .o(n_1695) );
in01f80 g748982 ( .a(n_31151), .o(n_31152) );
na02f80 g755129 ( .a(n_25374), .b(n_24469), .o(n_25501) );
oa12f80 g745565 ( .a(n_35480), .b(n_35479), .c(n_35478), .o(n_35926) );
in01f80 newInst_2950 ( .a(newNet_2949), .o(newNet_2950) );
na02f80 g780133 ( .a(n_1085), .b(n_1084), .o(n_1086) );
in01f80 FE_OCP_RBC3493_n_19390 ( .a(n_19390), .o(FE_OCP_RBN3493_n_19390) );
na02f80 FE_RC_2559_0 ( .a(n_6698), .b(n_6896), .o(FE_RN_1049_0) );
in01f80 g780905 ( .a(n_432), .o(n_448) );
in01f80 g745751 ( .a(n_34281), .o(n_34282) );
in01f80 g765690 ( .a(n_16338), .o(n_17336) );
in01f80 g766666 ( .a(n_13815), .o(n_13816) );
na02f80 g777259 ( .a(n_3492), .b(n_2764), .o(n_3493) );
no02f80 g768583 ( .a(n_12234), .b(n_11795), .o(n_12268) );
in01f80 FE_OCP_RBC3614_n_20249 ( .a(FE_OCP_RBN2670_n_20249), .o(FE_OCP_RBN3614_n_20249) );
in01f80 newInst_673 ( .a(newNet_672), .o(newNet_673) );
oa12f80 g768946 ( .a(n_11637), .b(n_11775), .c(n_11636), .o(n_11787) );
no02f80 g780754 ( .a(n_576), .b(n_568), .o(n_569) );
in01f80 newInst_2803 ( .a(newNet_298), .o(newNet_2803) );
in01f80 newInst_2329 ( .a(newNet_831), .o(newNet_2329) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_14_ ( .ck(newNet_3074), .d(n_1164), .o(delay_add_ln22_unr2_stage2_stallmux_q_14_) );
no02f80 g770139 ( .a(n_10711), .b(n_10391), .o(n_10738) );
in01f80 newInst_316 ( .a(newNet_315), .o(newNet_316) );
na02f80 FE_RC_2123_0 ( .a(FE_RN_738_0), .b(n_21090), .o(FE_RN_739_0) );
no02f80 g751851 ( .a(n_29073), .b(n_29044), .o(n_29102) );
oa12f80 g772988 ( .a(n_7773), .b(n_45846), .c(n_45871), .o(n_8091) );
in01f80 g766173 ( .a(n_14868), .o(n_14894) );
na02f80 g766330 ( .a(n_14400), .b(n_14319), .o(n_14436) );
no02f80 FE_RC_2315_0 ( .a(FE_RN_879_0), .b(n_35935), .o(FE_RN_880_0) );
in01f80 newInst_1004 ( .a(newNet_642), .o(newNet_1004) );
no02f80 g738058 ( .a(n_42092), .b(n_41906), .o(n_42120) );
ao12f80 g761362 ( .a(n_19954), .b(n_19980), .c(n_19900), .o(n_20898) );
no02f80 g768799 ( .a(n_12034), .b(n_12033), .o(n_12035) );
na02f80 g771557 ( .a(n_9365), .b(n_9334), .o(n_9526) );
in01f80 g749208 ( .a(n_30769), .o(n_30770) );
no02f80 g741808 ( .a(n_38342), .b(n_38142), .o(n_38425) );
in01f80 FE_RC_2033_0 ( .a(FE_OFN738_n_22641), .o(FE_RN_678_0) );
in01f80 FE_OFC779_n_17093 ( .a(FE_OFN777_n_17093), .o(FE_OFN779_n_17093) );
no02f80 g750542 ( .a(n_29407), .b(n_47251), .o(n_29429) );
na02f80 g760973 ( .a(n_19318), .b(n_19152), .o(n_19356) );
in01f80 g780499 ( .a(n_930), .o(n_931) );
in01f80 g757759 ( .a(n_46965), .o(n_22594) );
oa22f80 g773631 ( .a(n_7306), .b(n_7199), .c(n_7277), .d(n_7198), .o(n_7372) );
in01f80 newInst_3190 ( .a(newNet_1311), .o(newNet_3190) );
ao12f80 g742931 ( .a(n_37004), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n_37468) );
in01f80 newInst_165 ( .a(newNet_164), .o(newNet_165) );
in01f80 g740944 ( .a(n_39283), .o(n_39284) );
na02f80 g745243 ( .a(n_35939), .b(n_35996), .o(n_36025) );
na02f80 g751915 ( .a(n_28919), .b(n_29076), .o(n_29309) );
in01f80 newInst_2464 ( .a(newNet_2463), .o(newNet_2464) );
in01f80 newInst_1538 ( .a(newNet_1537), .o(newNet_1538) );
na02f80 g746993 ( .a(n_34104), .b(n_34103), .o(n_34105) );
in01f80 g748058 ( .a(n_31935), .o(n_31954) );
in01f80 g758046 ( .a(n_23053), .o(n_23054) );
in01f80 FE_OCP_RBC2496_n_8641 ( .a(FE_OCP_RBN2495_n_8641), .o(FE_OCP_RBN2496_n_8641) );
in01f80 newInst_3062 ( .a(newNet_3061), .o(newNet_3062) );
no02f80 g743085 ( .a(n_36923), .b(n_36922), .o(n_36924) );
in01f80 g767521 ( .a(n_13142), .o(n_13143) );
in01f80 FE_OCP_RBC2355_n_13858 ( .a(FE_OCP_RBN2353_n_13858), .o(FE_OCP_RBN2355_n_13858) );
in01f80 g738334 ( .a(n_41860), .o(n_41861) );
no02f80 g776256 ( .a(n_4846), .b(n_4369), .o(n_4866) );
in01f80 g772284 ( .a(n_8666), .o(n_8667) );
ao12f80 g751868 ( .a(n_28057), .b(n_28123), .c(n_28184), .o(n_28209) );
na02f80 g741278 ( .a(n_44944), .b(n_46951), .o(n_38988) );
no02f80 g767029 ( .a(n_14758), .b(n_14168), .o(n_14208) );
in01f80 newInst_2591 ( .a(newNet_2590), .o(newNet_2591) );
oa12f80 g748115 ( .a(n_31652), .b(n_31606), .c(FE_OCP_RBN3714_n_31466), .o(n_31744) );
in01f80 g767908 ( .a(n_12655), .o(n_12690) );
in01f80 FE_OCP_RBC3122_n_32239 ( .a(n_32239), .o(FE_OCP_RBN3122_n_32239) );
no02f80 g752938 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .o(n_27990) );
in01f80 newInst_2402 ( .a(newNet_1900), .o(newNet_2402) );
ao12f80 g755255 ( .a(n_24942), .b(n_24941), .c(n_24974), .o(n_26656) );
na02f80 g773982 ( .a(n_6919), .b(delay_add_ln22_unr5_stage3_stallmux_q_5_), .o(n_7011) );
oa22f80 g743764 ( .a(n_36047), .b(n_36260), .c(n_36074), .d(n_36261), .o(n_36340) );
oa22f80 g742584 ( .a(n_37499), .b(n_37504), .c(n_37520), .d(n_36768), .o(n_37636) );
in01f80 g772625 ( .a(n_8437), .o(n_8395) );
oa22f80 g764347 ( .a(n_16317), .b(n_14598), .c(n_16423), .d(n_14577), .o(n_16454) );
no02f80 g747436 ( .a(n_33815), .b(n_33763), .o(n_33816) );
na02f80 g761193 ( .a(n_19932), .b(n_19959), .o(n_19960) );
in01f80 g764387 ( .a(n_16675), .o(n_16676) );
na02f80 g765257 ( .a(n_15486), .b(n_15452), .o(n_15601) );
na02f80 g773822 ( .a(n_7090), .b(n_5777), .o(n_7146) );
in01f80 g744206 ( .a(n_36256), .o(n_36257) );
no03m80 FE_RC_1633_0 ( .a(n_17197), .b(FE_OCP_RBN1136_n_17040), .c(n_17245), .o(n_17561) );
oa12f80 g752436 ( .a(n_27848), .b(n_28378), .c(n_27903), .o(n_28397) );
oa22f80 FE_RC_1572_0 ( .a(FE_OCP_RBN3467_n_7886), .b(FE_OCP_RBN2467_n_8767), .c(FE_OCPN1011_n_7802), .d(n_8767), .o(n_8870) );
na02f80 g755434 ( .a(n_24751), .b(n_22484), .o(n_24806) );
na02f80 g773010 ( .a(n_7860), .b(n_7809), .o(n_7927) );
ao12f80 g747191 ( .a(n_32718), .b(n_32668), .c(n_32653), .o(n_32774) );
na02f80 g741749 ( .a(n_38474), .b(n_38159), .o(n_38476) );
in01f80 newInst_1813 ( .a(newNet_1812), .o(newNet_1813) );
in01f80 g772898 ( .a(n_7959), .o(n_8001) );
in01f80 newInst_2491 ( .a(newNet_2002), .o(newNet_2491) );
ao12f80 g738904 ( .a(n_41281), .b(n_41280), .c(n_41279), .o(n_41698) );
in01f80 g739943 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_4_), .o(n_40478) );
in01f80 g737502 ( .a(n_43037), .o(n_42714) );
oa22f80 FE_RC_3769_0 ( .a(FE_RN_1538_0), .b(FE_RN_1539_0), .c(FE_RN_1540_0), .d(n_32638), .o(n_32653) );
oa12f80 g750294 ( .a(n_30167), .b(n_30783), .c(n_30094), .o(n_30898) );
ao12f80 g773883 ( .a(n_6683), .b(n_7094), .c(n_6626), .o(n_7111) );
na02f80 g761818 ( .a(n_18641), .b(n_18431), .o(n_18821) );
na02f80 g772783 ( .a(n_8095), .b(n_8094), .o(n_8127) );
ao12f80 g753739 ( .a(n_26663), .b(n_26478), .c(n_26405), .o(n_26537) );
ao22s80 FE_RC_719_0 ( .a(n_37719), .b(n_37775), .c(n_37734), .d(n_37776), .o(n_37848) );
in01f80 newInst_2294 ( .a(newNet_1554), .o(newNet_2294) );
na02f80 g774823 ( .a(n_45475), .b(n_5469), .o(n_6414) );
in01f80 FE_RC_3666_0 ( .a(FE_RN_1610_0), .o(n_26586) );
na02f80 g768772 ( .a(n_11967), .b(n_11957), .o(n_12098) );
no02f80 FE_RC_3535_0 ( .a(n_17197), .b(FE_RN_1529_0), .o(n_17239) );
oa12f80 g752259 ( .a(n_28499), .b(FE_OCP_RBN2179_FE_RN_526_0), .c(n_28498), .o(n_28669) );
in01f80 FE_OCP_RBC2969_n_26398 ( .a(n_26398), .o(FE_OCP_RBN2969_n_26398) );
no02f80 g742446 ( .a(n_37629), .b(n_37300), .o(n_37694) );
na02f80 g751567 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_30_), .o(n_28741) );
na02f80 g751773 ( .a(n_29008), .b(n_28898), .o(n_29010) );
no02f80 g770045 ( .a(n_10766), .b(n_10469), .o(n_10800) );
na02f80 g738087 ( .a(n_42093), .b(n_42710), .o(n_42094) );
ao12f80 g758153 ( .a(n_22842), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_21_), .o(n_23150) );
in01f80 g755415 ( .a(n_24868), .o(n_24869) );
na02f80 g743651 ( .a(n_36351), .b(n_35782), .o(n_36412) );
no02f80 g758256 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_6_), .o(n_22647) );
in01f80 FE_OCP_RBC2775_n_10100 ( .a(FE_OCP_RBN3653_n_10100), .o(FE_OCP_RBN2775_n_10100) );
in01f80 g745950 ( .a(n_34083), .o(n_34084) );
no02f80 g764798 ( .a(n_15620), .b(n_15653), .o(n_15732) );
in01f80 g753145 ( .a(n_27047), .o(n_27013) );
in01f80 g774585 ( .a(n_6517), .o(n_6563) );
na02f80 g748750 ( .a(n_32503), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_0_), .o(n_32504) );
no02f80 FE_RC_3555_0 ( .a(n_12790), .b(n_13098), .o(FE_RN_1543_0) );
in01f80 FE_RC_709_0 ( .a(n_23047), .o(FE_RN_225_0) );
in01f80 newInst_81 ( .a(newNet_68), .o(newNet_81) );
na02f80 g784772 ( .a(FE_OCP_RBN3614_n_20249), .b(n_19131), .o(n_47258) );
in01f80 FE_OCP_RBC1178_n_18981 ( .a(FE_OCP_RBN1176_n_18981), .o(FE_OCP_RBN1178_n_18981) );
na02f80 g755374 ( .a(n_24766), .b(n_46963), .o(n_24920) );
na02f80 g768116 ( .a(n_12605), .b(delay_add_ln22_unr8_stage4_stallmux_q_18_), .o(n_12633) );
in01f80 g782632 ( .a(n_27885), .o(n_44025) );
in01f80 g775140 ( .a(n_6140), .o(n_6141) );
in01f80 g759687 ( .a(n_21867), .o(n_21868) );
na02f80 g763144 ( .a(n_17395), .b(n_17442), .o(n_17443) );
na02f80 g784400 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .o(n_46212) );
na02f80 g742115 ( .a(n_38049), .b(n_47252), .o(n_38160) );
in01f80 FE_OCP_RBC3447_n_37945 ( .a(FE_OCP_RBN3444_n_37945), .o(FE_OCP_RBN3447_n_37945) );
in01f80 g765283 ( .a(n_15828), .o(n_15929) );
in01f80 FE_OCP_RBC2543_n_9082 ( .a(n_9082), .o(FE_OCP_RBN2543_n_9082) );
in01f80 g752500 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n_27654) );
na02f80 g777939 ( .a(n_47021), .b(n_3080), .o(n_3175) );
na02f80 g744083 ( .a(n_35537), .b(n_35522), .o(n_35523) );
na02f80 g773633 ( .a(n_7288), .b(delay_add_ln22_unr5_stage3_stallmux_q_18_), .o(n_7360) );
in01f80 FE_OCP_RBC2767_n_4376 ( .a(n_4376), .o(FE_OCP_RBN2767_n_4376) );
no02f80 g762282 ( .a(n_18835), .b(n_18569), .o(n_19572) );
in01f80 g753885 ( .a(n_26327), .o(n_26328) );
in01f80 g780544 ( .a(n_831), .o(n_1002) );
in01f80 newInst_3094 ( .a(newNet_3093), .o(newNet_3094) );
na02f80 g778534 ( .a(n_2814), .b(n_2954), .o(n_3397) );
in01f80 g761024 ( .a(n_19350), .o(n_19375) );
no02f80 g771670 ( .a(n_9065), .b(n_44511), .o(n_10283) );
in01f80 g736640 ( .a(n_43156), .o(n_43118) );
na02f80 g750515 ( .a(n_30477), .b(n_30476), .o(n_30478) );
ao12f80 g739391 ( .a(n_40773), .b(FE_OCPN897_n_44776), .c(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n_41279) );
in01f80 g749609 ( .a(n_30285), .o(n_30286) );
no02f80 g758061 ( .a(n_22845), .b(n_22734), .o(n_22880) );
oa12f80 g774523 ( .a(n_6624), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_26_), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_25_), .o(n_6830) );
na02f80 g780402 ( .a(n_804), .b(n_45814), .o(n_876) );
in01f80 FE_RC_1850_0 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_1_), .o(FE_RN_564_0) );
na02f80 g767975 ( .a(n_12811), .b(n_12810), .o(n_13177) );
in01f80 newInst_1955 ( .a(newNet_855), .o(newNet_1955) );
ao12f80 g741561 ( .a(n_38670), .b(n_38669), .c(n_38668), .o(n_38712) );
ao12f80 g756621 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_25_), .c(delay_add_ln22_unr14_stage6_stallmux_q_24_), .o(n_23815) );
no02f80 g743560 ( .a(n_36148), .b(n_36504), .o(n_36547) );
no02f80 g760094 ( .a(n_20429), .b(FE_OCP_RBN1700_n_19353), .o(n_20534) );
in01f80 g736844 ( .a(n_43072), .o(n_43050) );
na02f80 g750035 ( .a(n_30007), .b(n_30049), .o(n_30139) );
no02f80 g750311 ( .a(n_30721), .b(n_30720), .o(n_30722) );
ao12f80 g781125 ( .a(n_218), .b(n_222), .c(n_217), .o(n_399) );
in01f80 g777198 ( .a(n_3635), .o(n_3579) );
na02f80 g736961 ( .a(n_43120), .b(n_43251), .o(n_43324) );
in01f80 g749273 ( .a(n_30739), .o(n_30763) );
no02f80 g739429 ( .a(FE_OCPN932_n_40736), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_21_), .o(n_40773) );
na02f80 g776216 ( .a(n_3993), .b(n_4668), .o(n_4795) );
in01f80 FE_OCP_DRV_C1583_n_30917 ( .a(n_30917), .o(FE_OCP_DRV_N1583_n_30917) );
ao12f80 g749659 ( .a(n_31542), .b(n_31459), .c(n_31311), .o(n_31543) );
no02f80 g776911 ( .a(n_3776), .b(n_3862), .o(n_3887) );
in01f80 g754597 ( .a(n_26793), .o(n_26707) );
in01f80 FE_RC_163_0 ( .a(n_11998), .o(FE_RN_49_0) );
in01f80 FE_RC_603_0 ( .a(FE_RN_191_0), .o(n_40736) );
no02f80 g780927 ( .a(n_403), .b(n_447), .o(n_452) );
no02f80 g762620 ( .a(FE_OCP_RBN2147_FE_OCPN861_n_45450), .b(delay_xor_ln21_unr12_stage5_stallmux_q_16_), .o(n_18137) );
na02f80 g761074 ( .a(n_19309), .b(n_19308), .o(n_19310) );
ao22s80 FE_RC_3707_0 ( .a(n_43542), .b(n_43875), .c(n_43541), .d(n_43874), .o(n_43902) );
in01f80 FE_OCP_RBC3714_n_31466 ( .a(FE_OCP_RBN3712_n_31466), .o(FE_OCP_RBN3714_n_31466) );
na02f80 g758058 ( .a(n_22920), .b(n_22951), .o(n_23342) );
in01f80 g743626 ( .a(n_36457), .o(n_36458) );
no02f80 g753971 ( .a(FE_OCP_RBN2882_n_26318), .b(n_23564), .o(n_26353) );
na02f80 g758721 ( .a(n_21656), .b(n_20059), .o(n_21687) );
in01f80 g762433 ( .a(n_18005), .o(n_18006) );
no02f80 g768877 ( .a(n_12124), .b(n_11871), .o(n_11872) );
ms00f80 cos_out_reg_29_ ( .ck(newNet_3702), .d(n_43897), .o(cos_out_29) );
no02f80 g743417 ( .a(n_37747), .b(n_36978), .o(n_37830) );
no02f80 g765338 ( .a(FE_OCP_RBN3621_n_15135), .b(n_14397), .o(n_15491) );
no02f80 g754357 ( .a(n_25731), .b(n_25824), .o(n_25765) );
oa12f80 g759704 ( .a(n_21406), .b(n_21751), .c(n_21750), .o(n_21799) );
na02f80 g748683 ( .a(n_31359), .b(n_31076), .o(n_31398) );
oa12f80 g750495 ( .a(n_30478), .b(n_30477), .c(n_30476), .o(n_31256) );
in01f80 g746518 ( .a(n_34777), .o(n_34721) );
ms00f80 delay_sub_ln23_0_unr19_stage7_stallmux_q_reg ( .ck(newNet_1666), .d(n_26896), .o(n_27014) );
no03m80 g757095 ( .a(n_23175), .b(n_23176), .c(delay_add_ln22_unr14_stage6_stallmux_q_7_), .o(n_23251) );
ao12f80 g742746 ( .a(n_37222), .b(n_37291), .c(n_37288), .o(n_37323) );
na02f80 g736812 ( .a(n_43424), .b(n_46935), .o(n_43313) );
ao12f80 g772225 ( .a(n_8487), .b(n_8632), .c(n_8535), .o(n_8711) );
in01f80 newInst_1467 ( .a(newNet_1466), .o(newNet_1467) );
in01f80 newInst_3696 ( .a(newNet_3695), .o(newNet_3696) );
oa12f80 g754504 ( .a(n_26932), .b(n_26931), .c(n_26930), .o(n_26996) );
na02f80 g773775 ( .a(n_7159), .b(n_7078), .o(n_7160) );
na02f80 g743833 ( .a(n_35920), .b(n_35919), .o(n_35921) );
in01f80 g745687 ( .a(n_34297), .o(n_34285) );
no02f80 g757546 ( .a(n_23298), .b(n_23295), .o(n_23299) );
ao12f80 g764932 ( .a(n_16066), .b(n_15874), .c(n_16246), .o(n_16353) );
na02f80 g777038 ( .a(n_3634), .b(n_3440), .o(n_3758) );
na02f80 FE_RC_4229_0 ( .a(n_13476), .b(n_15001), .o(FE_RN_1856_0) );
oa12f80 g768403 ( .a(n_12461), .b(n_12404), .c(FE_OCPN1002_n_45660), .o(n_12760) );
in01f80 newInst_2532 ( .a(newNet_2531), .o(newNet_2532) );
no02f80 g774077 ( .a(n_6723), .b(n_6653), .o(n_6777) );
no02f80 g773618 ( .a(n_7381), .b(n_7173), .o(n_7420) );
no02f80 g772397 ( .a(n_8518), .b(n_8027), .o(n_8606) );
in01f80 newInst_1837 ( .a(newNet_1836), .o(newNet_1837) );
no02f80 g740025 ( .a(n_40006), .b(FE_OCP_RBN3717_n_39913), .o(n_40154) );
in01f80 g769971 ( .a(n_10965), .o(n_10966) );
na02f80 FE_RC_2130_0 ( .a(n_15036), .b(FE_RN_743_0), .o(n_15321) );
oa22f80 FE_RC_706_0 ( .a(n_38214), .b(n_38520), .c(n_38215), .d(n_38519), .o(n_38583) );
in01f80 FE_OCP_RBC1847_n_22068 ( .a(FE_OCP_RBN1846_n_22068), .o(FE_OCP_RBN1847_n_22068) );
in01f80 g756602 ( .a(n_23580), .o(n_23663) );
no02f80 g764585 ( .a(n_16144), .b(FE_OCPN1734_n_16143), .o(n_16271) );
in01f80 g736569 ( .a(n_43571), .o(n_43572) );
ao12f80 g750168 ( .a(n_29791), .b(n_29790), .c(n_29789), .o(n_29842) );
no02f80 g747131 ( .a(n_32926), .b(n_32967), .o(n_32983) );
oa22f80 g752853 ( .a(n_27988), .b(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .c(n_27762), .d(delay_sub_ln23_0_unr20_stage7_stallmux_q_3_), .o(n_28021) );
in01f80 g744971 ( .a(n_34978), .o(n_34996) );
na02f80 g739110 ( .a(n_40946), .b(n_40798), .o(n_40997) );
no02f80 g773458 ( .a(n_7522), .b(n_7521), .o(n_7531) );
no02f80 g755988 ( .a(n_24165), .b(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24185) );
in01f80 g740195 ( .a(n_40214), .o(n_40215) );
oa12f80 g756288 ( .a(n_24008), .b(n_24588), .c(n_24074), .o(n_24676) );
in01f80 g774848 ( .a(n_6341), .o(n_6342) );
oa22f80 g784558 ( .a(FE_OFN800_n_46285), .b(n_10959), .c(FE_OCP_RBN3709_n_46337), .d(n_10928), .o(n_46379) );
na02f80 g764621 ( .a(n_15951), .b(n_14588), .o(n_16048) );
na02f80 g759640 ( .a(n_21752), .b(n_21831), .o(n_21832) );
na02f80 g760509 ( .a(n_20044), .b(n_19994), .o(n_20073) );
in01f80 g773243 ( .a(n_7735), .o(n_7736) );
in01f80 g740021 ( .a(n_40120), .o(n_40148) );
no02f80 g777796 ( .a(n_3328), .b(n_3321), .o(n_3405) );
na02f80 g775584 ( .a(n_5308), .b(n_4182), .o(n_5451) );
in01f80 g773970 ( .a(n_7008), .o(n_7009) );
no02f80 g760870 ( .a(n_19450), .b(n_19552), .o(n_19553) );
no02f80 g740140 ( .a(n_39816), .b(n_39785), .o(n_39845) );
no02f80 g766594 ( .a(n_13931), .b(FE_OCP_RBN2363_n_13785), .o(n_13952) );
in01f80 fopt783571 ( .a(n_2408), .o(n_45194) );
in01f80 g760366 ( .a(n_20209), .o(n_20210) );
na02f80 g773506 ( .a(n_7508), .b(n_7117), .o(n_7560) );
na02f80 g768888 ( .a(n_12088), .b(n_12087), .o(n_12089) );
in01f80 newInst_1268 ( .a(newNet_1182), .o(newNet_1268) );
in01f80 g760731 ( .a(n_19639), .o(n_19658) );
no02f80 g764386 ( .a(n_16632), .b(n_16062), .o(n_16677) );
no02f80 g744398 ( .a(n_35501), .b(FE_OCP_DRV_N1582_n_35500), .o(n_35516) );
no02f80 g754577 ( .a(n_25404), .b(n_25212), .o(n_25430) );
in01f80 newInst_1608 ( .a(newNet_1607), .o(newNet_1608) );
in01f80 FE_OCP_RBC1194_n_22542 ( .a(n_22542), .o(FE_OCP_RBN1194_n_22542) );
in01f80 g756875 ( .a(n_24063), .o(n_24046) );
in01f80 g744487 ( .a(n_35429), .o(n_35430) );
oa12f80 g775106 ( .a(n_6066), .b(n_6127), .c(n_6069), .o(n_6128) );
in01f80 g772305 ( .a(n_8548), .o(n_8549) );
in01f80 g776140 ( .a(n_4990), .o(n_5107) );
ao12f80 g746521 ( .a(n_34473), .b(n_34697), .c(n_34696), .o(n_34698) );
na02f80 g774968 ( .a(n_6125), .b(n_5980), .o(n_6156) );
na02f80 g776455 ( .a(n_4542), .b(n_4688), .o(n_4753) );
na02f80 g744131 ( .a(n_35590), .b(n_35615), .o(n_35638) );
na02f80 g778025 ( .a(n_3008), .b(n_2985), .o(n_2986) );
ao22s80 FE_RC_741_0 ( .a(FE_OCPN1011_n_7802), .b(FE_OCP_RBN2476_n_8599), .c(n_8599), .d(FE_OCP_RBN3468_n_7886), .o(n_8727) );
na04m80 g762179 ( .a(n_18813), .b(n_18841), .c(n_18840), .d(n_18839), .o(n_18931) );
oa12f80 g768440 ( .a(n_12251), .b(n_12412), .c(n_12186), .o(n_12467) );
in01f80 g769072 ( .a(n_11775), .o(n_11665) );
in01f80 g780949 ( .a(n_420), .o(n_580) );
no02f80 g741966 ( .a(n_37957), .b(n_38016), .o(n_38017) );
in01f80 FE_OCP_RBC1724_n_21004 ( .a(FE_OCP_RBN1723_n_21004), .o(FE_OCP_RBN1724_n_21004) );
oa12f80 g753612 ( .a(n_26625), .b(n_26624), .c(n_26623), .o(n_26693) );
in01f80 newInst_3465 ( .a(newNet_3464), .o(newNet_3465) );
oa22f80 FE_RC_3343_0 ( .a(n_25562), .b(n_25845), .c(n_25563), .d(n_25846), .o(n_25934) );
na02f80 g739579 ( .a(n_40615), .b(n_44610), .o(n_40647) );
no02f80 g738293 ( .a(n_41865), .b(n_41480), .o(n_41844) );
in01f80 FE_OCPC981_n_31961 ( .a(FE_OCP_RBN3085_n_31819), .o(FE_OCPN981_n_31961) );
in01f80 g762126 ( .a(n_18218), .o(n_18219) );
in01f80 g747187 ( .a(n_32903), .o(n_32904) );
no02f80 g777394 ( .a(n_3549), .b(n_3548), .o(n_3576) );
in01f80 newInst_2389 ( .a(newNet_2388), .o(newNet_2389) );
in01f80 g761118 ( .a(n_19301), .o(n_20430) );
na02f80 g777120 ( .a(n_3696), .b(n_3670), .o(n_3802) );
na02f80 g765937 ( .a(n_14774), .b(FE_OCP_RBN2272_n_13489), .o(n_14851) );
no02f80 g775615 ( .a(n_5477), .b(n_5476), .o(n_5506) );
no02f80 g771301 ( .a(n_9785), .b(n_9784), .o(n_9905) );
na02f80 g743012 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_37075) );
in01f80 g772552 ( .a(FE_OCP_RBN2440_n_8402), .o(n_8452) );
na02f80 g767863 ( .a(n_12773), .b(n_12723), .o(n_12793) );
na02f80 g751612 ( .a(n_29249), .b(n_29103), .o(n_29250) );
no03m80 FE_RC_645_0 ( .a(FE_OCP_RBN3373_n_6745), .b(n_6716), .c(n_6710), .o(n_6711) );
in01f80 g763438 ( .a(n_17027), .o(n_17069) );
no02f80 g746943 ( .a(n_32857), .b(n_32275), .o(n_32920) );
in01f80 g778362 ( .a(n_2583), .o(n_2584) );
in01f80 newInst_2626 ( .a(newNet_973), .o(newNet_2626) );
na02f80 g748186 ( .a(n_31503), .b(FE_OCP_RBN3712_n_31466), .o(n_31562) );
in01f80 fopt784455 ( .a(n_37082), .o(n_46256) );
no02f80 g757491 ( .a(FE_OCP_RBN3823_n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_6_), .o(n_23227) );
no02f80 g775617 ( .a(n_5307), .b(FE_OCP_RBN2734_n_4219), .o(n_5370) );
na02f80 g759990 ( .a(FE_OCP_RBN3840_n_19513), .b(n_20533), .o(n_20581) );
ao12f80 g776869 ( .a(n_3975), .b(n_4209), .c(n_4208), .o(n_4210) );
na02f80 g774966 ( .a(n_6186), .b(n_6234), .o(n_6203) );
na02f80 FE_RC_3831_0 ( .a(FE_RN_1669_0), .b(FE_RN_1670_0), .o(FE_RN_1671_0) );
in01f80 g752985 ( .a(n_27276), .o(n_27310) );
oa22f80 FE_RC_3915_0 ( .a(n_22270), .b(n_22639), .c(n_22307), .d(FE_OCP_RBN1850_n_22639), .o(n_22829) );
oa22f80 FE_RC_3412_0 ( .a(n_22961), .b(n_22631), .c(n_20252), .d(n_22611), .o(n_22704) );
no02f80 g737194 ( .a(n_42947), .b(delay_sub_ln23_0_unr30_stage10_stallmux_q), .o(n_42965) );
oa22f80 FE_RC_193_0 ( .a(n_17385), .b(n_17693), .c(n_17384), .d(n_17658), .o(n_17812) );
in01f80 newInst_118 ( .a(newNet_117), .o(newNet_118) );
ao12f80 g779187 ( .a(n_1630), .b(n_44811), .c(n_1586), .o(n_1885) );
in01f80 g751194 ( .a(n_29974), .o(n_29975) );
in01f80 g761467 ( .a(n_20254), .o(n_20009) );
oa12f80 g776825 ( .a(n_3586), .b(n_3724), .c(n_3539), .o(n_3822) );
in01f80 g753459 ( .a(n_27586), .o(n_27587) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_12_ ( .ck(newNet_668), .d(n_46362), .o(delay_xor_ln21_unr9_stage4_stallmux_q_12_) );
ao22s80 g752217 ( .a(n_28479), .b(n_28315), .c(n_28480), .d(n_28314), .o(n_28987) );
no02f80 g776317 ( .a(n_4429), .b(n_4182), .o(n_4550) );
in01f80 g776746 ( .a(n_4011), .o(n_4012) );
in01f80 FE_OCP_RBC2724_n_4219 ( .a(n_4219), .o(FE_OCP_RBN2724_n_4219) );
no02f80 FE_RC_2652_0 ( .a(n_12323), .b(n_12542), .o(FE_RN_1106_0) );
no02f80 g749550 ( .a(n_30357), .b(n_30076), .o(n_30388) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_24_ ( .ck(newNet_1604), .d(n_27447), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_24_) );
in01f80 FE_OCP_RBC3332_n_44962 ( .a(n_44962), .o(FE_OCP_RBN3332_n_44962) );
in01f80 newInst_1121 ( .a(newNet_1120), .o(newNet_1121) );
na02f80 g776321 ( .a(n_4771), .b(n_4171), .o(n_4846) );
ao22s80 FE_RC_1891_0 ( .a(n_45312), .b(FE_RN_589_0), .c(n_45311), .d(n_23000), .o(n_23193) );
na02f80 g751327 ( .a(n_29601), .b(n_29581), .o(n_29582) );
no02f80 g740322 ( .a(n_39733), .b(n_39742), .o(n_39770) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_29_ ( .ck(newNet_1484), .d(n_32379), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_29_) );
in01f80 g773380 ( .a(n_7590), .o(n_7591) );
in01f80 g780354 ( .a(n_947), .o(n_1019) );
no02f80 g762106 ( .a(n_46972), .b(n_16830), .o(n_18263) );
oa22f80 FE_RC_3266_0 ( .a(FE_OFN803_n_46285), .b(n_12068), .c(FE_OCP_RBN3043_n_46337), .d(n_12064), .o(n_46354) );
oa12f80 g756404 ( .a(n_23843), .b(n_24011), .c(delay_add_ln22_unr14_stage6_stallmux_q_30_), .o(n_24012) );
in01f80 newInst_428 ( .a(newNet_168), .o(newNet_428) );
in01f80 FE_OCP_RBC3660_n_15233 ( .a(n_15233), .o(FE_OCP_RBN3660_n_15233) );
oa22f80 g763861 ( .a(n_46979), .b(n_17584), .c(n_16634), .d(n_16338), .o(n_16700) );
ao22s80 FE_RC_853_0 ( .a(n_23917), .b(n_24424), .c(n_23918), .d(n_24423), .o(n_24518) );
ao12f80 g737485 ( .a(n_42247), .b(n_42555), .c(n_42259), .o(n_42639) );
in01f80 FE_OCP_RBC1174_n_18981 ( .a(n_18981), .o(FE_OCP_RBN1174_n_18981) );
no02f80 g742677 ( .a(n_37497), .b(n_37496), .o(n_37498) );
na02f80 g746482 ( .a(n_34865), .b(n_34811), .o(n_34866) );
na02f80 g772417 ( .a(n_8686), .b(n_8652), .o(n_8774) );
no02f80 g760124 ( .a(n_20332), .b(n_20369), .o(n_20370) );
oa22f80 g784348 ( .a(FE_OFN774_n_46137), .b(n_6280), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_6301), .o(n_46154) );
in01f80 g753134 ( .a(n_27496), .o(n_27497) );
in01f80 newInst_1378 ( .a(newNet_1377), .o(newNet_1378) );
in01f80 g771705 ( .a(n_9234), .o(n_9235) );
oa12f80 g750929 ( .a(n_30208), .b(n_30130), .c(n_29944), .o(n_30233) );
na02f80 g776220 ( .a(n_4630), .b(n_4699), .o(n_4743) );
no02f80 g766128 ( .a(n_14595), .b(n_14572), .o(n_14657) );
no02f80 g776624 ( .a(n_3981), .b(n_3029), .o(n_4055) );
no02f80 g778303 ( .a(n_2586), .b(n_2557), .o(n_2718) );
in01f80 g775452 ( .a(n_5526), .o(n_5540) );
oa22f80 g744877 ( .a(n_36403), .b(n_35886), .c(n_36404), .d(n_35887), .o(n_36453) );
na02f80 g739919 ( .a(n_40231), .b(n_39974), .o(n_40260) );
in01f80 g738493 ( .a(n_41701), .o(n_41670) );
in01f80 g771769 ( .a(n_9097), .o(n_9127) );
in01f80 g759263 ( .a(n_20984), .o(n_21011) );
na02f80 g765528 ( .a(n_15719), .b(n_15711), .o(n_15784) );
no02f80 g767807 ( .a(n_12764), .b(n_13017), .o(n_13350) );
in01f80 newInst_3585 ( .a(newNet_3584), .o(newNet_3585) );
na02f80 g752672 ( .a(n_28261), .b(n_28132), .o(n_28262) );
na02f80 g737752 ( .a(n_42293), .b(n_42258), .o(n_42357) );
in01f80 g774046 ( .a(n_7196), .o(n_7197) );
in01f80 g750075 ( .a(n_30216), .o(n_30261) );
na02f80 g740277 ( .a(n_39857), .b(n_40045), .o(n_39858) );
in01f80 FE_OCPC896_n_44776 ( .a(n_44776), .o(FE_OCPN896_n_44776) );
na02f80 g780597 ( .a(n_713), .b(n_731), .o(n_771) );
na02f80 g745015 ( .a(n_45185), .b(n_34429), .o(n_34833) );
in01f80 g761536 ( .a(n_18799), .o(n_18871) );
in01f80 newInst_2816 ( .a(newNet_376), .o(newNet_2816) );
in01f80 g770522 ( .a(n_10499), .o(n_10500) );
in01f80 g776847 ( .a(n_4254), .o(n_4255) );
in01f80 g777814 ( .a(n_3318), .o(n_3270) );
na02f80 g776230 ( .a(n_4812), .b(n_4345), .o(n_4933) );
na02f80 g741469 ( .a(n_38792), .b(n_38791), .o(n_38802) );
ao12f80 g760314 ( .a(n_19989), .b(n_20835), .c(n_20053), .o(n_20929) );
no02f80 g741876 ( .a(n_38191), .b(n_38062), .o(n_38262) );
na02f80 g748812 ( .a(n_32420), .b(n_32419), .o(n_32803) );
in01f80 g768544 ( .a(n_12346), .o(n_12347) );
ao22s80 FE_RC_1812_0 ( .a(FE_RN_537_0), .b(n_11909), .c(FE_OCP_RBN2138_n_11909), .d(n_11770), .o(n_12128) );
in01f80 newInst_37 ( .a(newNet_1), .o(newNet_37) );
oa22f80 g784550 ( .a(FE_OFN801_n_46285), .b(n_11307), .c(FE_OCP_RBN3044_n_46337), .d(n_11282), .o(n_46371) );
na02f80 g775988 ( .a(n_4957), .b(n_4763), .o(n_5002) );
oa12f80 g780808 ( .a(n_381), .b(n_380), .c(n_379), .o(n_1108) );
ao12f80 g736388 ( .a(n_43681), .b(n_43822), .c(n_43522), .o(n_43842) );
in01f80 g756713 ( .a(n_23595), .o(n_23596) );
in01f80 newInst_613 ( .a(newNet_612), .o(newNet_613) );
ao12f80 g744445 ( .a(n_35227), .b(n_35475), .c(n_35148), .o(n_35487) );
oa22f80 g784565 ( .a(FE_OFN801_n_46285), .b(n_11411), .c(FE_OCP_RBN3044_n_46337), .d(n_11396), .o(n_46386) );
ao12f80 g737356 ( .a(n_42551), .b(n_42808), .c(n_42530), .o(n_42864) );
no02f80 g757340 ( .a(n_23105), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_3_), .o(n_23127) );
no02f80 g768987 ( .a(n_11656), .b(n_47279), .o(n_11729) );
ao22s80 g765408 ( .a(n_16245), .b(n_15788), .c(n_15874), .d(n_14112), .o(n_16346) );
ao22s80 g761646 ( .a(n_19540), .b(n_18838), .c(n_19526), .d(n_18837), .o(n_19986) );
in01f80 g747219 ( .a(n_32755), .o(n_32756) );
na02f80 FE_RC_4035_0 ( .a(n_21200), .b(FE_RN_1752_0), .o(n_21394) );
in01f80 g754756 ( .a(n_25365), .o(n_25403) );
no02f80 g762243 ( .a(n_18835), .b(n_18834), .o(n_18836) );
in01f80 FE_OCP_RBC1689_n_18986 ( .a(FE_OCP_RBN1687_n_18986), .o(FE_OCP_RBN1689_n_18986) );
in01f80 g756345 ( .a(n_24478), .o(n_24587) );
no02f80 g740071 ( .a(n_40112), .b(n_40111), .o(n_40139) );
in01f80 g775298 ( .a(n_5691), .o(n_5692) );
na02f80 g741464 ( .a(n_44165), .b(n_38730), .o(n_38789) );
oa12f80 g774174 ( .a(n_6673), .b(n_6672), .c(n_6671), .o(n_7673) );
oa22f80 FE_RC_1238_0 ( .a(n_44570), .b(FE_OCP_RBN3557_n_8687), .c(n_8687), .d(n_44568), .o(n_9001) );
in01f80 newInst_864 ( .a(newNet_570), .o(newNet_864) );
in01f80 g776239 ( .a(n_4894), .o(n_4895) );
na02f80 g757937 ( .a(n_22924), .b(n_22851), .o(n_22925) );
ao12f80 g757362 ( .a(n_22972), .b(n_44084), .c(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .o(n_22998) );
no02f80 g777229 ( .a(n_3741), .b(n_3714), .o(n_3899) );
in01f80 g772930 ( .a(n_7936), .o(n_7937) );
in01f80 FE_RC_2887_0 ( .a(FE_RN_1250_0), .o(n_14625) );
no02f80 FE_RC_2558_0 ( .a(n_6698), .b(n_6896), .o(FE_RN_1048_0) );
na02f80 g759718 ( .a(n_20755), .b(n_20787), .o(n_20838) );
ao12f80 g773955 ( .a(n_7271), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .o(n_7289) );
in01f80 g754570 ( .a(n_26790), .o(n_26791) );
in01f80 newInst_3129 ( .a(newNet_3128), .o(newNet_3129) );
in01f80 g757409 ( .a(n_23095), .o(n_23096) );
in01f80 g741171 ( .a(n_38885), .o(n_38922) );
ao12f80 g738133 ( .a(n_42019), .b(n_42018), .c(n_42017), .o(n_42321) );
in01f80 g745229 ( .a(n_36250), .o(n_36251) );
no02f80 g741000 ( .a(n_39063), .b(n_38993), .o(n_39064) );
na02f80 g765278 ( .a(n_15668), .b(n_15783), .o(n_15785) );
in01f80 g761731 ( .a(n_18714), .o(n_18715) );
in01f80 FE_OCP_RBC1129_n_24179 ( .a(n_24179), .o(FE_OCP_RBN1129_n_24179) );
in01f80 g745727 ( .a(n_35432), .o(n_35451) );
na02f80 g750372 ( .a(n_29739), .b(n_29737), .o(n_29727) );
in01f80 g749403 ( .a(delay_sub_ln23_0_unr24_stage8_stallmux_q_9_), .o(n_32034) );
oa12f80 g775562 ( .a(n_5710), .b(n_5638), .c(n_5709), .o(n_5739) );
in01f80 FE_OCP_RBC2447_n_14114 ( .a(n_14114), .o(FE_OCP_RBN2447_n_14114) );
na02f80 g764323 ( .a(n_16677), .b(n_15973), .o(n_16722) );
oa12f80 g762059 ( .a(n_18105), .b(n_18247), .c(n_18067), .o(n_18267) );
ao12f80 g743547 ( .a(n_37612), .b(n_36727), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37699) );
in01f80 g740629 ( .a(n_39592), .o(n_39593) );
no02f80 g738739 ( .a(n_41483), .b(n_41142), .o(n_41529) );
na02f80 g743958 ( .a(n_36303), .b(n_35699), .o(n_36318) );
no02f80 g741065 ( .a(n_38956), .b(FE_OCP_RBN2553_n_44921), .o(n_39054) );
no02f80 FE_RC_3521_0 ( .a(n_34490), .b(n_34514), .o(FE_RN_1521_0) );
no02f80 g770340 ( .a(n_10597), .b(n_10508), .o(n_10660) );
ao12f80 g766532 ( .a(n_13922), .b(n_13994), .c(n_14064), .o(n_14026) );
in01f80 g757054 ( .a(n_23704), .o(n_23672) );
in01f80 g768136 ( .a(n_12721), .o(n_13004) );
in01f80 g766248 ( .a(n_14591), .o(n_14592) );
oa22f80 g739852 ( .a(n_40400), .b(n_40317), .c(n_40401), .d(n_40316), .o(n_40441) );
in01f80 FE_RC_1007_0 ( .a(n_17355), .o(FE_RN_291_0) );
na02f80 g754724 ( .a(FE_OCP_RBN2966_n_26231), .b(n_26542), .o(n_26708) );
in01f80 g747584 ( .a(n_32382), .o(n_32383) );
in01f80 newInst_734 ( .a(newNet_733), .o(newNet_734) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_18_ ( .ck(newNet_1122), .d(n_10840), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_18_) );
no02f80 g746273 ( .a(n_33589), .b(n_33588), .o(n_33591) );
na02f80 g764268 ( .a(n_16453), .b(n_16454), .o(n_16512) );
oa12f80 g751421 ( .a(n_28958), .b(n_29177), .c(n_28878), .o(n_29226) );
in01f80 g775376 ( .a(n_5717), .o(n_5754) );
na02f80 g744569 ( .a(n_35329), .b(n_35223), .o(n_35387) );
na02f80 g763837 ( .a(n_16640), .b(n_16656), .o(n_16703) );
ao12f80 g779648 ( .a(n_1451), .b(n_1452), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .o(n_1482) );
na03f80 g743597 ( .a(n_37541), .b(n_37475), .c(n_37540), .o(n_37543) );
in01f80 g768233 ( .a(n_12721), .o(n_12739) );
no02f80 g746967 ( .a(FE_OCP_RBN2168_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .o(n_33158) );
in01f80 g780612 ( .a(n_664), .o(n_687) );
no02f80 g743946 ( .a(n_47267), .b(n_36036), .o(n_36037) );
na02f80 g750555 ( .a(n_29496), .b(n_29495), .o(n_29497) );
ao12f80 g754815 ( .a(n_25246), .b(n_25247), .c(n_25144), .o(n_25336) );
in01f80 g765376 ( .a(n_16300), .o(n_16301) );
in01f80 g739731 ( .a(n_40491), .o(n_40492) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_0_ ( .ck(newNet_2226), .d(n_46055), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_0_) );
in01f80 newInst_2436 ( .a(newNet_962), .o(newNet_2436) );
in01f80 g771310 ( .a(n_9639), .o(n_9686) );
in01f80 g741312 ( .a(n_38852), .o(n_39246) );
ao12f80 g769740 ( .a(n_10211), .b(n_11267), .c(n_11266), .o(n_11268) );
na02f80 g767981 ( .a(n_12765), .b(n_12701), .o(n_12786) );
in01f80 FE_RC_4220_0 ( .a(n_30018), .o(FE_RN_1849_0) );
ao22s80 FE_RC_1548_0 ( .a(n_23029), .b(n_23263), .c(n_23030), .d(n_23246), .o(n_23347) );
ao12f80 g751361 ( .a(n_28320), .b(n_28536), .c(n_28344), .o(n_28612) );
na02f80 g769822 ( .a(n_11029), .b(n_44498), .o(n_11065) );
in01f80 FE_OCP_RBC2819_n_4872 ( .a(n_4872), .o(FE_OCP_RBN2819_n_4872) );
no02f80 g742828 ( .a(n_37276), .b(n_37110), .o(n_37368) );
no02f80 g753978 ( .a(n_26212), .b(n_26186), .o(n_26294) );
in01f80 g737635 ( .a(n_42762), .o(n_42763) );
na02f80 g775015 ( .a(n_6147), .b(n_6001), .o(n_6179) );
in01f80 newInst_3730 ( .a(newNet_3729), .o(newNet_3730) );
na02f80 g777928 ( .a(n_3075), .b(n_2408), .o(n_3107) );
in01f80 g765834 ( .a(n_14929), .o(n_14930) );
no02f80 g754372 ( .a(n_26941), .b(n_26232), .o(n_26646) );
in01f80 g752413 ( .a(n_27781), .o(n_27752) );
no03m80 FE_RC_700_0 ( .a(n_40655), .b(n_40649), .c(n_40637), .o(n_40659) );
in01f80 newInst_2033 ( .a(newNet_2032), .o(newNet_2033) );
in01f80 g780619 ( .a(n_985), .o(n_986) );
na02f80 g749036 ( .a(n_31004), .b(n_31003), .o(n_31005) );
oa12f80 g757523 ( .a(n_22305), .b(n_22720), .c(n_22221), .o(n_22721) );
in01f80 g749219 ( .a(n_30871), .o(n_30906) );
na02f80 g766724 ( .a(n_13778), .b(n_13777), .o(n_13779) );
na02f80 FE_RC_1045_0 ( .a(FE_RN_303_0), .b(FE_RN_304_0), .o(FE_RN_305_0) );
na02f80 g747210 ( .a(n_32671), .b(n_32670), .o(n_32735) );
na02f80 g769205 ( .a(n_11798), .b(n_11797), .o(n_12153) );
in01f80 newInst_2103 ( .a(newNet_379), .o(newNet_2103) );
oa22f80 FE_RC_1428_0 ( .a(n_22801), .b(n_22715), .c(n_22793), .d(n_22670), .o(n_22770) );
in01f80 newInst_1963 ( .a(newNet_1962), .o(newNet_1963) );
in01f80 g747036 ( .a(n_32860), .o(n_32892) );
in01f80 g764272 ( .a(n_16407), .o(n_16434) );
in01f80 newInst_2302 ( .a(newNet_46), .o(newNet_2302) );
no02f80 g749925 ( .a(n_30318), .b(n_30294), .o(n_30320) );
oa12f80 g767399 ( .a(n_13522), .b(n_13521), .c(n_13520), .o(n_13975) );
in01f80 g774382 ( .a(n_6922), .o(n_6923) );
no02f80 g763070 ( .a(n_17452), .b(n_17451), .o(n_17453) );
in01f80 newInst_2656 ( .a(newNet_2655), .o(newNet_2656) );
no02f80 g739452 ( .a(n_44769), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_28_), .o(n_40901) );
in01f80 FE_RC_2245_0 ( .a(n_37205), .o(FE_RN_824_0) );
oa12f80 g744155 ( .a(n_46223), .b(n_46222), .c(n_36898), .o(n_36882) );
no02f80 g755142 ( .a(n_25373), .b(FE_OCP_RBN2421_n_24505), .o(n_25644) );
na02f80 g757814 ( .a(n_23183), .b(n_23119), .o(n_23182) );
in01f80 g738501 ( .a(n_41743), .o(n_41744) );
in01f80 newInst_1634 ( .a(newNet_256), .o(newNet_1634) );
in01f80 g778659 ( .a(n_2425), .o(n_2426) );
in01f80 newInst_3687 ( .a(newNet_3686), .o(newNet_3687) );
in01f80 g780464 ( .a(n_821), .o(n_805) );
in01f80 FE_RC_1331_0 ( .a(n_39426), .o(FE_RN_394_0) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_22_ ( .ck(newNet_3527), .d(n_22709), .o(delay_add_ln22_unr14_stage6_stallmux_q_22_) );
na02f80 FE_RC_2316_0 ( .a(FE_RN_880_0), .b(n_36476), .o(n_36513) );
oa12f80 g784616 ( .a(n_42567), .b(n_42552), .c(n_42314), .o(n_46944) );
in01f80 g773757 ( .a(n_45889), .o(n_7193) );
in01f80 newInst_2602 ( .a(newNet_995), .o(newNet_2602) );
no02f80 g747984 ( .a(n_33085), .b(n_33084), .o(n_33086) );
na02f80 g760433 ( .a(n_20033), .b(n_20032), .o(n_20034) );
in01f80 g743304 ( .a(n_36725), .o(n_36739) );
oa12f80 g778930 ( .a(n_1751), .b(n_2143), .c(n_1801), .o(n_2170) );
oa22f80 FE_RC_1114_0 ( .a(n_38198), .b(n_38532), .c(n_38197), .d(n_38531), .o(n_38586) );
in01f80 g779334 ( .a(n_1701), .o(n_1702) );
in01f80 FE_OCP_RBC2221_n_13010 ( .a(n_13010), .o(FE_OCP_RBN2221_n_13010) );
in01f80 g764452 ( .a(n_16272), .o(n_16364) );
no02f80 g771599 ( .a(n_9168), .b(n_9203), .o(n_9268) );
no02f80 g760623 ( .a(n_19810), .b(n_19809), .o(n_19811) );
na02f80 g742392 ( .a(n_37745), .b(FE_OCPN1778_n_37744), .o(n_37799) );
no02f80 FE_RC_2440_0 ( .a(n_29915), .b(n_30298), .o(n_30375) );
no02f80 g746343 ( .a(n_33473), .b(n_33019), .o(n_33504) );
oa22f80 g742963 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_31_), .c(n_37082), .d(n_36650), .o(n_37054) );
na02f80 FE_RC_3483_0 ( .a(n_37133), .b(FE_RN_1497_0), .o(FE_RN_1498_0) );
in01f80 g745211 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .o(n_36353) );
in01f80 g764161 ( .a(n_16557), .o(n_16558) );
oa12f80 g752977 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n_28016) );
na02f80 g760896 ( .a(n_19460), .b(n_19427), .o(n_19585) );
no02f80 g769990 ( .a(n_10826), .b(n_10860), .o(n_10919) );
na02f80 g761921 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_23_), .o(n_18400) );
na02f80 g768435 ( .a(n_12390), .b(n_12431), .o(n_12666) );
in01f80 g742532 ( .a(n_37598), .o(n_37623) );
in01f80 newInst_983 ( .a(newNet_982), .o(newNet_983) );
ao22s80 g736479 ( .a(n_43713), .b(n_43586), .c(n_43712), .d(n_43585), .o(n_43748) );
in01f80 FE_RC_3485_0 ( .a(FE_RN_1500_0), .o(FE_RN_1499_0) );
in01f80 FE_RC_4066_0 ( .a(n_26516), .o(FE_RN_1770_0) );
no02f80 g742881 ( .a(n_37208), .b(n_37115), .o(n_37366) );
no02f80 g776550 ( .a(n_4218), .b(n_3848), .o(n_4341) );
no02f80 g774281 ( .a(n_6696), .b(n_6733), .o(n_6767) );
in01f80 FE_OCPC1471_n_13434 ( .a(n_13434), .o(FE_OCPN1471_n_13434) );
in01f80 g762338 ( .a(n_18834), .o(n_18807) );
no02f80 g746705 ( .a(n_33083), .b(n_32963), .o(n_33386) );
na02f80 g749069 ( .a(n_30933), .b(n_27131), .o(n_30964) );
in01f80 newInst_1028 ( .a(newNet_82), .o(newNet_1028) );
in01f80 g743913 ( .a(n_35954), .o(n_35985) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_14_ ( .ck(newNet_2968), .d(n_5972), .o(delay_add_ln22_unr5_stage3_stallmux_q_14_) );
ao12f80 g741936 ( .a(n_37905), .b(n_37991), .c(n_37867), .o(n_38074) );
no02f80 g750844 ( .a(n_29039), .b(n_28678), .o(n_29095) );
in01f80 g764075 ( .a(n_17093), .o(n_17101) );
in01f80 FE_OCP_RBC2608_n_3807 ( .a(FE_OCP_RBN2607_n_3807), .o(FE_OCP_RBN2608_n_3807) );
na02f80 g778291 ( .a(n_2676), .b(n_2543), .o(n_2763) );
ao12f80 g757077 ( .a(n_23550), .b(n_23549), .c(n_23548), .o(n_24023) );
no02f80 g751439 ( .a(n_28510), .b(n_28494), .o(n_28530) );
na02f80 g747468 ( .a(n_32367), .b(n_44962), .o(n_32578) );
no02f80 g772505 ( .a(n_8456), .b(n_8457), .o(n_8533) );
no02f80 g765820 ( .a(n_14888), .b(n_14864), .o(n_14988) );
in01f80 newInst_2661 ( .a(newNet_1278), .o(newNet_2661) );
no02f80 g749121 ( .a(n_30914), .b(n_27366), .o(n_30996) );
na02f80 g773096 ( .a(n_7646), .b(n_45821), .o(n_7647) );
na02f80 g776070 ( .a(n_5102), .b(n_5078), .o(n_5253) );
in01f80 g759209 ( .a(n_21312), .o(n_21367) );
in01f80 g763691 ( .a(n_16760), .o(n_16761) );
in01f80 newInst_531 ( .a(newNet_530), .o(newNet_531) );
no02f80 g770603 ( .a(n_10267), .b(n_10201), .o(n_10411) );
in01f80 FE_OCP_RBC3725_n_16975 ( .a(FE_OCP_RBN3723_n_16975), .o(FE_OCP_RBN3725_n_16975) );
oa12f80 g767366 ( .a(n_13450), .b(n_13449), .c(n_13448), .o(n_15207) );
in01f80 newInst_2074 ( .a(newNet_1318), .o(newNet_2074) );
na02f80 g770818 ( .a(n_10014), .b(n_9894), .o(n_10091) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_17_ ( .ck(newNet_2869), .d(n_11356), .o(delay_add_ln22_unr8_stage4_stallmux_q_17_) );
in01f80 FE_OCPC1467_n_12968 ( .a(n_12968), .o(FE_OCPN1467_n_12968) );
no02f80 g776962 ( .a(n_3561), .b(n_2797), .o(n_3633) );
ms00f80 mux_while_ln12_psv_q_reg_2_ ( .ck(newNet_121), .d(n_173), .o(mux_while_ln12_psv_q_2_) );
in01f80 g773848 ( .a(n_7129), .o(n_7130) );
in01f80 g751472 ( .a(n_28569), .o(n_28570) );
in01f80 g775864 ( .a(n_5142), .o(n_5143) );
na02f80 g759750 ( .a(n_21775), .b(n_21826), .o(n_21957) );
no02f80 g748246 ( .a(FE_OCP_RBN3083_n_31819), .b(FE_OCPN3793_n_31804), .o(n_31902) );
in01f80 FE_OCP_RBC3382_n_12365 ( .a(n_12365), .o(FE_OCP_RBN3382_n_12365) );
no02f80 FE_RC_1922_0 ( .a(n_29379), .b(n_29091), .o(FE_RN_607_0) );
na02f80 g763811 ( .a(n_17159), .b(n_17158), .o(n_17160) );
no02f80 g759548 ( .a(n_20846), .b(FE_OCPN1444_n_45050), .o(n_20879) );
no02f80 g773077 ( .a(n_8058), .b(n_8012), .o(n_8735) );
no02f80 g772361 ( .a(n_8677), .b(n_8676), .o(n_8714) );
in01f80 g755453 ( .a(n_24659), .o(n_24660) );
no02f80 g755705 ( .a(n_24520), .b(n_24519), .o(n_24521) );
in01f80 g752757 ( .a(n_27957), .o(n_27958) );
in01f80 FE_OCP_RBC2160_n_1675 ( .a(n_1675), .o(FE_OCP_RBN2160_n_1675) );
na02f80 g776167 ( .a(n_47008), .b(FE_OCP_RBN2723_n_4219), .o(n_4660) );
no02f80 g739931 ( .a(n_40336), .b(n_40195), .o(n_40335) );
in01f80 g768025 ( .a(n_12992), .o(n_12993) );
in01f80 g767462 ( .a(n_13232), .o(n_13272) );
na02f80 g739154 ( .a(n_40958), .b(n_40873), .o(n_40959) );
in01f80 g752528 ( .a(n_27693), .o(n_27666) );
no02f80 g756825 ( .a(n_23958), .b(n_23910), .o(n_23959) );
no02f80 g774514 ( .a(n_6585), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_10_), .o(n_6658) );
in01f80 g746141 ( .a(n_33937), .o(n_33938) );
no02f80 g740386 ( .a(n_39803), .b(n_39878), .o(n_39880) );
oa22f80 g744499 ( .a(n_36684), .b(n_36176), .c(n_36683), .d(n_36177), .o(n_36729) );
ao12f80 g760374 ( .a(n_20004), .b(n_20030), .c(n_19979), .o(n_20081) );
in01f80 g740580 ( .a(n_39691), .o(n_39692) );
in01f80 newInst_2194 ( .a(newNet_2193), .o(newNet_2194) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_7_ ( .ck(newNet_2995), .d(n_1018), .o(delay_add_ln22_unr2_stage2_stallmux_q_7_) );
no02f80 g749764 ( .a(n_31322), .b(n_31321), .o(n_31323) );
na02f80 g756943 ( .a(n_24215), .b(n_23904), .o(n_24383) );
no02f80 g744900 ( .a(n_35047), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35093) );
ao12f80 g784689 ( .a(n_3360), .b(n_3340), .c(n_3152), .o(n_47019) );
in01f80 newInst_2766 ( .a(newNet_2765), .o(newNet_2766) );
in01f80 g757205 ( .a(n_23378), .o(n_23113) );
in01f80 newInst_412 ( .a(newNet_131), .o(newNet_412) );
na02f80 g771600 ( .a(n_9239), .b(n_9264), .o(n_9334) );
in01f80 g775960 ( .a(n_5234), .o(n_5235) );
in01f80 newInst_850 ( .a(newNet_849), .o(newNet_850) );
ao12f80 g768513 ( .a(n_12180), .b(n_12341), .c(n_12273), .o(n_12412) );
no02f80 g742383 ( .a(n_37707), .b(n_37709), .o(n_37710) );
no02f80 g750098 ( .a(n_29857), .b(n_28889), .o(n_29986) );
na02f80 g778471 ( .a(n_2570), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .o(n_2666) );
no02f80 g745609 ( .a(n_34369), .b(n_34504), .o(n_34704) );
in01f80 newInst_3293 ( .a(newNet_3292), .o(newNet_3293) );
in01f80 g754073 ( .a(n_26167), .o(n_26196) );
in01f80 g764468 ( .a(n_16423), .o(n_16317) );
no03m80 g748771 ( .a(n_32413), .b(n_32502), .c(n_32441), .o(n_32535) );
na02f80 g755353 ( .a(n_24839), .b(n_24838), .o(n_24860) );
no02f80 g767085 ( .a(n_13718), .b(n_13717), .o(n_13719) );
oa12f80 g779049 ( .a(n_2089), .b(n_2105), .c(n_2088), .o(n_2161) );
no02f80 g780634 ( .a(n_923), .b(n_658), .o(n_929) );
in01f80 g748529 ( .a(n_31466), .o(n_31730) );
in01f80 g755596 ( .a(n_24711), .o(n_24712) );
in01f80 newInst_321 ( .a(newNet_320), .o(newNet_321) );
na02f80 g745369 ( .a(n_36049), .b(n_35391), .o(n_36122) );
oa22f80 g749442 ( .a(n_31939), .b(n_31621), .c(n_31940), .d(n_31622), .o(n_32005) );
in01f80 g749532 ( .a(n_30452), .o(n_30471) );
na02f80 g736515 ( .a(n_43654), .b(n_43235), .o(n_43664) );
ao12f80 g751011 ( .a(n_28529), .b(n_28853), .c(n_28511), .o(n_28871) );
no02f80 g780492 ( .a(n_819), .b(n_884), .o(n_895) );
no02f80 g757794 ( .a(n_22411), .b(n_22555), .o(n_22593) );
in01f80 FE_OCP_RBC1060_n_24473 ( .a(n_24473), .o(FE_OCP_RBN1060_n_24473) );
ao12f80 g745087 ( .a(n_34898), .b(n_34897), .c(n_34896), .o(n_34966) );
na02f80 g764227 ( .a(n_16460), .b(n_16485), .o(n_16582) );
in01f80 fopt783266 ( .a(n_36410), .o(n_44835) );
in01f80 newInst_1391 ( .a(newNet_1390), .o(newNet_1391) );
no02f80 g767496 ( .a(n_13291), .b(n_13290), .o(n_13292) );
in01f80 g758760 ( .a(n_21620), .o(n_21680) );
oa22f80 g748854 ( .a(n_32316), .b(n_31579), .c(n_44764), .d(n_31578), .o(n_32379) );
in01f80 g780972 ( .a(n_420), .o(n_457) );
in01f80 fopt784023 ( .a(n_45760), .o(n_45758) );
no02f80 g761316 ( .a(n_19954), .b(n_19899), .o(n_20053) );
in01f80 newInst_1993 ( .a(newNet_1992), .o(newNet_1993) );
oa12f80 g751704 ( .a(n_28247), .b(n_28303), .c(n_28223), .o(n_28391) );
in01f80 g739952 ( .a(n_40049), .o(n_40087) );
na02f80 g751403 ( .a(n_28580), .b(n_28632), .o(n_28651) );
in01f80 g739811 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n_40499) );
no02f80 g748441 ( .a(n_31474), .b(FE_OCPN1446_n_31473), .o(n_31499) );
in01f80 g779664 ( .a(delay_xor_ln21_unr3_stage2_stallmux_q_0_), .o(n_1362) );
na02f80 g769289 ( .a(n_11456), .b(n_11398), .o(n_11511) );
in01f80 g768766 ( .a(n_12117), .o(n_12113) );
na02f80 g756048 ( .a(n_25139), .b(n_25132), .o(n_25197) );
na02f80 g766569 ( .a(n_13925), .b(n_13424), .o(n_14021) );
in01f80 g772645 ( .a(n_8335), .o(n_8336) );
in01f80 g778266 ( .a(n_3014), .o(n_3015) );
in01f80 g763750 ( .a(n_16706), .o(n_16707) );
na02f80 g777619 ( .a(n_3519), .b(n_3479), .o(n_3542) );
in01f80 g779630 ( .a(n_1764), .o(n_1765) );
in01f80 g754111 ( .a(n_26978), .o(n_26950) );
na02f80 FE_RC_1279_0 ( .a(FE_RN_377_0), .b(n_2915), .o(n_47023) );
in01f80 g780018 ( .a(n_1270), .o(n_1271) );
ao12f80 g771477 ( .a(n_7622), .b(n_8818), .c(n_7633), .o(n_8943) );
no02f80 g740546 ( .a(n_39647), .b(n_39621), .o(n_39690) );
na02f80 g745764 ( .a(n_34115), .b(n_34148), .o(n_34209) );
in01f80 g759837 ( .a(n_22280), .o(n_24620) );
oa12f80 g751208 ( .a(n_28780), .b(n_28791), .c(n_28779), .o(n_28830) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_12_ ( .ck(newNet_2589), .d(n_27279), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_) );
na02f80 g749699 ( .a(n_31431), .b(n_31415), .o(n_31453) );
in01f80 newInst_827 ( .a(newNet_826), .o(newNet_827) );
in01f80 g748659 ( .a(n_31486), .o(n_31487) );
no02f80 g739190 ( .a(n_40857), .b(n_40883), .o(n_40936) );
oa22f80 FE_RC_265_0 ( .a(n_22039), .b(n_21985), .c(n_22038), .d(n_44296), .o(n_22066) );
no02f80 g736438 ( .a(n_43721), .b(n_43444), .o(n_43731) );
in01f80 fopt782793 ( .a(n_32360), .o(n_44213) );
in01f80 FE_RC_1110_0 ( .a(delay_xor_ln22_unr6_stage3_stallmux_q_3_), .o(FE_RN_333_0) );
no02f80 g742797 ( .a(n_37310), .b(n_37147), .o(n_37333) );
ao22s80 g761897 ( .a(n_18704), .b(n_17724), .c(n_18284), .d(delay_sub_ln21_0_unr11_stage5_stallmux_q_31_), .o(n_18912) );
oa12f80 g737854 ( .a(n_42214), .b(FE_OCPN1232_n_42201), .c(n_42212), .o(n_42534) );
in01f80 FE_RC_675_0 ( .a(n_17581), .o(FE_RN_216_0) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_4_ ( .ck(newNet_153), .d(n_46375), .o(delay_xor_ln22_unr9_stage4_stallmux_q_4_) );
no02f80 g757944 ( .a(n_22138), .b(n_22081), .o(n_22139) );
in01f80 g740552 ( .a(FE_OCP_RBN2945_FE_RN_1269_0), .o(n_39665) );
no02f80 g778385 ( .a(n_2430), .b(n_2442), .o(n_2443) );
oa12f80 g736351 ( .a(n_298), .b(n_43838), .c(FE_OFN1_n_43918), .o(n_43869) );
oa12f80 g752711 ( .a(n_28054), .b(n_27954), .c(n_27923), .o(n_28615) );
in01f80 newInst_2569 ( .a(newNet_2568), .o(newNet_2569) );
na02f80 g773899 ( .a(n_7050), .b(n_5438), .o(n_7107) );
in01f80 FE_OCP_RBC1692_n_19052 ( .a(FE_OCPN1738_n_19052), .o(FE_OCP_RBN1692_n_19052) );
na02f80 g744219 ( .a(n_36096), .b(n_36089), .o(n_36236) );
no02f80 g748934 ( .a(n_31136), .b(n_31108), .o(n_31156) );
in01f80 newInst_1522 ( .a(newNet_1521), .o(newNet_1522) );
oa12f80 g746877 ( .a(n_34105), .b(n_34104), .c(n_34103), .o(n_34667) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_11_ ( .ck(newNet_3566), .d(n_21967), .o(delay_add_ln22_unr14_stage6_stallmux_q_11_) );
in01f80 g776956 ( .a(n_3968), .o(n_3969) );
in01f80 FE_RC_4052_0 ( .a(n_14768), .o(FE_RN_1762_0) );
na02f80 g753124 ( .a(n_27463), .b(n_27462), .o(n_27502) );
na02f80 g769333 ( .a(FE_OCP_RBN2002_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_2_), .o(n_11548) );
in01f80 newInst_150 ( .a(newNet_20), .o(newNet_150) );
na02f80 FE_RC_2373_0 ( .a(FE_RN_921_0), .b(n_42285), .o(FE_RN_922_0) );
in01f80 FE_OFC734_n_22641 ( .a(n_22641), .o(FE_OFN734_n_22641) );
in01f80 g746335 ( .a(n_33673), .o(n_33708) );
in01f80 FE_OCP_RBC3112_n_32254 ( .a(n_32254), .o(FE_OCP_RBN3112_n_32254) );
no02f80 g771081 ( .a(n_9907), .b(n_9906), .o(n_9959) );
na02f80 g777733 ( .a(n_3426), .b(n_3488), .o(n_3509) );
in01f80 g740675 ( .a(FE_OCP_RBN2871_n_39542), .o(n_39555) );
ao22s80 g780997 ( .a(n_284), .b(n_139), .c(n_281), .d(n_138), .o(n_495) );
in01f80 g772329 ( .a(n_8806), .o(n_8807) );
in01f80 newInst_287 ( .a(newNet_286), .o(newNet_287) );
in01f80 g755948 ( .a(n_24254), .o(n_24267) );
na02f80 g767751 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_24_), .o(n_13238) );
oa12f80 g760292 ( .a(n_20106), .b(n_20081), .c(n_19967), .o(n_20174) );
oa22f80 FE_RC_1486_0 ( .a(n_27630), .b(n_27267), .c(n_27268), .d(n_27631), .o(n_27727) );
in01f80 FE_OCP_RBC3625_n_38870 ( .a(FE_OCP_RBN2685_n_38870), .o(FE_OCP_RBN3625_n_38870) );
no02f80 g746834 ( .a(n_33449), .b(n_33102), .o(n_33482) );
na02f80 g762114 ( .a(n_18702), .b(n_18500), .o(n_18847) );
na02f80 g775795 ( .a(n_5070), .b(n_5097), .o(n_5255) );
ms00f80 delay_sub_ln23_0_unr27_stage10_stallmux_q_reg ( .ck(newNet_1444), .d(delay_sub_ln23_0_unr27_stage10_stallmux_z), .o(n_44610) );
in01f80 g769797 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_14_), .o(n_12468) );
oa12f80 g741556 ( .a(n_38687), .b(n_38686), .c(n_38685), .o(n_39675) );
in01f80 g755650 ( .a(n_24436), .o(n_24450) );
na02f80 g741039 ( .a(n_39245), .b(n_39304), .o(n_39331) );
na02f80 g773917 ( .a(n_7017), .b(n_7016), .o(n_7208) );
oa22f80 g744857 ( .a(n_36405), .b(n_36157), .c(n_36406), .d(n_36158), .o(n_36454) );
in01f80 FE_OCP_RBC3429_n_13245 ( .a(n_13245), .o(FE_OCP_RBN3429_n_13245) );
in01f80 g762825 ( .a(n_17822), .o(n_17823) );
na02f80 g739379 ( .a(n_40807), .b(n_40873), .o(n_41130) );
in01f80 newInst_3388 ( .a(newNet_3387), .o(newNet_3388) );
no02f80 g740252 ( .a(n_39934), .b(n_39969), .o(n_39970) );
in01f80 g738251 ( .a(n_41982), .o(n_41992) );
ao12f80 g744200 ( .a(n_35265), .b(n_35532), .c(FE_OCP_RBN2809_n_35285), .o(n_35550) );
ao12f80 g763859 ( .a(n_17297), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n_17602) );
no02f80 FE_RC_3960_0 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .b(n_23599), .o(FE_RN_1715_0) );
in01f80 g764208 ( .a(n_16885), .o(n_16886) );
ao12f80 g762986 ( .a(n_17391), .b(n_17350), .c(n_17331), .o(n_17495) );
in01f80 newInst_2720 ( .a(newNet_2719), .o(newNet_2720) );
no02f80 g775132 ( .a(n_5943), .b(n_5964), .o(n_5997) );
no02f80 g748896 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_13_), .o(n_32443) );
in01f80 g749428 ( .a(n_30541), .o(n_31864) );
no02f80 g751186 ( .a(n_29837), .b(n_29312), .o(n_29878) );
na02f80 g748562 ( .a(n_31365), .b(n_31384), .o(n_31474) );
na02f80 g741786 ( .a(n_38510), .b(n_38483), .o(n_38511) );
in01f80 FE_OCP_RBC3455_FE_OCPN1240_n_7721 ( .a(FE_OCP_RBN3454_FE_OCPN1240_n_7721), .o(FE_OCP_RBN3455_FE_OCPN1240_n_7721) );
na02f80 g753287 ( .a(FE_OCPN964_n_27287), .b(n_26653), .o(n_27327) );
oa22f80 g743716 ( .a(n_36277), .b(n_35638), .c(n_36247), .d(n_35639), .o(n_36345) );
na02f80 g751898 ( .a(n_28897), .b(n_29041), .o(n_29070) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_4_ ( .ck(newNet_2908), .d(n_4828), .o(delay_add_ln22_unr5_stage3_stallmux_q_4_) );
in01f80 g763522 ( .a(n_16902), .o(n_16942) );
na02f80 g764928 ( .a(n_15679), .b(n_15678), .o(n_15723) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_16_ ( .ck(newNet_2964), .d(n_6063), .o(delay_add_ln22_unr5_stage3_stallmux_q_16_) );
in01f80 FE_RC_3851_0 ( .a(FE_RN_1681_0), .o(n_19724) );
no02f80 g777842 ( .a(n_3198), .b(n_2426), .o(n_3230) );
no02f80 g737710 ( .a(n_42394), .b(n_42172), .o(n_42469) );
na02f80 g755442 ( .a(n_24750), .b(n_24691), .o(n_24783) );
in01f80 g771447 ( .a(n_9404), .o(n_9405) );
oa12f80 g759813 ( .a(n_21335), .b(n_21714), .c(n_21244), .o(n_22057) );
no02f80 g761005 ( .a(n_19274), .b(n_18851), .o(n_19327) );
no02f80 g736635 ( .a(n_43441), .b(n_43371), .o(n_43481) );
no02f80 g751628 ( .a(n_28405), .b(delay_add_ln22_unr17_stage7_stallmux_q_12_), .o(n_28423) );
in01f80 g777955 ( .a(n_4662), .o(n_3118) );
na02f80 g776932 ( .a(n_4023), .b(n_4022), .o(n_4175) );
no02f80 FE_RC_2889_0 ( .a(FE_OCPN1858_n_22207), .b(n_24684), .o(FE_RN_1251_0) );
oa22f80 g736908 ( .a(n_43230), .b(FE_OCP_RBN2915_n_42947), .c(FE_OCP_RBN3074_n_43230), .d(n_42961), .o(n_43634) );
na02f80 g748326 ( .a(n_31755), .b(n_31799), .o(n_31838) );
in01f80 FE_OCP_RBC1197_n_30619 ( .a(n_30619), .o(FE_OCP_RBN1197_n_30619) );
ao12f80 g750259 ( .a(n_29737), .b(n_29736), .c(n_29602), .o(n_29738) );
na02f80 g761470 ( .a(n_19980), .b(n_19794), .o(n_20196) );
in01f80 newInst_1306 ( .a(newNet_1305), .o(newNet_1306) );
in01f80 g748591 ( .a(n_32674), .o(n_32675) );
in01f80 FE_OCPC961_n_28506 ( .a(n_28506), .o(FE_OCPN961_n_28506) );
in01f80 g755779 ( .a(n_25371), .o(n_25342) );
na02f80 FE_RC_1780_0 ( .a(FE_RN_518_0), .b(n_2240), .o(FE_RN_519_0) );
in01f80 g771462 ( .a(n_9290), .o(n_9291) );
in01f80 g768049 ( .a(n_12882), .o(n_12883) );
na02f80 g736554 ( .a(n_43638), .b(n_43286), .o(n_43661) );
oa22f80 g745334 ( .a(n_36049), .b(n_35842), .c(FE_OCP_RBN2995_n_35539), .d(n_35476), .o(n_36213) );
in01f80 FE_OCP_RBC2950_n_21363 ( .a(n_21363), .o(FE_OCP_RBN2950_n_21363) );
no02f80 g776670 ( .a(n_4053), .b(n_4077), .o(n_4283) );
no02f80 g762837 ( .a(n_17598), .b(n_17036), .o(n_17657) );
na02f80 g779343 ( .a(n_1608), .b(n_1633), .o(n_1634) );
na02f80 g744283 ( .a(FE_OCPN1510_n_44174), .b(n_35025), .o(n_36090) );
in01f80 newInst_1532 ( .a(newNet_540), .o(newNet_1532) );
no02f80 g762015 ( .a(n_18309), .b(n_18337), .o(n_18357) );
na02f80 g743920 ( .a(n_36099), .b(n_36037), .o(n_36270) );
oa12f80 g738324 ( .a(n_41475), .b(n_41596), .c(n_41426), .o(n_41648) );
na02f80 g738486 ( .a(n_41582), .b(n_41590), .o(n_41680) );
in01f80 newInst_1192 ( .a(newNet_1191), .o(newNet_1192) );
no02f80 g742206 ( .a(n_44887), .b(n_37884), .o(n_38296) );
ao12f80 g750892 ( .a(n_30156), .b(n_30183), .c(n_29852), .o(n_30235) );
na02f80 g764491 ( .a(FE_OCP_RBN3686_n_16074), .b(n_14618), .o(n_16224) );
ao12f80 g743713 ( .a(n_37361), .b(n_37405), .c(n_46235), .o(n_37472) );
oa12f80 g780155 ( .a(n_1123), .b(n_1139), .c(n_1122), .o(n_1164) );
in01f80 newInst_2084 ( .a(newNet_2083), .o(newNet_2084) );
in01f80 newInst_1137 ( .a(newNet_1136), .o(newNet_1137) );
in01f80 g761846 ( .a(n_18551), .o(n_19893) );
na02f80 g772935 ( .a(n_8009), .b(n_7850), .o(n_8010) );
no02f80 g745850 ( .a(n_34138), .b(n_34137), .o(n_34157) );
in01f80 fopt782677 ( .a(n_44066), .o(n_44071) );
no02f80 g760726 ( .a(n_19588), .b(FE_OCPN1426_n_18099), .o(n_19698) );
ao12f80 g765231 ( .a(n_15874), .b(n_15969), .c(n_15512), .o(n_15970) );
in01f80 g757033 ( .a(n_23986), .o(n_23934) );
na02f80 g780091 ( .a(n_1184), .b(n_1171), .o(n_1172) );
no02f80 g737772 ( .a(n_42227), .b(n_42226), .o(n_42537) );
ao22s80 g760850 ( .a(n_19387), .b(FE_OCP_RBN1351_n_19148), .c(n_19386), .d(n_19164), .o(n_19563) );
na02f80 g739230 ( .a(n_40887), .b(n_40886), .o(n_41260) );
in01f80 g758186 ( .a(n_22194), .o(n_22214) );
na02f80 g751971 ( .a(n_28897), .b(n_28939), .o(n_29025) );
na02f80 g742553 ( .a(FE_OCP_RBN2174_n_37559), .b(n_37557), .o(n_37558) );
in01f80 g760820 ( .a(n_19537), .o(n_19558) );
in01f80 g743500 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_28_), .o(n_36625) );
in01f80 newInst_18 ( .a(newNet_9), .o(newNet_18) );
ao12f80 g751399 ( .a(n_29227), .b(n_29226), .c(n_29225), .o(n_29311) );
na02f80 g771693 ( .a(n_9126), .b(n_8269), .o(n_9355) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_4_ ( .ck(newNet_493), .d(n_22716), .o(delay_xor_ln22_unr15_stage6_stallmux_q_4_) );
in01f80 g754501 ( .a(n_25601), .o(n_25567) );
oa12f80 g755317 ( .a(n_25578), .b(n_25577), .c(n_25576), .o(n_26310) );
na02f80 g773904 ( .a(n_7021), .b(delay_add_ln22_unr5_stage3_stallmux_q_8_), .o(n_7086) );
in01f80 fopt783250 ( .a(FE_OCP_RBN3411_n_33547), .o(n_44814) );
in01f80 g774742 ( .a(n_6350), .o(n_6351) );
no02f80 g742058 ( .a(FE_OCP_RBN2257_n_37844), .b(n_37385), .o(n_38016) );
ao12f80 g741846 ( .a(n_38361), .b(n_38360), .c(n_38359), .o(n_38469) );
oa12f80 g750448 ( .a(n_30000), .b(n_30552), .c(n_30381), .o(n_30590) );
in01f80 g766910 ( .a(n_13575), .o(n_13576) );
in01f80 FE_OCPC931_n_40736 ( .a(n_40736), .o(FE_OCPN931_n_40736) );
na02f80 g773903 ( .a(n_7051), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .o(n_7106) );
in01f80 FE_OCP_RBC3854_n_20848 ( .a(FE_OCP_RBN3853_n_20848), .o(FE_OCP_RBN3854_n_20848) );
in01f80 g780586 ( .a(n_675), .o(n_667) );
no02f80 g776308 ( .a(n_4704), .b(n_4274), .o(n_4830) );
in01f80 FE_OCPC1417_n_31504 ( .a(n_31504), .o(FE_OCPN1417_n_31504) );
na02f80 g749483 ( .a(n_30452), .b(n_30240), .o(n_30455) );
na02f80 g743895 ( .a(n_35710), .b(n_35709), .o(n_35711) );
ao22s80 g768000 ( .a(n_12646), .b(n_12429), .c(n_12645), .d(n_12430), .o(n_12905) );
in01f80 newInst_1148 ( .a(newNet_706), .o(newNet_1148) );
in01f80 g746318 ( .a(n_33589), .o(n_33774) );
na02f80 g774795 ( .a(n_6214), .b(n_5523), .o(n_6265) );
oa12f80 g761835 ( .a(n_18126), .b(n_18318), .c(n_18127), .o(n_18376) );
no02f80 g755334 ( .a(n_24879), .b(n_24878), .o(n_24880) );
no02f80 g741703 ( .a(n_38535), .b(n_38200), .o(n_38577) );
na02f80 g748422 ( .a(n_31730), .b(n_30871), .o(n_31725) );
ao12f80 g762980 ( .a(n_17543), .b(n_17939), .c(n_17301), .o(n_17990) );
ao12f80 g745467 ( .a(n_35510), .b(n_35509), .c(n_35508), .o(n_36019) );
na02f80 g767416 ( .a(n_13367), .b(FE_OCPN1854_n_13366), .o(n_13383) );
oa22f80 g780858 ( .a(n_420), .b(n_376), .c(n_457), .d(n_384), .o(n_564) );
oa22f80 g746410 ( .a(n_33429), .b(n_33304), .c(n_33331), .d(n_33303), .o(n_34296) );
in01f80 g778071 ( .a(n_3000), .o(n_2996) );
no02f80 g765942 ( .a(n_14697), .b(n_14698), .o(n_14773) );
oa22f80 FE_RC_1419_0 ( .a(FE_OFN806_n_46196), .b(n_6643), .c(FE_OFN84_n_46137), .d(n_6587), .o(n_46189) );
no02f80 FE_RC_1843_0 ( .a(n_44223), .b(FE_RN_558_0), .o(FE_RN_559_0) );
in01f80 g753445 ( .a(n_27006), .o(n_27007) );
no02f80 g762378 ( .a(FE_OCP_RBN3410_n_45120), .b(n_18492), .o(n_18528) );
na02f80 g741984 ( .a(n_38216), .b(n_38217), .o(n_38218) );
in01f80 g773031 ( .a(n_7686), .o(n_7687) );
na02f80 g778628 ( .a(n_2745), .b(n_2744), .o(n_2746) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_23_ ( .ck(newNet_814), .d(n_1317), .o(delay_xor_ln21_unr3_stage2_stallmux_q_23_) );
in01f80 g755054 ( .a(n_25585), .o(n_25586) );
in01f80 FE_OCP_RBC3116_n_22710 ( .a(n_22710), .o(FE_OCP_RBN3116_n_22710) );
in01f80 FE_OCP_RBC2857_n_10399 ( .a(n_10399), .o(FE_OCP_RBN2857_n_10399) );
na02f80 g753713 ( .a(n_26442), .b(FE_RN_1667_0), .o(n_26504) );
in01f80 g762388 ( .a(n_18658), .o(n_18610) );
na02f80 g767702 ( .a(n_13314), .b(n_13236), .o(n_13797) );
in01f80 newInst_3705 ( .a(newNet_3704), .o(newNet_3705) );
in01f80 g745101 ( .a(n_34753), .o(n_34754) );
oa12f80 g776609 ( .a(n_4402), .b(n_4401), .c(n_4400), .o(n_4491) );
na02f80 g776211 ( .a(n_4734), .b(n_4629), .o(n_4906) );
in01f80 g748304 ( .a(n_31895), .o(n_31896) );
oa12f80 g780116 ( .a(n_1086), .b(n_1085), .c(n_1084), .o(n_1135) );
in01f80 FE_OCP_RBC3548_n_44575 ( .a(FE_OCP_RBN3543_n_44575), .o(FE_OCP_RBN3548_n_44575) );
no02f80 g759164 ( .a(n_21013), .b(n_20977), .o(n_21082) );
in01f80 fopt783286 ( .a(n_5048), .o(n_44862) );
na02f80 g757980 ( .a(n_22083), .b(n_22046), .o(n_22138) );
in01f80 g747253 ( .a(n_32786), .o(n_32787) );
na02f80 g770616 ( .a(n_10379), .b(FE_OCP_RBN3558_n_8687), .o(n_10393) );
in01f80 g768657 ( .a(n_12294), .o(n_12227) );
no02f80 g740138 ( .a(n_39781), .b(n_39800), .o(n_39801) );
oa12f80 g751622 ( .a(FE_OCP_RBN2216_FE_OCPN950_n_28595), .b(n_28795), .c(n_27778), .o(n_28798) );
no02f80 g741120 ( .a(n_38994), .b(n_38993), .o(n_39285) );
no02f80 g764952 ( .a(FE_OCP_RBN2743_n_15319), .b(FE_OCPN1007_n_13962), .o(n_15393) );
no02f80 g784699 ( .a(n_20250), .b(n_20229), .o(n_47175) );
no02f80 g772805 ( .a(n_8041), .b(n_7782), .o(n_8097) );
in01f80 g743854 ( .a(n_37166), .o(n_37167) );
no02f80 g748017 ( .a(n_31974), .b(n_31852), .o(n_31997) );
in01f80 newInst_2096 ( .a(newNet_384), .o(newNet_2096) );
in01f80 g736804 ( .a(n_43516), .o(n_43517) );
in01f80 g773211 ( .a(n_7759), .o(n_7760) );
ao12f80 g746174 ( .a(n_34037), .b(n_33752), .c(n_33728), .o(n_33849) );
na02f80 g755060 ( .a(n_25499), .b(n_25531), .o(n_25552) );
na02f80 g747082 ( .a(n_32930), .b(n_32732), .o(n_33015) );
na02f80 g777398 ( .a(n_3521), .b(n_2759), .o(n_3551) );
in01f80 FE_OCPC1468_n_12968 ( .a(FE_OCPN1467_n_12968), .o(FE_OCPN1468_n_12968) );
no02f80 g750922 ( .a(n_29012), .b(n_29011), .o(n_29013) );
na02f80 g781015 ( .a(cos_out_1), .b(FE_OFN5_n_43918), .o(n_321) );
oa12f80 g780077 ( .a(n_841), .b(n_1199), .c(n_793), .o(n_1215) );
na02f80 g737032 ( .a(n_43082), .b(n_43121), .o(n_43084) );
in01f80 FE_OCP_RBC3636_n_47260 ( .a(FE_OCP_RBN3635_n_47260), .o(FE_OCP_RBN3636_n_47260) );
in01f80 g771995 ( .a(n_10081), .o(n_10036) );
in01f80 g744042 ( .a(n_35699), .o(n_35744) );
no03m80 g738175 ( .a(n_41600), .b(n_42007), .c(n_41614), .o(n_42079) );
no02f80 g762091 ( .a(n_18355), .b(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n_18589) );
in01f80 FE_OCP_DRV_C1560_n_34288 ( .a(FE_OCP_DRV_N1559_n_34288), .o(FE_OCP_DRV_N1560_n_34288) );
in01f80 FE_RC_2614_0 ( .a(n_14558), .o(FE_RN_1088_0) );
in01f80 g766239 ( .a(n_14444), .o(n_14464) );
oa22f80 FE_RC_1158_0 ( .a(n_11806), .b(n_12027), .c(n_11807), .d(FE_OCP_RBN3737_n_12027), .o(n_12240) );
in01f80 g747515 ( .a(n_33721), .o(n_34211) );
in01f80 g744753 ( .a(n_35303), .o(n_35304) );
no02f80 g778735 ( .a(n_2438), .b(n_2596), .o(n_2612) );
no02f80 FE_RC_2263_0 ( .a(FE_RN_838_0), .b(FE_RN_837_0), .o(FE_RN_839_0) );
in01f80 g775045 ( .a(n_6169), .o(n_6170) );
in01f80 FE_RC_2271_0 ( .a(n_33680), .o(FE_RN_845_0) );
na02f80 g763382 ( .a(FE_OCP_RBN3725_n_16975), .b(n_15762), .o(n_17328) );
in01f80 g745968 ( .a(n_33966), .o(n_33967) );
no02f80 g738206 ( .a(n_41972), .b(n_41803), .o(n_42009) );
no02f80 g752724 ( .a(n_27883), .b(n_27988), .o(n_27933) );
oa22f80 FE_RC_4264_0 ( .a(n_32730), .b(n_32815), .c(n_32729), .d(n_32816), .o(n_32906) );
in01f80 g751083 ( .a(n_29852), .o(n_30207) );
na02f80 g779403 ( .a(n_1509), .b(n_1486), .o(n_1525) );
ao12f80 g779413 ( .a(n_1502), .b(n_1501), .c(n_1515), .o(n_1565) );
ao12f80 g763422 ( .a(FE_OCP_RBN3360_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .b(n_17577), .c(n_17496), .o(n_17578) );
no02f80 g755601 ( .a(n_24473), .b(n_24344), .o(n_24474) );
na02f80 g766834 ( .a(n_13658), .b(n_13705), .o(n_13748) );
no02f80 g781326 ( .a(n_1), .b(beta_4), .o(n_78) );
in01f80 g744728 ( .a(n_35235), .o(n_35183) );
na02f80 g757015 ( .a(n_24188), .b(n_23978), .o(n_24215) );
in01f80 FE_OCP_RBC2541_n_8800 ( .a(n_8800), .o(FE_OCP_RBN2541_n_8800) );
in01f80 newInst_3130 ( .a(newNet_3129), .o(newNet_3130) );
na02f80 g738830 ( .a(n_41311), .b(n_41319), .o(n_41341) );
ao12f80 g746751 ( .a(n_32743), .b(n_32924), .c(n_32775), .o(n_32980) );
na02f80 g751415 ( .a(n_29255), .b(n_29254), .o(n_29256) );
no02f80 g774804 ( .a(n_6244), .b(n_6240), .o(n_6334) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_7_ ( .ck(newNet_773), .d(n_1324), .o(delay_xor_ln21_unr3_stage2_stallmux_q_7_) );
in01f80 FE_OCP_RBC2562_n_34905 ( .a(n_34905), .o(FE_OCP_RBN2562_n_34905) );
oa12f80 g749888 ( .a(n_29807), .b(n_29816), .c(n_29775), .o(n_29875) );
no02f80 g778594 ( .a(n_2449), .b(n_2448), .o(n_2985) );
oa12f80 g768480 ( .a(n_12411), .b(n_12360), .c(FE_OCPN1002_n_45660), .o(n_12606) );
in01f80 g754130 ( .a(n_26176), .o(n_26139) );
no02f80 g761039 ( .a(n_19208), .b(n_19181), .o(n_19271) );
na02f80 g741622 ( .a(n_38596), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38626) );
in01f80 newInst_1365 ( .a(newNet_1364), .o(newNet_1365) );
oa12f80 g738381 ( .a(n_41432), .b(n_41431), .c(n_41430), .o(n_41515) );
in01f80 g750367 ( .a(n_30662), .o(n_30687) );
na02f80 g766816 ( .a(n_13943), .b(n_13941), .o(n_13942) );
na02f80 g738166 ( .a(n_42003), .b(n_42001), .o(n_42002) );
na02f80 g739983 ( .a(n_39849), .b(n_39795), .o(n_39929) );
na02f80 g754545 ( .a(n_26638), .b(n_26710), .o(n_26738) );
in01f80 g773394 ( .a(n_7588), .o(n_7589) );
in01f80 g772264 ( .a(n_8709), .o(n_8710) );
oa12f80 g745202 ( .a(n_34290), .b(n_34573), .c(n_34353), .o(n_34594) );
in01f80 g742215 ( .a(n_38271), .o(n_38272) );
in01f80 g737917 ( .a(n_42558), .o(n_42559) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_18_ ( .ck(newNet_2660), .d(n_46965), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_) );
oa22f80 FE_RC_2896_0 ( .a(FE_OCP_RBN2898_n_45484), .b(n_5315), .c(n_45484), .d(n_5316), .o(n_5454) );
in01f80 newInst_2839 ( .a(newNet_2266), .o(newNet_2839) );
na02f80 g741253 ( .a(FE_OCP_RBN2636_n_38806), .b(n_38563), .o(n_39007) );
in01f80 g754304 ( .a(n_25900), .o(n_25901) );
no02f80 g756282 ( .a(n_24117), .b(n_24119), .o(n_24389) );
na02f80 g757187 ( .a(n_23209), .b(n_23190), .o(n_23366) );
in01f80 FE_OCPC1864_n_26171 ( .a(FE_OCPN1863_n_26171), .o(FE_OCPN1864_n_26171) );
in01f80 newInst_334 ( .a(newNet_240), .o(newNet_334) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_13_ ( .ck(newNet_588), .d(n_17755), .o(delay_xor_ln22_unr12_stage5_stallmux_q_13_) );
no02f80 g745580 ( .a(n_34297), .b(n_34294), .o(n_34357) );
no02f80 g748252 ( .a(n_30499), .b(n_31835), .o(n_31869) );
in01f80 g749896 ( .a(n_31249), .o(n_31374) );
in01f80 newInst_1114 ( .a(newNet_1113), .o(newNet_1114) );
na02f80 g755874 ( .a(n_24955), .b(n_24930), .o(n_25060) );
in01f80 g750088 ( .a(n_29894), .o(n_29895) );
no02f80 g739424 ( .a(n_44769), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_), .o(n_40806) );
na02f80 g744035 ( .a(n_44223), .b(n_34707), .o(n_36298) );
in01f80 FE_OCP_RBC1921_n_22476 ( .a(FE_OCP_RBN1920_n_22476), .o(FE_OCP_RBN1921_n_22476) );
no02f80 g745093 ( .a(n_34824), .b(n_34823), .o(n_34825) );
in01f80 FE_OCP_RBC3206_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3206_n_44365) );
na02f80 g756639 ( .a(n_23626), .b(n_23635), .o(n_23651) );
na02f80 g760507 ( .a(n_19976), .b(n_19975), .o(n_19977) );
in01f80 g774120 ( .a(n_7198), .o(n_7199) );
na02f80 g770555 ( .a(n_10287), .b(n_10398), .o(n_10433) );
in01f80 g746504 ( .a(n_33223), .o(n_33224) );
in01f80 g768620 ( .a(n_12211), .o(n_12151) );
no02f80 g781123 ( .a(n_236), .b(n_264), .o(n_243) );
in01f80 g742596 ( .a(n_37716), .o(n_37529) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_9_ ( .ck(newNet_603), .d(n_46386), .o(delay_xor_ln21_unr9_stage4_stallmux_q_9_) );
in01f80 newInst_2362 ( .a(newNet_697), .o(newNet_2362) );
no02f80 g765844 ( .a(n_14853), .b(n_14854), .o(n_14924) );
oa22f80 g784542 ( .a(n_11731), .b(FE_OFN802_n_46285), .c(n_11682), .d(FE_OCP_RBN3043_n_46337), .o(n_46363) );
in01f80 g740104 ( .a(n_40283), .o(n_40284) );
in01f80 FE_OCP_RBC2830_n_10198 ( .a(n_10198), .o(FE_OCP_RBN2830_n_10198) );
no02f80 g755390 ( .a(n_24659), .b(n_24704), .o(n_24705) );
in01f80 newInst_1863 ( .a(newNet_1862), .o(newNet_1863) );
no02f80 g759288 ( .a(n_44158), .b(n_21030), .o(n_21181) );
in01f80 g774376 ( .a(n_6962), .o(n_6963) );
no02f80 FE_RC_1949_0 ( .a(FE_OCP_RBN2596_n_25181), .b(FE_RN_624_0), .o(FE_RN_625_0) );
in01f80 newInst_1338 ( .a(newNet_48), .o(newNet_1338) );
in01f80 g780483 ( .a(FE_OFN759_n_45813), .o(n_1203) );
in01f80 g763448 ( .a(n_17319), .o(n_17320) );
no02f80 g771785 ( .a(n_8905), .b(n_8936), .o(n_8966) );
na02f80 g739740 ( .a(n_40538), .b(n_40248), .o(n_40539) );
oa22f80 g779887 ( .a(n_44652), .b(n_1065), .c(n_44623), .d(n_1049), .o(n_1304) );
no02f80 g749133 ( .a(n_30958), .b(n_27315), .o(n_31025) );
in01f80 g775754 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_8_), .o(n_5438) );
in01f80 g774564 ( .a(n_6524), .o(n_6521) );
ao12f80 g756889 ( .a(n_23803), .b(n_23899), .c(n_24023), .o(n_23984) );
na02f80 g746165 ( .a(FE_OCP_RBN2234_n_33648), .b(n_33197), .o(n_33676) );
no02f80 g748764 ( .a(n_31328), .b(n_31327), .o(n_31356) );
in01f80 FE_RC_3622_0 ( .a(FE_RN_1585_0), .o(FE_RN_1586_0) );
in01f80 FE_OCP_RBC3490_n_3390 ( .a(FE_OCP_RBN3488_n_3390), .o(FE_OCP_RBN3490_n_3390) );
na02f80 g769880 ( .a(n_47199), .b(n_11076), .o(n_11187) );
na02f80 g738678 ( .a(FE_OCPN1013_n_41478), .b(n_41605), .o(n_41759) );
in01f80 newInst_637 ( .a(newNet_636), .o(newNet_637) );
in01f80 newInst_1432 ( .a(newNet_1431), .o(newNet_1432) );
in01f80 g743754 ( .a(n_37328), .o(n_37329) );
in01f80 FE_OCP_RBC2784_n_9859 ( .a(n_9859), .o(FE_OCP_RBN2784_n_9859) );
in01f80 newInst_245 ( .a(newNet_244), .o(newNet_245) );
in01f80 g763348 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_), .o(n_17186) );
in01f80 FE_OCPC1447_n_27463 ( .a(n_27463), .o(FE_OCPN1447_n_27463) );
na02f80 g779257 ( .a(n_1815), .b(n_1814), .o(n_1949) );
no02f80 g756265 ( .a(n_24069), .b(n_23681), .o(n_24096) );
in01f80 newInst_855 ( .a(newNet_387), .o(newNet_855) );
in01f80 newInst_1205 ( .a(newNet_1204), .o(newNet_1205) );
ao12f80 g745780 ( .a(n_34845), .b(n_35408), .c(n_34775), .o(n_35435) );
no02f80 g762099 ( .a(n_18208), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_16_), .o(n_18311) );
na02f80 g765320 ( .a(FE_OCP_RBN3514_n_13960), .b(FE_OCP_RBN3619_n_15135), .o(n_15230) );
in01f80 g756914 ( .a(n_23361), .o(n_23393) );
no02f80 g767527 ( .a(n_13096), .b(n_13095), .o(n_13227) );
no02f80 g765577 ( .a(n_15171), .b(n_15133), .o(n_15332) );
in01f80 g738792 ( .a(n_41716), .o(n_41713) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_15_ ( .ck(newNet_1131), .d(n_10744), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_) );
in01f80 g762036 ( .a(n_18323), .o(n_18324) );
in01f80 g767452 ( .a(n_13334), .o(n_13301) );
in01f80 g761506 ( .a(n_18945), .o(n_18978) );
na02f80 g763530 ( .a(FE_OCP_RBN1210_n_16814), .b(n_16089), .o(n_16941) );
na02f80 g744600 ( .a(n_35275), .b(n_35238), .o(n_35276) );
in01f80 g762827 ( .a(n_17907), .o(n_17908) );
na02f80 g765140 ( .a(n_15836), .b(n_15830), .o(n_15883) );
no02f80 g761228 ( .a(n_19013), .b(n_18990), .o(n_19077) );
in01f80 fopt783489 ( .a(n_45066), .o(n_45069) );
na02f80 g742736 ( .a(n_37302), .b(n_37301), .o(n_37303) );
ao12f80 g737628 ( .a(n_42566), .b(n_42392), .c(n_42286), .o(n_42661) );
in01f80 g761618 ( .a(n_19649), .o(n_19647) );
in01f80 g777337 ( .a(n_4216), .o(n_4217) );
na02f80 g777134 ( .a(n_4779), .b(n_4796), .o(n_4871) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_11_ ( .ck(newNet_3345), .d(n_31750), .o(delay_add_ln22_unr20_stage8_stallmux_q_11_) );
ao12f80 g756728 ( .a(n_23499), .b(n_23514), .c(n_23498), .o(n_24943) );
ao12f80 g758026 ( .a(n_21910), .b(n_21999), .c(n_21947), .o(n_22080) );
na02f80 g772855 ( .a(n_46991), .b(n_7730), .o(n_8029) );
no02f80 g767773 ( .a(n_13025), .b(n_13024), .o(n_13083) );
no02f80 g779731 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .o(n_1748) );
no02f80 FE_RC_2665_0 ( .a(n_2258), .b(FE_RN_1113_0), .o(n_2508) );
na02f80 g760250 ( .a(FE_OCP_RBN1332_n_20249), .b(n_19236), .o(n_20302) );
no02f80 g763787 ( .a(n_16683), .b(FE_OCP_RBN3060_FE_RN_640_0), .o(n_16749) );
no02f80 g750595 ( .a(n_29329), .b(FE_OCP_RBN2215_FE_OCPN950_n_28595), .o(n_29354) );
na02f80 g744885 ( .a(n_34933), .b(n_30588), .o(n_34985) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_9_ ( .ck(newNet_1783), .d(n_16549), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_9_) );
na02f80 g751579 ( .a(n_28447), .b(n_27637), .o(n_28549) );
no02f80 g745657 ( .a(n_35432), .b(n_34885), .o(n_35461) );
in01f80 g742621 ( .a(n_37587), .o(n_37588) );
in01f80 newInst_466 ( .a(newNet_465), .o(newNet_466) );
no02f80 g775915 ( .a(n_4959), .b(FE_OCPN846_n_4046), .o(n_5200) );
na02f80 g736590 ( .a(n_43447), .b(n_43495), .o(n_43627) );
na02f80 g750390 ( .a(n_29634), .b(n_29612), .o(n_29635) );
no02f80 g736767 ( .a(n_43271), .b(n_43147), .o(n_43148) );
ao12f80 g751069 ( .a(n_29975), .b(n_30303), .c(n_29534), .o(n_30548) );
oa12f80 g736398 ( .a(n_327), .b(n_43758), .c(FE_OFN3_n_43918), .o(n_43803) );
na02f80 g772027 ( .a(n_8950), .b(n_47243), .o(n_9030) );
na02f80 g752144 ( .a(n_28638), .b(n_28637), .o(n_28639) );
no02f80 g755449 ( .a(n_24826), .b(n_24825), .o(n_24892) );
in01f80 FE_RC_2561_0 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_3_), .o(FE_RN_1050_0) );
in01f80 FE_OCP_RBC2491_n_3338 ( .a(FE_OCP_RBN2489_n_3338), .o(FE_OCP_RBN2491_n_3338) );
na02f80 g753529 ( .a(n_26821), .b(n_26820), .o(n_26912) );
in01f80 g758679 ( .a(n_21812), .o(n_21899) );
ao12f80 g775905 ( .a(n_4848), .b(n_4853), .c(n_4841), .o(n_5011) );
na02f80 g758937 ( .a(n_21236), .b(n_45081), .o(n_21291) );
in01f80 g779309 ( .a(FE_OFN812_n_2405), .o(n_1758) );
in01f80 g779170 ( .a(n_1901), .o(n_1902) );
in01f80 newInst_2672 ( .a(newNet_2671), .o(newNet_2672) );
in01f80 newInst_3480 ( .a(newNet_3479), .o(newNet_3480) );
oa12f80 g780427 ( .a(n_834), .b(n_1098), .c(FE_OFN50_n_1045), .o(n_937) );
na02f80 g752924 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_20_), .o(n_27813) );
oa22f80 FE_RC_2825_0 ( .a(n_9856), .b(n_9801), .c(n_9800), .d(n_9857), .o(n_10015) );
in01f80 g748147 ( .a(n_32161), .o(n_32162) );
in01f80 newInst_2205 ( .a(newNet_2204), .o(newNet_2205) );
na02f80 g739727 ( .a(n_40511), .b(n_40409), .o(n_40543) );
in01f80 g748885 ( .a(n_32414), .o(n_32415) );
na02f80 g750980 ( .a(n_30182), .b(n_29944), .o(n_30231) );
na02f80 g764988 ( .a(n_15607), .b(n_15580), .o(n_15753) );
no02f80 g743979 ( .a(n_35624), .b(n_35597), .o(n_35919) );
oa22f80 g774716 ( .a(n_6317), .b(n_5416), .c(n_6316), .d(n_5415), .o(n_6384) );
na02f80 g760098 ( .a(n_20275), .b(n_20293), .o(n_20914) );
in01f80 g768089 ( .a(n_13031), .o(n_13032) );
na02f80 g768755 ( .a(n_12177), .b(n_12176), .o(n_12178) );
na02f80 g741493 ( .a(n_38765), .b(n_38764), .o(n_38790) );
no02f80 g745275 ( .a(n_35606), .b(n_35635), .o(n_36681) );
in01f80 FE_RC_85_0 ( .a(FE_RN_26_0), .o(n_17395) );
na02f80 g773488 ( .a(n_7493), .b(n_6813), .o(n_7527) );
na02f80 g776127 ( .a(n_4524), .b(n_4534), .o(n_4692) );
in01f80 g778044 ( .a(n_3104), .o(n_3105) );
no02f80 g778061 ( .a(n_3016), .b(n_3494), .o(n_3028) );
no02f80 g748159 ( .a(n_32326), .b(n_32020), .o(n_32099) );
na02f80 g778690 ( .a(FE_OCP_RBN2295_n_2438), .b(n_2596), .o(n_2736) );
na02f80 g761050 ( .a(n_19183), .b(n_19154), .o(n_19270) );
in01f80 g745813 ( .a(n_34477), .o(n_34478) );
oa12f80 g756229 ( .a(n_24735), .b(n_24734), .c(n_24733), .o(n_24813) );
oa12f80 g736527 ( .a(n_43411), .b(n_43661), .c(n_43328), .o(n_43701) );
in01f80 newInst_3743 ( .a(newNet_3742), .o(newNet_3743) );
in01f80 g737828 ( .a(n_42216), .o(n_42367) );
oa12f80 g742855 ( .a(n_37238), .b(n_37237), .c(n_37236), .o(n_37274) );
ao22s80 g779024 ( .a(n_2163), .b(n_1932), .c(n_2147), .d(n_1931), .o(n_2204) );
no02f80 g779733 ( .a(n_1416), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_3_), .o(n_1521) );
na02f80 g776492 ( .a(n_4431), .b(n_4144), .o(n_4571) );
no02f80 g751833 ( .a(n_28264), .b(n_28371), .o(n_28369) );
na02f80 g745938 ( .a(n_35321), .b(n_35320), .o(n_35322) );
no02f80 g756552 ( .a(n_23678), .b(delay_add_ln22_unr14_stage6_stallmux_q_26_), .o(n_23853) );
ao12f80 g757631 ( .a(n_22308), .b(FE_OCP_RBN1195_n_22542), .c(n_22131), .o(n_22618) );
ao12f80 g738196 ( .a(n_41585), .b(n_41977), .c(n_41814), .o(n_41980) );
in01f80 FE_OCPC906_n_44561 ( .a(FE_OCP_RBN2617_n_44561), .o(FE_OCPN906_n_44561) );
no02f80 g767963 ( .a(n_13150), .b(n_12917), .o(n_13602) );
ao12f80 g766976 ( .a(n_13768), .b(n_13767), .c(n_13766), .o(n_13846) );
na02f80 g770234 ( .a(n_10629), .b(FE_OFN756_n_44461), .o(n_10735) );
in01f80 newInst_3673 ( .a(newNet_3672), .o(newNet_3673) );
ao12f80 g748679 ( .a(n_44042), .b(n_32451), .c(FE_OCPN1229_n_46101), .o(n_32645) );
no02f80 FE_RC_4233_0 ( .a(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .b(FE_RN_1858_0), .o(FE_RN_1859_0) );
in01f80 FE_RC_3031_0 ( .a(n_11810), .o(FE_RN_1327_0) );
oa12f80 g749672 ( .a(n_31639), .b(n_31638), .c(n_31637), .o(n_31689) );
no02f80 g769182 ( .a(n_12083), .b(n_12082), .o(n_12157) );
in01f80 FE_RC_3566_0 ( .a(FE_RN_1549_0), .o(n_29859) );
ao12f80 g756916 ( .a(n_23170), .b(n_23270), .c(n_23199), .o(n_23334) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_20_ ( .ck(newNet_721), .d(n_46182), .o(delay_xor_ln21_unr6_stage3_stallmux_q_20_) );
ao12f80 g758591 ( .a(n_21663), .b(n_21849), .c(n_21664), .o(n_21903) );
no02f80 g767059 ( .a(FE_OCP_RBN2458_n_13765), .b(n_13324), .o(n_13937) );
na02f80 g741200 ( .a(FE_OCP_RBN2685_n_38870), .b(FE_OCP_RBN2349_n_38515), .o(n_39100) );
oa22f80 FE_RC_2760_0 ( .a(n_32582), .b(n_32520), .c(FE_OCP_RBN1344_n_32520), .d(n_32522), .o(n_32638) );
no02f80 g748907 ( .a(n_32393), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_4_), .o(n_32391) );
na02f80 g771207 ( .a(n_9492), .b(n_9415), .o(n_9493) );
no02f80 g775344 ( .a(n_5909), .b(FE_OCPN1050_n_4459), .o(n_5982) );
na02f80 g737446 ( .a(n_42689), .b(n_42427), .o(n_42731) );
in01f80 newInst_722 ( .a(newNet_241), .o(newNet_722) );
na02f80 g768309 ( .a(n_12516), .b(n_12348), .o(n_12518) );
na02f80 g780600 ( .a(n_694), .b(n_719), .o(n_753) );
no02f80 g749410 ( .a(n_30514), .b(FE_OCP_RBN2634_n_30213), .o(n_30544) );
na02f80 g779793 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_15_), .o(n_1506) );
no02f80 g779092 ( .a(n_2061), .b(FE_OCP_RBN2199_n_2032), .o(n_2351) );
no02f80 g737926 ( .a(n_42270), .b(n_42500), .o(n_42514) );
na02f80 g780528 ( .a(n_677), .b(n_669), .o(n_689) );
na02f80 g778609 ( .a(n_2913), .b(n_2807), .o(n_2877) );
in01f80 FE_OCP_RBC2900_n_44853 ( .a(n_44853), .o(FE_OCP_RBN2900_n_44853) );
na02f80 g744986 ( .a(n_34921), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_34952) );
in01f80 g764337 ( .a(n_16741), .o(n_16768) );
no02f80 g747843 ( .a(n_33571), .b(n_33651), .o(n_33792) );
in01f80 g754485 ( .a(n_25597), .o(n_25631) );
no02f80 g759099 ( .a(n_21277), .b(n_21220), .o(n_21318) );
in01f80 FE_OCP_RBC2259_n_18899 ( .a(n_18899), .o(FE_OCP_RBN2259_n_18899) );
no02f80 g760461 ( .a(n_20094), .b(FE_RN_1248_0), .o(n_20160) );
no02f80 g744257 ( .a(FE_OCPN1510_n_44174), .b(n_36091), .o(n_36135) );
na02f80 g767949 ( .a(n_12775), .b(n_12774), .o(n_12788) );
no02f80 g738944 ( .a(n_41246), .b(n_40850), .o(n_41247) );
in01f80 g750415 ( .a(n_29615), .o(n_29626) );
in01f80 g774754 ( .a(n_6485), .o(n_6480) );
in01f80 g767192 ( .a(n_14730), .o(n_14805) );
in01f80 g768054 ( .a(n_13078), .o(n_13033) );
in01f80 g746829 ( .a(n_33100), .o(n_33101) );
no02f80 g775782 ( .a(n_5367), .b(n_5290), .o(n_5291) );
na02f80 g737616 ( .a(n_42239), .b(n_42223), .o(n_42251) );
no02f80 g739922 ( .a(n_40336), .b(n_40116), .o(n_40338) );
na02f80 g736792 ( .a(n_43054), .b(n_43036), .o(n_43068) );
no02f80 FE_RC_3061_0 ( .a(n_20404), .b(FE_OCP_RBN1696_n_19206), .o(FE_RN_1343_0) );
no02f80 FE_RC_2813_0 ( .a(FE_RN_1203_0), .b(FE_RN_1204_0), .o(n_9898) );
in01f80 g780683 ( .a(n_660), .o(n_661) );
na02f80 g776946 ( .a(n_3945), .b(n_3944), .o(n_3977) );
na02f80 g736745 ( .a(n_43187), .b(n_43315), .o(n_43188) );
no02f80 g760355 ( .a(n_20161), .b(n_20204), .o(n_20238) );
in01f80 newInst_175 ( .a(newNet_174), .o(newNet_175) );
in01f80 FE_OCP_RBC2345_FE_OCPN870_n_2737 ( .a(FE_OCP_RBN2343_FE_OCPN870_n_2737), .o(FE_OCP_RBN2345_FE_OCPN870_n_2737) );
na02f80 g742024 ( .a(n_37944), .b(n_37903), .o(n_38034) );
no02f80 g765515 ( .a(n_15565), .b(n_15564), .o(n_16135) );
na02f80 g762648 ( .a(n_18020), .b(n_17917), .o(n_18039) );
in01f80 g770184 ( .a(n_11013), .o(n_11014) );
no02f80 g742494 ( .a(n_37656), .b(n_37655), .o(n_37687) );
ao12f80 g779434 ( .a(n_1503), .b(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_7_), .o(n_1534) );
in01f80 g758850 ( .a(n_21505), .o(n_21548) );
oa12f80 g740880 ( .a(n_39145), .b(n_39113), .c(n_39062), .o(n_39220) );
in01f80 g751841 ( .a(n_29126), .o(n_29127) );
in01f80 g777670 ( .a(n_3414), .o(n_3389) );
no02f80 g759767 ( .a(n_21748), .b(n_21694), .o(n_21667) );
oa12f80 g776537 ( .a(n_4574), .b(n_4573), .c(n_4572), .o(n_4623) );
na02f80 g751946 ( .a(n_28167), .b(n_28222), .o(n_28300) );
oa12f80 g741729 ( .a(n_38051), .b(n_38421), .c(n_38087), .o(n_38499) );
in01f80 newInst_34 ( .a(newNet_32), .o(newNet_34) );
in01f80 g745084 ( .a(n_34870), .o(n_34871) );
na02f80 g764696 ( .a(n_15808), .b(n_15375), .o(n_15809) );
in01f80 g759023 ( .a(n_21238), .o(n_21237) );
in01f80 FE_OCP_RBC3427_n_44881 ( .a(FE_OCP_RBN3425_n_44881), .o(FE_OCP_RBN3427_n_44881) );
in01f80 FE_OCP_RBC2817_n_4458 ( .a(n_4458), .o(FE_OCP_RBN2817_n_4458) );
no02f80 g748432 ( .a(FE_OCP_RBN3712_n_31466), .b(n_31017), .o(n_31680) );
na02f80 g778396 ( .a(n_2467), .b(n_2466), .o(n_2505) );
ao12f80 g760476 ( .a(n_19949), .b(n_19950), .c(n_19948), .o(n_21763) );
no02f80 FE_RC_2655_0 ( .a(FE_RN_1107_0), .b(FE_RN_1108_0), .o(FE_RN_1109_0) );
in01f80 g774724 ( .a(n_6363), .o(n_6382) );
no02f80 g738148 ( .a(n_42025), .b(n_41770), .o(n_42105) );
in01f80 newInst_2276 ( .a(newNet_2275), .o(newNet_2276) );
in01f80 g777100 ( .a(n_3778), .o(n_3774) );
ao22s80 g736500 ( .a(n_43665), .b(n_43557), .c(n_43670), .d(n_43556), .o(n_43704) );
in01f80 g773645 ( .a(n_7307), .o(n_7308) );
no02f80 g740792 ( .a(n_39349), .b(n_39365), .o(n_39442) );
in01f80 g762993 ( .a(n_17417), .o(n_17494) );
na02f80 g771606 ( .a(n_44056), .b(n_9284), .o(n_9394) );
no02f80 g780449 ( .a(n_855), .b(n_521), .o(n_802) );
in01f80 newInst_2516 ( .a(newNet_2515), .o(newNet_2516) );
in01f80 newInst_348 ( .a(newNet_251), .o(newNet_348) );
in01f80 g774072 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n_7651) );
in01f80 newInst_641 ( .a(newNet_640), .o(newNet_641) );
in01f80 newInst_376 ( .a(newNet_375), .o(newNet_376) );
na02f80 g736533 ( .a(n_43661), .b(n_43409), .o(n_43709) );
no02f80 g751908 ( .a(n_28919), .b(n_29068), .o(n_29100) );
no02f80 g747593 ( .a(n_32198), .b(n_31703), .o(n_32243) );
no02f80 g746945 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_), .o(n_32961) );
na02f80 g746082 ( .a(n_33938), .b(FE_OCPN1766_n_33447), .o(n_33974) );
no02f80 FE_RC_1319_0 ( .a(FE_RN_389_0), .b(n_43162), .o(n_43287) );
ao12f80 g759559 ( .a(n_21797), .b(n_21800), .c(n_21714), .o(n_21883) );
in01f80 newInst_3214 ( .a(newNet_3213), .o(newNet_3214) );
in01f80 FE_OCP_RBC2554_n_44576 ( .a(FE_OCP_RBN3543_n_44575), .o(FE_OCP_RBN2554_n_44576) );
na02f80 g746155 ( .a(n_33807), .b(n_33305), .o(n_33852) );
oa22f80 FE_RC_1561_0 ( .a(n_28675), .b(n_28965), .c(n_28674), .d(n_28966), .o(n_29055) );
na02f80 g742719 ( .a(n_37369), .b(n_37368), .o(n_37370) );
in01f80 FE_RC_3863_0 ( .a(n_21847), .o(FE_RN_1688_0) );
ao12f80 g742165 ( .a(n_38274), .b(n_44887), .c(n_38273), .o(n_38390) );
in01f80 g760395 ( .a(n_20169), .o(n_20212) );
oa12f80 g784393 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_16_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46203) );
na02f80 g744098 ( .a(n_35612), .b(n_44174), .o(n_35663) );
na02f80 g737070 ( .a(n_43230), .b(n_43179), .o(n_43482) );
no02f80 g745995 ( .a(n_34427), .b(n_34037), .o(n_34038) );
no02f80 g745949 ( .a(n_35277), .b(n_34808), .o(n_35336) );
in01f80 g777748 ( .a(n_5178), .o(n_3380) );
no02f80 g765482 ( .a(n_15077), .b(n_14758), .o(n_15110) );
in01f80 g736493 ( .a(n_43689), .o(n_43690) );
in01f80 g767992 ( .a(n_12668), .o(n_12688) );
in01f80 g769666 ( .a(n_46986), .o(n_11412) );
no02f80 g769965 ( .a(n_10955), .b(n_10958), .o(n_10997) );
in01f80 newInst_3712 ( .a(newNet_3711), .o(newNet_3712) );
na02f80 g751998 ( .a(n_28897), .b(n_28987), .o(n_29023) );
in01f80 g761972 ( .a(n_19049), .o(n_19050) );
in01f80 newInst_326 ( .a(newNet_325), .o(newNet_326) );
no02f80 g747195 ( .a(n_33893), .b(n_33892), .o(n_33894) );
in01f80 fopt783235 ( .a(n_44769), .o(n_44775) );
in01f80 newInst_3038 ( .a(newNet_1646), .o(newNet_3038) );
oa12f80 g750520 ( .a(n_30002), .b(n_30441), .c(n_29998), .o(n_30475) );
na02f80 g747221 ( .a(n_32813), .b(n_32845), .o(n_32886) );
in01f80 newInst_2562 ( .a(newNet_970), .o(newNet_2562) );
no02f80 g763035 ( .a(n_17132), .b(n_17453), .o(n_17513) );
in01f80 FE_OCP_RBC2325_n_13616 ( .a(n_13616), .o(FE_OCP_RBN2325_n_13616) );
na02f80 g740430 ( .a(FE_OCP_RBN3031_n_39942), .b(n_39427), .o(n_40266) );
no02f80 g777292 ( .a(n_3604), .b(n_5062), .o(n_3714) );
in01f80 FE_OCP_RBC2535_n_47018 ( .a(FE_OCP_RBN2533_n_47018), .o(FE_OCP_RBN2535_n_47018) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_15_ ( .ck(newNet_3248), .d(n_36423), .o(delay_add_ln22_unr23_stage9_stallmux_q_15_) );
no02f80 g753832 ( .a(n_26338), .b(n_26337), .o(n_26413) );
oa12f80 g762170 ( .a(n_18066), .b(n_18194), .c(n_18016), .o(n_18247) );
in01f80 g755554 ( .a(n_24718), .o(n_24745) );
no02f80 g747665 ( .a(n_32169), .b(n_32168), .o(n_32170) );
in01f80 newInst_711 ( .a(newNet_710), .o(newNet_711) );
oa12f80 g758972 ( .a(n_22054), .b(n_22053), .c(n_22052), .o(n_22115) );
in01f80 newInst_1116 ( .a(newNet_224), .o(newNet_1116) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_21_ ( .ck(newNet_3416), .d(n_27728), .o(delay_add_ln22_unr17_stage7_stallmux_q_21_) );
na02f80 g760843 ( .a(n_19474), .b(n_19120), .o(n_19516) );
oa22f80 g780059 ( .a(n_1225), .b(n_825), .c(n_1226), .d(n_826), .o(n_1234) );
in01f80 g763743 ( .a(n_16733), .o(n_16734) );
in01f80 g781152 ( .a(n_206), .o(n_208) );
in01f80 g771135 ( .a(n_9664), .o(n_9665) );
ao12f80 g766570 ( .a(n_14393), .b(n_14435), .c(n_14392), .o(n_15669) );
na02f80 FE_RC_2254_0 ( .a(FE_RN_830_0), .b(n_18013), .o(FE_RN_831_0) );
no02f80 g774368 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_18_), .o(n_7097) );
na02f80 g775698 ( .a(n_5357), .b(n_5402), .o(n_5478) );
in01f80 newInst_2059 ( .a(newNet_2058), .o(newNet_2059) );
no02f80 g752816 ( .a(n_28280), .b(n_27953), .o(n_28278) );
na02f80 g760302 ( .a(n_20081), .b(n_20106), .o(n_20107) );
no02f80 g771655 ( .a(n_8885), .b(n_7571), .o(n_8939) );
in01f80 FE_OCPC1008_n_28439 ( .a(n_28439), .o(FE_OCPN1008_n_28439) );
in01f80 g742189 ( .a(n_38229), .o(n_38230) );
no02f80 g740826 ( .a(n_39402), .b(n_39074), .o(n_39464) );
oa12f80 g781109 ( .a(n_234), .b(n_233), .c(n_232), .o(n_417) );
na02f80 g754696 ( .a(n_26160), .b(n_25685), .o(n_26864) );
in01f80 g763471 ( .a(n_17025), .o(n_17026) );
no02f80 g752677 ( .a(n_28136), .b(n_28135), .o(n_28137) );
in01f80 newInst_2291 ( .a(newNet_2290), .o(newNet_2291) );
oa12f80 g765071 ( .a(n_15378), .b(n_15526), .c(n_15457), .o(n_15529) );
in01f80 newInst_1770 ( .a(newNet_1769), .o(newNet_1770) );
in01f80 newInst_769 ( .a(newNet_768), .o(newNet_769) );
na02f80 g763282 ( .a(n_17230), .b(n_17229), .o(n_17393) );
in01f80 newInst_3069 ( .a(newNet_3068), .o(newNet_3069) );
in01f80 newInst_1419 ( .a(newNet_1418), .o(newNet_1419) );
na02f80 g740179 ( .a(FE_OCP_RBN3719_n_39913), .b(n_40009), .o(n_40179) );
na02f80 g741719 ( .a(n_38478), .b(n_38085), .o(n_38479) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_9_ ( .ck(newNet_3267), .d(n_31561), .o(delay_add_ln22_unr20_stage8_stallmux_q_9_) );
na02f80 g747098 ( .a(n_32794), .b(n_32793), .o(n_32833) );
in01f80 FE_OCP_RBC3538_n_8597 ( .a(n_8597), .o(FE_OCP_RBN3538_n_8597) );
in01f80 newInst_510 ( .a(newNet_509), .o(newNet_510) );
na02f80 g775824 ( .a(n_5049), .b(FE_OCP_RBN2728_n_4219), .o(n_5070) );
in01f80 g754944 ( .a(n_25668), .o(n_25669) );
ao12f80 g769242 ( .a(n_11709), .b(n_11707), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_12_), .o(n_12241) );
na02f80 g747001 ( .a(n_32990), .b(n_32989), .o(n_33052) );
oa22f80 g744914 ( .a(n_34990), .b(n_34743), .c(n_34991), .d(n_34744), .o(n_35092) );
na02f80 g770653 ( .a(n_10307), .b(n_10260), .o(n_10465) );
no02f80 g771443 ( .a(n_9317), .b(n_9269), .o(n_9406) );
in01f80 g770588 ( .a(n_47263), .o(n_10276) );
in01f80 g761086 ( .a(n_20039), .o(n_20040) );
oa12f80 g753434 ( .a(n_26387), .b(n_26987), .c(n_26985), .o(n_27008) );
no02f80 g780068 ( .a(n_1222), .b(n_843), .o(n_1223) );
na02f80 g772330 ( .a(n_8771), .b(n_8715), .o(n_8806) );
oa22f80 g749536 ( .a(n_31752), .b(n_31535), .c(n_31780), .d(n_31534), .o(n_31856) );
na02f80 g760185 ( .a(n_20429), .b(n_19472), .o(n_20712) );
no02f80 g770883 ( .a(n_10013), .b(n_9636), .o(n_10014) );
in01f80 newInst_2017 ( .a(newNet_980), .o(newNet_2017) );
ao22s80 g736449 ( .a(n_43718), .b(n_43321), .c(n_43717), .d(n_43322), .o(n_43757) );
in01f80 g758629 ( .a(n_21918), .o(n_21919) );
in01f80 g765978 ( .a(n_14754), .o(n_14698) );
in01f80 g759417 ( .a(n_20917), .o(n_20918) );
na02f80 g777806 ( .a(n_3224), .b(n_2735), .o(n_3306) );
oa12f80 g747143 ( .a(n_32713), .b(n_32707), .c(n_32711), .o(n_32794) );
no02f80 g737663 ( .a(n_42392), .b(n_42562), .o(n_42583) );
in01f80 newInst_566 ( .a(newNet_565), .o(newNet_566) );
na02f80 g755664 ( .a(n_24522), .b(n_24552), .o(n_24683) );
na02f80 g779373 ( .a(n_1585), .b(delay_add_ln22_unr2_stage2_stallmux_q_1_), .o(n_1608) );
in01f80 g768894 ( .a(n_11944), .o(n_12724) );
na02f80 g772320 ( .a(n_8722), .b(n_8721), .o(n_8723) );
na02f80 g737437 ( .a(n_42703), .b(n_42577), .o(n_42736) );
in01f80 g756475 ( .a(n_23881), .o(n_23882) );
no02f80 g767311 ( .a(n_13496), .b(n_13495), .o(n_13569) );
in01f80 g738052 ( .a(n_42144), .o(n_42350) );
in01f80 FE_OCP_RBC3554_n_44575 ( .a(FE_OCP_RBN3546_n_44575), .o(FE_OCP_RBN3554_n_44575) );
na02f80 g744952 ( .a(n_34974), .b(n_34952), .o(n_35046) );
in01f80 FE_OCP_RBC1846_n_22068 ( .a(n_22068), .o(FE_OCP_RBN1846_n_22068) );
in01f80 newInst_3233 ( .a(newNet_3027), .o(newNet_3233) );
no02f80 g737431 ( .a(n_42671), .b(n_42575), .o(n_42690) );
in01f80 g743917 ( .a(n_35869), .o(n_35870) );
na02f80 g745318 ( .a(n_36117), .b(n_35722), .o(n_36167) );
in01f80 g758933 ( .a(n_21542), .o(n_21577) );
in01f80 newInst_3079 ( .a(newNet_209), .o(newNet_3079) );
no02f80 g742128 ( .a(n_37891), .b(n_37809), .o(n_37951) );
no03m80 FE_RC_1659_0 ( .a(n_33717), .b(n_34560), .c(n_33828), .o(n_33882) );
no02f80 FE_RC_2413_0 ( .a(n_1976), .b(FE_RN_951_0), .o(FE_RN_952_0) );
na02f80 g750775 ( .a(n_29164), .b(n_28734), .o(n_29218) );
na02f80 g771070 ( .a(n_9715), .b(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .o(n_9743) );
in01f80 g746761 ( .a(n_33203), .o(n_33188) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_20_ ( .ck(newNet_821), .d(n_1354), .o(delay_xor_ln21_unr3_stage2_stallmux_q_20_) );
no02f80 g741054 ( .a(n_39004), .b(n_38548), .o(n_39005) );
in01f80 g741127 ( .a(n_39046), .o(n_39047) );
na02f80 g776113 ( .a(n_44862), .b(n_4466), .o(n_4994) );
na02f80 g755086 ( .a(n_25717), .b(n_25716), .o(n_25718) );
in01f80 newInst_2906 ( .a(newNet_1915), .o(newNet_2906) );
no02f80 g770131 ( .a(n_10810), .b(n_44464), .o(n_10823) );
in01f80 FE_RC_1185_0 ( .a(n_13689), .o(FE_RN_358_0) );
in01f80 newInst_3645 ( .a(newNet_3554), .o(newNet_3645) );
na02f80 g737556 ( .a(n_42266), .b(n_42267), .o(n_42268) );
na02f80 g746246 ( .a(n_35072), .b(n_35071), .o(n_35073) );
no02f80 g743260 ( .a(n_36844), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_1_), .o(n_36883) );
na02f80 g738849 ( .a(n_41288), .b(n_41287), .o(n_41289) );
na02f80 g745822 ( .a(n_44104), .b(n_34160), .o(n_34177) );
no02f80 g737476 ( .a(n_42565), .b(n_42661), .o(n_42686) );
in01f80 newInst_2731 ( .a(newNet_2730), .o(newNet_2731) );
na02f80 g749314 ( .a(n_30758), .b(n_29441), .o(n_30799) );
in01f80 g745479 ( .a(FE_OCP_RBN2995_n_35539), .o(n_36049) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_11_ ( .ck(newNet_525), .d(n_22908), .o(delay_xor_ln22_unr15_stage6_stallmux_q_11_) );
in01f80 g780537 ( .a(n_855), .o(n_764) );
no02f80 g750744 ( .a(n_29299), .b(n_29267), .o(n_29268) );
na02f80 FE_RC_2945_0 ( .a(FE_RN_1283_0), .b(FE_OCP_RBN2752_n_15461), .o(FE_RN_1285_0) );
na02f80 g769356 ( .a(n_11507), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_9_), .o(n_11570) );
no02f80 g750455 ( .a(n_29524), .b(n_30191), .o(n_29575) );
oa12f80 g752745 ( .a(n_28204), .b(n_27880), .c(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27959) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_24_ ( .ck(newNet_2089), .d(n_6435), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_) );
in01f80 g741087 ( .a(n_39107), .o(n_39051) );
in01f80 FE_OCP_RBC1849_n_22639 ( .a(n_22639), .o(FE_OCP_RBN1849_n_22639) );
na02f80 g771831 ( .a(n_9728), .b(n_9730), .o(n_10491) );
in01f80 g744860 ( .a(n_35099), .o(n_35100) );
in01f80 g776755 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n_4373) );
na02f80 g765641 ( .a(n_15019), .b(n_15043), .o(n_15044) );
in01f80 g767821 ( .a(n_13381), .o(n_13280) );
in01f80 FE_OCP_DRV_C1562_n_19562 ( .a(FE_OCP_DRV_N1561_n_19562), .o(FE_OCP_DRV_N1562_n_19562) );
ao12f80 g751004 ( .a(n_28505), .b(n_28853), .c(n_28474), .o(n_28872) );
in01f80 FE_OCP_RBC2305_n_7817 ( .a(FE_OCP_RBN2303_n_7817), .o(FE_OCP_RBN2305_n_7817) );
in01f80 g772563 ( .a(n_8426), .o(n_8427) );
in01f80 g757267 ( .a(n_23488), .o(n_23489) );
ao12f80 g745394 ( .a(n_34490), .b(n_34404), .c(n_34369), .o(n_34491) );
na02f80 g749604 ( .a(n_31582), .b(n_31222), .o(n_31672) );
ao12f80 g753921 ( .a(n_26126), .b(n_26267), .c(n_26127), .o(n_26412) );
oa12f80 g738281 ( .a(n_41889), .b(n_41888), .c(n_41887), .o(n_41947) );
in01f80 FE_OCP_RBC2783_n_9859 ( .a(n_9859), .o(FE_OCP_RBN2783_n_9859) );
na02f80 g778228 ( .a(n_2718), .b(n_2717), .o(n_2816) );
in01f80 newInst_3144 ( .a(newNet_978), .o(newNet_3144) );
oa12f80 g745252 ( .a(n_34265), .b(n_34275), .c(n_34264), .o(n_34327) );
no02f80 g768545 ( .a(n_12316), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_8_), .o(n_12346) );
na02f80 g744484 ( .a(n_35424), .b(n_35358), .o(n_35458) );
no03m80 FE_RC_3002_0 ( .a(n_15114), .b(n_15356), .c(n_15358), .o(n_15510) );
in01f80 newInst_762 ( .a(newNet_761), .o(newNet_762) );
na02f80 g763155 ( .a(n_17789), .b(n_17788), .o(n_17790) );
na02f80 FE_RC_1324_0 ( .a(FE_RN_390_0), .b(FE_RN_391_0), .o(FE_RN_392_0) );
no02f80 g741139 ( .a(n_39129), .b(n_38981), .o(n_39151) );
no02f80 g747419 ( .a(FE_OCP_RBN3331_n_44962), .b(delay_xor_ln21_unr21_stage8_stallmux_q_5_), .o(n_32436) );
no02f80 g748302 ( .a(n_31560), .b(n_31559), .o(n_31608) );
in01f80 g754336 ( .a(n_26688), .o(n_26689) );
in01f80 FE_OCPC1745_n_29420 ( .a(n_29420), .o(FE_OCPN1745_n_29420) );
in01f80 fopt783663 ( .a(n_45312), .o(n_45311) );
in01f80 g743179 ( .a(n_45896), .o(n_38193) );
in01f80 FE_OCP_RBC2254_n_33729 ( .a(n_33729), .o(FE_OCP_RBN2254_n_33729) );
na02f80 g744134 ( .a(n_36188), .b(n_35588), .o(n_36240) );
oa12f80 g767910 ( .a(n_12765), .b(n_12700), .c(FE_OCP_RBN1925_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_12863) );
no02f80 g767793 ( .a(n_12744), .b(n_11868), .o(n_12870) );
in01f80 newInst_2966 ( .a(newNet_2965), .o(newNet_2966) );
no02f80 g744148 ( .a(n_47265), .b(n_35974), .o(n_36004) );
na02f80 g771225 ( .a(n_9639), .b(n_9447), .o(n_9793) );
in01f80 newInst_690 ( .a(newNet_496), .o(newNet_690) );
in01f80 g775805 ( .a(n_5549), .o(n_5550) );
no02f80 g738043 ( .a(n_42110), .b(n_42119), .o(n_42323) );
na02f80 g754079 ( .a(n_26069), .b(n_25624), .o(n_26071) );
no02f80 g738568 ( .a(n_41534), .b(n_41879), .o(n_41618) );
ao12f80 g762631 ( .a(n_18257), .b(n_18256), .c(n_18255), .o(n_18521) );
in01f80 FE_OCP_RBC2474_n_8664 ( .a(FE_OCP_RBN2473_n_8664), .o(FE_OCP_RBN2474_n_8664) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_3_ ( .ck(newNet_700), .d(n_46156), .o(delay_xor_ln21_unr6_stage3_stallmux_q_3_) );
no02f80 g746931 ( .a(n_32863), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_15_), .o(n_32949) );
na02f80 g751271 ( .a(n_29758), .b(n_29757), .o(n_29759) );
ao12f80 g760161 ( .a(n_20014), .b(n_20929), .c(n_19906), .o(n_20988) );
in01f80 g769995 ( .a(n_11055), .o(n_11098) );
na02f80 FE_RC_2330_0 ( .a(FE_RN_885_0), .b(FE_RN_889_0), .o(n_33484) );
in01f80 g763180 ( .a(n_18479), .o(n_18744) );
oa12f80 g743939 ( .a(n_36900), .b(n_36556), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37434) );
na02f80 g761273 ( .a(n_19931), .b(n_19787), .o(n_19956) );
na02f80 g763350 ( .a(n_17708), .b(n_17665), .o(n_17710) );
in01f80 newInst_2668 ( .a(newNet_2667), .o(newNet_2668) );
in01f80 FE_OCP_RBC3484_n_13667 ( .a(FE_OCP_RBN3483_n_13667), .o(FE_OCP_RBN3484_n_13667) );
in01f80 g739831 ( .a(n_40450), .o(n_40451) );
oa12f80 g766802 ( .a(n_13864), .b(n_13943), .c(n_13939), .o(n_14011) );
in01f80 g740533 ( .a(n_39685), .o(n_39686) );
in01f80 newInst_584 ( .a(newNet_583), .o(newNet_584) );
in01f80 g763534 ( .a(n_16976), .o(n_17022) );
na02f80 g761927 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_25_), .o(n_18467) );
oa22f80 g763130 ( .a(n_17199), .b(n_17336), .c(n_17142), .d(n_17753), .o(n_17291) );
in01f80 g739962 ( .a(n_40228), .o(n_40196) );
no02f80 g758112 ( .a(n_44277), .b(FE_OCP_RBN1913_n_20965), .o(n_22099) );
in01f80 FE_RC_144_0 ( .a(n_12038), .o(FE_RN_42_0) );
in01f80 FE_OCP_RBC2955_n_26231 ( .a(FE_OCP_RBN2954_n_26231), .o(FE_OCP_RBN2955_n_26231) );
in01f80 g754849 ( .a(n_25509), .o(n_25510) );
in01f80 newInst_402 ( .a(newNet_289), .o(newNet_402) );
oa12f80 g748729 ( .a(n_46107), .b(n_32405), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_27_), .o(n_32538) );
oa22f80 FE_RC_405_0 ( .a(n_13332), .b(FE_OCP_RBN3429_n_13245), .c(n_13245), .d(n_13294), .o(n_13398) );
in01f80 g738947 ( .a(n_41195), .o(n_41196) );
ms00f80 delay_xor_ln22_unr28_stage10_stallmux_q_reg_0_ ( .ck(newNet_386), .d(n_40580), .o(delay_xor_ln22_unr28_stage10_stallmux_q_0_) );
na02f80 g746586 ( .a(n_34612), .b(n_34227), .o(n_34776) );
no02f80 g752038 ( .a(n_28118), .b(n_28028), .o(n_28168) );
in01f80 g775897 ( .a(n_5121), .o(n_5122) );
in01f80 newInst_1057 ( .a(newNet_180), .o(newNet_1057) );
in01f80 FE_OFC774_n_46137 ( .a(FE_OFN773_n_46137), .o(FE_OFN774_n_46137) );
oa12f80 g778005 ( .a(n_2389), .b(n_3008), .c(n_2449), .o(n_3045) );
no02f80 g749710 ( .a(n_31349), .b(n_31224), .o(n_31351) );
in01f80 g753557 ( .a(n_27449), .o(n_27450) );
in01f80 newInst_1894 ( .a(newNet_1175), .o(newNet_1894) );
na02f80 g750687 ( .a(n_30359), .b(n_30358), .o(n_30360) );
in01f80 g750218 ( .a(n_29846), .o(n_29869) );
no02f80 g766873 ( .a(n_14347), .b(n_14345), .o(n_14346) );
no02f80 g737332 ( .a(n_42832), .b(n_42841), .o(n_43181) );
in01f80 g749541 ( .a(n_30496), .o(n_30497) );
in01f80 newInst_505 ( .a(newNet_504), .o(newNet_505) );
no02f80 g738929 ( .a(n_41197), .b(n_40995), .o(n_41273) );
na02f80 g776240 ( .a(n_4811), .b(n_4287), .o(n_4894) );
na02f80 g773156 ( .a(n_7576), .b(n_7321), .o(n_7654) );
oa22f80 FE_RC_19_0 ( .a(FE_OFN806_n_46196), .b(n_6720), .c(FE_OFN84_n_46137), .d(n_44823), .o(n_46192) );
in01f80 fopt783493 ( .a(n_45066), .o(n_45101) );
no02f80 g770708 ( .a(n_10098), .b(n_10061), .o(n_10270) );
na02f80 g746579 ( .a(n_34666), .b(n_34580), .o(n_35041) );
in01f80 g751590 ( .a(n_28543), .o(n_28626) );
na02f80 g754212 ( .a(n_25939), .b(n_25919), .o(n_25972) );
oa12f80 g771500 ( .a(n_9559), .b(n_9595), .c(n_9558), .o(n_9653) );
in01f80 newInst_274 ( .a(newNet_273), .o(newNet_274) );
no02f80 g748760 ( .a(n_31057), .b(n_29678), .o(n_31162) );
na02f80 g745261 ( .a(n_34513), .b(n_34491), .o(n_34591) );
oa12f80 g742725 ( .a(n_37303), .b(n_37302), .c(n_37301), .o(n_37849) );
oa22f80 g784345 ( .a(FE_OCP_RBN3077_FE_OFN807_n_46195), .b(n_6248), .c(FE_OFN774_n_46137), .d(n_6206), .o(n_46151) );
no02f80 g781309 ( .a(beta_31), .b(beta_9), .o(n_57) );
na02f80 g778708 ( .a(n_2365), .b(n_2432), .o(n_2710) );
na02f80 g758012 ( .a(n_22225), .b(n_22232), .o(n_22338) );
no02f80 g778369 ( .a(n_2782), .b(delay_add_ln22_unr2_stage2_stallmux_q_27_), .o(n_2818) );
oa12f80 g778644 ( .a(n_2241), .b(n_2240), .c(n_2239), .o(n_3084) );
oa12f80 g749628 ( .a(n_30227), .b(n_30226), .c(n_30225), .o(n_30299) );
in01f80 newInst_1803 ( .a(newNet_1802), .o(newNet_1803) );
oa22f80 g763873 ( .a(n_17158), .b(FE_OCP_RBN3359_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .c(n_17256), .d(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_), .o(n_17788) );
in01f80 FE_OCP_RBC1345_n_19270 ( .a(n_19270), .o(FE_OCP_RBN1345_n_19270) );
in01f80 g748741 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_3_), .o(n_31181) );
no02f80 g773435 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_27_), .o(n_7614) );
no02f80 g767617 ( .a(n_13100), .b(n_12842), .o(n_13136) );
no02f80 g741479 ( .a(n_38753), .b(n_38752), .o(n_38761) );
oa22f80 g746730 ( .a(n_32951), .b(n_32831), .c(n_32980), .d(n_32832), .o(n_34182) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_16_ ( .ck(newNet_3546), .d(n_22479), .o(delay_add_ln22_unr14_stage6_stallmux_q_16_) );
ao12f80 g762457 ( .a(n_18051), .b(FE_OCP_RBN2142_FE_OCPN861_n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_13_), .o(n_18001) );
no02f80 g778121 ( .a(n_2805), .b(n_2227), .o(n_2806) );
in01f80 FE_RC_2466_0 ( .a(n_13970), .o(FE_RN_991_0) );
in01f80 g778410 ( .a(n_2664), .o(n_3274) );
ao12f80 g760104 ( .a(n_20029), .b(n_20107), .c(n_20006), .o(n_20195) );
na02f80 g760663 ( .a(FE_OCP_RBN1181_n_19726), .b(n_19557), .o(n_19860) );
in01f80 newInst_652 ( .a(newNet_651), .o(newNet_652) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_26_ ( .ck(newNet_1496), .d(n_32291), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_26_) );
na02f80 g766100 ( .a(n_14636), .b(n_14579), .o(n_14659) );
in01f80 g777145 ( .a(n_3695), .o(n_3696) );
no02f80 g776581 ( .a(n_4050), .b(n_4033), .o(n_4138) );
in01f80 g764012 ( .a(n_18119), .o(n_18140) );
in01f80 g781193 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_24105) );
in01f80 FE_OCP_RBC3358_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(FE_OCP_RBN3296_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3358_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
in01f80 g769019 ( .a(n_11698), .o(n_11654) );
no02f80 g771334 ( .a(n_9564), .b(n_9609), .o(n_9794) );
no02f80 g767581 ( .a(n_13178), .b(n_13177), .o(n_13179) );
in01f80 newInst_1830 ( .a(newNet_1829), .o(newNet_1830) );
in01f80 g754878 ( .a(n_25247), .o(n_25280) );
na02f80 g739973 ( .a(n_40023), .b(n_40045), .o(n_40085) );
no02f80 g760954 ( .a(n_19282), .b(n_19331), .o(n_19467) );
na02f80 g758271 ( .a(FE_OCPN992_n_22249), .b(FE_OCP_RBN1712_n_21087), .o(n_22375) );
ao12f80 g757929 ( .a(FE_OCP_RBN2112_n_22650), .b(n_22785), .c(n_22728), .o(n_22854) );
in01f80 g776173 ( .a(n_4717), .o(n_4676) );
in01f80 newInst_3407 ( .a(newNet_3406), .o(newNet_3407) );
in01f80 g739160 ( .a(n_40957), .o(n_40989) );
ao22s80 FE_RC_993_0 ( .a(n_44061), .b(FE_OCP_RBN2051_delay_xor_ln22_unr15_stage6_stallmux_q_2_), .c(delay_xor_ln22_unr15_stage6_stallmux_q_2_), .d(FE_OCP_RBN3823_n_44061), .o(n_22771) );
no02f80 FE_RC_1010_0 ( .a(FE_RN_293_0), .b(n_17736), .o(n_17787) );
no02f80 g740057 ( .a(n_40042), .b(n_40001), .o(n_40040) );
na02f80 g777176 ( .a(n_4599), .b(n_4739), .o(n_5413) );
no02f80 g740256 ( .a(n_39912), .b(n_39965), .o(n_39966) );
in01f80 newInst_3357 ( .a(newNet_1680), .o(newNet_3357) );
na02f80 FE_RC_1746_0 ( .a(n_12293), .b(FE_RN_490_0), .o(FE_RN_491_0) );
in01f80 FE_OCP_RBC2668_n_4158 ( .a(FE_OCP_RBN2667_n_4158), .o(FE_OCP_RBN2668_n_4158) );
in01f80 newInst_2796 ( .a(newNet_975), .o(newNet_2796) );
no02f80 g737683 ( .a(n_42392), .b(n_42112), .o(n_42527) );
na02f80 g750373 ( .a(n_29667), .b(n_29666), .o(n_29668) );
na02f80 g756039 ( .a(n_24981), .b(n_24980), .o(n_24997) );
no02f80 g753487 ( .a(n_26851), .b(n_26850), .o(n_26960) );
in01f80 g760958 ( .a(n_19255), .o(n_19256) );
in01f80 FE_OCP_RBC2196_n_2103 ( .a(n_2103), .o(FE_OCP_RBN2196_n_2103) );
na02f80 g756776 ( .a(n_23396), .b(n_23144), .o(n_23425) );
no02f80 g767065 ( .a(FE_OCP_RBN2459_n_13765), .b(n_13893), .o(n_13897) );
in01f80 g744966 ( .a(n_35905), .o(n_34954) );
ao12f80 g784613 ( .a(n_42752), .b(n_42734), .c(n_42712), .o(n_46941) );
na02f80 g779744 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n_1751) );
no02f80 g749943 ( .a(n_30116), .b(n_29167), .o(n_30117) );
no02f80 FE_RC_2591_0 ( .a(FE_RN_1071_0), .b(FE_RN_1070_0), .o(FE_RN_1072_0) );
na02f80 g753585 ( .a(n_26629), .b(n_26592), .o(n_26698) );
na02f80 FE_RC_3038_0 ( .a(n_11476), .b(FE_RN_1330_0), .o(n_11582) );
no02f80 g754495 ( .a(n_26714), .b(n_26644), .o(n_26715) );
in01f80 newInst_2616 ( .a(newNet_2615), .o(newNet_2616) );
in01f80 newInst_2266 ( .a(newNet_1228), .o(newNet_2266) );
no02f80 g774076 ( .a(n_6724), .b(n_6652), .o(n_6790) );
in01f80 g748917 ( .a(n_32390), .o(n_32448) );
no02f80 g736862 ( .a(n_43304), .b(n_43508), .o(n_43613) );
no02f80 g745999 ( .a(n_34003), .b(n_34033), .o(n_34034) );
in01f80 g762441 ( .a(n_18071), .o(n_18072) );
in01f80 g772614 ( .a(n_8337), .o(n_8324) );
no02f80 g746160 ( .a(n_33697), .b(n_34037), .o(n_33717) );
in01f80 g780317 ( .a(n_979), .o(n_980) );
in01f80 g769976 ( .a(n_11043), .o(n_11044) );
oa22f80 FE_RC_3921_0 ( .a(n_27681), .b(n_27399), .c(n_27682), .d(n_27398), .o(n_27772) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_15_ ( .ck(newNet_507), .d(n_22947), .o(delay_xor_ln22_unr15_stage6_stallmux_q_15_) );
ao22s80 FE_RC_120_0 ( .a(n_45065), .b(n_20325), .c(n_20326), .d(n_45066), .o(n_20435) );
na02f80 FE_RC_2658_0 ( .a(n_7802), .b(FE_RN_1110_0), .o(FE_RN_1111_0) );
in01f80 newInst_2527 ( .a(newNet_2206), .o(newNet_2527) );
no02f80 g759429 ( .a(n_20973), .b(FE_OCP_RBN2739_n_20432), .o(n_20972) );
no02f80 g761654 ( .a(n_19494), .b(n_18883), .o(n_19545) );
in01f80 g757069 ( .a(n_23359), .o(n_23360) );
na02f80 g740448 ( .a(n_39717), .b(n_39689), .o(n_39726) );
na02f80 g749201 ( .a(n_30739), .b(n_30386), .o(n_30828) );
no02f80 g760144 ( .a(n_20456), .b(FE_OCP_RBN1703_n_19560), .o(n_20667) );
oa22f80 FE_RC_899_0 ( .a(n_25380), .b(n_25632), .c(n_25354), .d(n_25600), .o(n_25731) );
na02f80 g770757 ( .a(FE_OCP_RBN3653_n_10100), .b(n_9162), .o(n_10245) );
no03m80 g743786 ( .a(n_46205), .b(n_46253), .c(n_46221), .o(n_37284) );
na02f80 g769319 ( .a(FE_OCPN858_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_20_), .o(n_12016) );
oa12f80 g763138 ( .a(n_17790), .b(n_17789), .c(n_17788), .o(n_17859) );
no02f80 g778467 ( .a(n_2570), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_), .o(n_2601) );
na02f80 g781045 ( .a(cos_out_18), .b(n_43918), .o(n_315) );
no02f80 g779150 ( .a(n_1993), .b(n_1706), .o(n_2025) );
oa12f80 g751872 ( .a(n_28247), .b(n_28221), .c(n_28220), .o(n_28362) );
na02f80 g758141 ( .a(n_22463), .b(n_22330), .o(n_22464) );
na02f80 g752808 ( .a(n_28156), .b(n_28174), .o(n_28710) );
na02f80 g758175 ( .a(n_44268), .b(n_21264), .o(n_22216) );
in01f80 g756249 ( .a(n_24139), .o(n_24140) );
no02f80 FE_RC_1052_0 ( .a(FE_RN_306_0), .b(FE_RN_307_0), .o(FE_RN_308_0) );
no02f80 g749688 ( .a(n_31395), .b(n_31346), .o(n_31418) );
no02f80 g736981 ( .a(FE_OCPN1246_n_43120), .b(n_43061), .o(n_43504) );
in01f80 newInst_617 ( .a(newNet_616), .o(newNet_617) );
in01f80 g770725 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .o(n_10371) );
ao12f80 g754478 ( .a(n_26381), .b(n_26418), .c(FE_OCP_RBN2957_n_26231), .o(n_26514) );
in01f80 g752947 ( .a(n_27926), .o(n_27810) );
no02f80 g756276 ( .a(n_24665), .b(n_24664), .o(n_24666) );
in01f80 newInst_1250 ( .a(newNet_1249), .o(newNet_1250) );
no02f80 g773212 ( .a(n_7730), .b(n_7690), .o(n_7759) );
oa12f80 g746868 ( .a(n_32877), .b(n_32876), .c(n_32875), .o(n_34085) );
in01f80 FE_RC_1997_0 ( .a(n_24281), .o(FE_RN_654_0) );
in01f80 newInst_2426 ( .a(newNet_2425), .o(newNet_2426) );
no02f80 g759909 ( .a(n_21053), .b(n_21052), .o(n_21172) );
in01f80 g771680 ( .a(n_10124), .o(n_10210) );
in01f80 g739341 ( .a(n_40692), .o(n_40730) );
in01f80 g750403 ( .a(n_29658), .o(n_29659) );
in01f80 g748190 ( .a(n_31524), .o(n_31525) );
in01f80 g745429 ( .a(n_35839), .o(n_35996) );
na02f80 g783824 ( .a(FE_OCP_RBN3356_delay_xor_ln22_unr28_stage10_stallmux_q_0_), .b(n_44610), .o(n_45511) );
in01f80 g765947 ( .a(n_15128), .o(n_15210) );
in01f80 newInst_629 ( .a(newNet_628), .o(newNet_629) );
in01f80 g778403 ( .a(n_2537), .o(n_2585) );
na02f80 g745765 ( .a(n_34053), .b(n_34069), .o(n_34054) );
na02f80 g764376 ( .a(n_16231), .b(FE_OCPN3775_n_14730), .o(n_16373) );
ao12f80 g754734 ( .a(n_25214), .b(n_25366), .c(n_25183), .o(n_25432) );
in01f80 g775978 ( .a(n_5169), .o(n_5170) );
no02f80 g741327 ( .a(FE_OCP_RBN2546_n_44944), .b(FE_OCP_RBN2452_n_38537), .o(n_39120) );
no03m80 FE_RC_1685_0 ( .a(n_33782), .b(FE_OCP_RBN1355_n_44259), .c(FE_OCP_RBN2261_n_33691), .o(n_33784) );
oa12f80 g739023 ( .a(n_41179), .b(n_41178), .c(n_41177), .o(n_41218) );
no03m80 FE_RC_1132_0 ( .a(FE_OCPN1020_n_23078), .b(n_23047), .c(FE_RN_155_0), .o(n_23194) );
no02f80 g759430 ( .a(n_21144), .b(n_21056), .o(n_21207) );
na02f80 g775728 ( .a(n_5550), .b(n_4076), .o(n_5658) );
in01f80 FE_OCPC853_n_45450 ( .a(n_45450), .o(FE_OCPN853_n_45450) );
in01f80 g742561 ( .a(n_37593), .o(n_37594) );
in01f80 FE_OCP_RBC3419_n_12739 ( .a(FE_OCP_RBN3417_n_12739), .o(FE_OCP_RBN3419_n_12739) );
no02f80 g755401 ( .a(n_24894), .b(n_24893), .o(n_24913) );
no02f80 g740679 ( .a(n_39553), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39570) );
in01f80 g759697 ( .a(n_20640), .o(n_20639) );
na02f80 g761871 ( .a(n_47246), .b(n_18470), .o(n_18513) );
in01f80 newInst_2861 ( .a(newNet_971), .o(newNet_2861) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_8_ ( .ck(newNet_606), .d(n_46374), .o(delay_xor_ln21_unr9_stage4_stallmux_q_8_) );
na02f80 g778205 ( .a(n_2750), .b(n_2816), .o(n_2969) );
no02f80 g746240 ( .a(n_33531), .b(n_33104), .o(n_33595) );
no02f80 g745875 ( .a(n_35356), .b(n_35355), .o(n_35357) );
oa22f80 FE_RC_2961_0 ( .a(n_10845), .b(n_10905), .c(n_10904), .d(n_10846), .o(n_11017) );
na02f80 g739057 ( .a(n_41075), .b(n_41074), .o(n_41076) );
in01f80 FE_OCP_RBC2124_n_45224 ( .a(FE_OCP_RBN2122_n_45224), .o(FE_OCP_RBN2124_n_45224) );
in01f80 newInst_3552 ( .a(newNet_3551), .o(newNet_3552) );
ao12f80 g742885 ( .a(n_37082), .b(n_44021), .c(n_36470), .o(n_37081) );
no02f80 g750345 ( .a(n_29686), .b(n_29701), .o(n_29766) );
in01f80 g740493 ( .a(n_39787), .o(n_39803) );
no02f80 g743371 ( .a(n_37830), .b(n_46243), .o(n_37805) );
in01f80 g750968 ( .a(n_30183), .o(n_30184) );
no02f80 g768638 ( .a(n_12199), .b(n_12198), .o(n_12200) );
in01f80 g765075 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_2_), .o(n_17018) );
na02f80 g771141 ( .a(n_9623), .b(FE_OCPN3769_FE_OCP_RBN2375_n_8221), .o(n_9740) );
oa22f80 g764185 ( .a(n_16824), .b(n_16306), .c(n_16848), .d(n_16307), .o(n_16849) );
no02f80 g738698 ( .a(n_41716), .b(n_41401), .o(n_41760) );
no02f80 g739304 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n_40988) );
na02f80 g770229 ( .a(n_10709), .b(n_44463), .o(n_10727) );
in01f80 FE_OCP_RBC3374_n_6745 ( .a(FE_OCP_RBN2127_n_6745), .o(FE_OCP_RBN3374_n_6745) );
no02f80 g747161 ( .a(n_33952), .b(n_33933), .o(n_33934) );
na02f80 g737392 ( .a(n_42780), .b(n_43132), .o(n_42781) );
in01f80 FE_OCP_RBC2883_n_26292 ( .a(n_26292), .o(FE_OCP_RBN2883_n_26292) );
na02f80 g755231 ( .a(n_44445), .b(n_24804), .o(n_25019) );
no02f80 g777278 ( .a(FE_OCP_RBN2731_n_4219), .b(n_4537), .o(n_4685) );
in01f80 g741691 ( .a(n_38539), .o(n_38540) );
no02f80 g757817 ( .a(n_22357), .b(n_22172), .o(n_22482) );
in01f80 g753587 ( .a(n_26670), .o(n_26671) );
no02f80 g778666 ( .a(n_45903), .b(n_1565), .o(n_2273) );
in01f80 newInst_1683 ( .a(newNet_1682), .o(newNet_1683) );
in01f80 g775259 ( .a(n_5895), .o(n_5896) );
in01f80 g744772 ( .a(n_35262), .o(n_35281) );
na02f80 g763832 ( .a(n_16612), .b(n_16464), .o(n_16648) );
in01f80 g739442 ( .a(n_40805), .o(n_40900) );
na02f80 g763416 ( .a(n_16838), .b(n_16758), .o(n_16910) );
ao12f80 g748841 ( .a(n_32441), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_19_), .o(n_33088) );
in01f80 g736891 ( .a(n_43589), .o(n_43590) );
in01f80 g774391 ( .a(n_6529), .o(n_6519) );
na02f80 g773175 ( .a(n_7817), .b(n_7908), .o(n_7919) );
in01f80 g772278 ( .a(n_8471), .o(n_8523) );
in01f80 g773198 ( .a(n_7805), .o(n_7806) );
in01f80 g770981 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_), .o(n_12061) );
na02f80 g764200 ( .a(n_16471), .b(FE_OCP_RBN2653_n_14684), .o(n_16564) );
in01f80 FE_OCPC1449_n_20443 ( .a(n_20443), .o(FE_OCPN1449_n_20443) );
no02f80 g744833 ( .a(n_34981), .b(delay_sub_ln23_0_unr22_stage8_stallmux_q), .o(n_35039) );
in01f80 newInst_57 ( .a(newNet_56), .o(newNet_57) );
in01f80 g761524 ( .a(n_18974), .o(n_20876) );
na02f80 g768112 ( .a(n_12733), .b(n_12696), .o(n_12755) );
na02f80 g781037 ( .a(cos_out_22), .b(n_43918), .o(n_347) );
in01f80 g737738 ( .a(n_42386), .o(n_42410) );
na02f80 g762930 ( .a(n_18034), .b(n_18033), .o(n_18035) );
na02f80 g743107 ( .a(n_36950), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37095) );
in01f80 newInst_2986 ( .a(newNet_2174), .o(newNet_2986) );
in01f80 g737481 ( .a(n_42637), .o(n_42650) );
oa12f80 g751428 ( .a(n_28427), .b(n_28426), .c(n_28425), .o(n_28476) );
no02f80 g776615 ( .a(n_4055), .b(n_4094), .o(n_4252) );
in01f80 g775831 ( .a(n_5516), .o(n_5583) );
no04s80 FE_RC_2520_0 ( .a(n_40942), .b(n_40963), .c(n_40941), .d(n_40824), .o(n_40979) );
na02f80 g768354 ( .a(n_12466), .b(n_12446), .o(n_12530) );
na02f80 g779600 ( .a(n_1721), .b(n_1715), .o(n_2176) );
na02f80 g771812 ( .a(FE_OCP_RBN2541_n_8800), .b(n_8562), .o(n_8849) );
in01f80 newInst_3125 ( .a(newNet_3124), .o(newNet_3125) );
in01f80 g774020 ( .a(n_7250), .o(n_7251) );
in01f80 newInst_1733 ( .a(newNet_986), .o(newNet_1733) );
in01f80 FE_OCP_RBC2917_n_10644 ( .a(n_10644), .o(FE_OCP_RBN2917_n_10644) );
na02f80 g761538 ( .a(n_18866), .b(FE_OFN778_n_17093), .o(n_18867) );
in01f80 FE_OCP_RBC3663_n_20750 ( .a(FE_OCP_RBN3662_n_20750), .o(FE_OCP_RBN3663_n_20750) );
in01f80 g752664 ( .a(n_28856), .o(n_28203) );
no02f80 g755798 ( .a(n_24320), .b(n_24319), .o(n_24321) );
no02f80 g781333 ( .a(n_1), .b(beta_7), .o(n_49) );
no02f80 g777802 ( .a(n_3238), .b(n_2504), .o(n_3252) );
in01f80 g747874 ( .a(n_32032), .o(n_32033) );
in01f80 g743742 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_11_), .o(n_36435) );
no02f80 g741626 ( .a(n_38595), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38649) );
no02f80 g749834 ( .a(n_31311), .b(n_30474), .o(n_31510) );
in01f80 g775515 ( .a(n_5348), .o(n_5349) );
in01f80 g738773 ( .a(n_41386), .o(n_41378) );
in01f80 g742089 ( .a(n_38181), .o(n_38182) );
no02f80 g762189 ( .a(n_18153), .b(n_18152), .o(n_18171) );
in01f80 newInst_2634 ( .a(newNet_2633), .o(newNet_2634) );
no02f80 g736968 ( .a(FE_OCPN1246_n_43120), .b(n_42968), .o(n_43508) );
na02f80 g761284 ( .a(n_19011), .b(FE_OCP_DRV_N1552_n_19010), .o(n_19037) );
oa22f80 g780173 ( .a(n_1093), .b(n_1203), .c(n_1094), .d(FE_OFN794_n_45813), .o(n_1163) );
no02f80 g765050 ( .a(n_15463), .b(n_15462), .o(n_15496) );
in01f80 g781289 ( .a(n_63), .o(n_64) );
in01f80 g763050 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_20_), .o(n_17416) );
no02f80 g748232 ( .a(n_31765), .b(n_31770), .o(n_31772) );
na02f80 g743908 ( .a(n_36199), .b(n_36198), .o(n_36200) );
na02f80 g758984 ( .a(n_21535), .b(n_21269), .o(n_21576) );
oa12f80 g757665 ( .a(n_22439), .b(n_22705), .c(n_22667), .o(n_22707) );
in01f80 g766207 ( .a(n_14505), .o(n_14506) );
no02f80 g746283 ( .a(n_33528), .b(FE_OCP_RBN3411_n_33547), .o(n_33644) );
in01f80 g745553 ( .a(n_34533), .o(n_34534) );
no02f80 g778569 ( .a(n_2441), .b(n_2439), .o(n_2440) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_24_ ( .ck(newNet_2843), .d(n_12131), .o(delay_add_ln22_unr8_stage4_stallmux_q_24_) );
no02f80 g755867 ( .a(n_25164), .b(n_25604), .o(n_25218) );
na02f80 FE_RC_347_0 ( .a(FE_RN_99_0), .b(FE_OCP_RBN2135_n_11780), .o(FE_RN_101_0) );
in01f80 newInst_1724 ( .a(newNet_1723), .o(newNet_1724) );
no02f80 g779556 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .o(n_1664) );
no02f80 g758919 ( .a(n_21332), .b(n_21239), .o(n_21399) );
in01f80 g741715 ( .a(n_38919), .o(n_38548) );
in01f80 FE_OCP_RBC2450_n_14114 ( .a(FE_OCP_RBN2449_n_14114), .o(FE_OCP_RBN2450_n_14114) );
in01f80 g757159 ( .a(n_23743), .o(n_23803) );
no02f80 g775553 ( .a(n_5352), .b(n_5293), .o(n_5456) );
in01f80 newInst_3597 ( .a(newNet_3596), .o(newNet_3597) );
no02f80 g753780 ( .a(n_26436), .b(n_26406), .o(n_26516) );
in01f80 g761943 ( .a(n_18431), .o(n_18594) );
in01f80 g763595 ( .a(n_17577), .o(n_17503) );
ao12f80 g780339 ( .a(n_874), .b(n_1079), .c(n_919), .o(n_967) );
in01f80 g766473 ( .a(n_14169), .o(n_14224) );
in01f80 g741932 ( .a(n_38187), .o(n_38188) );
na02f80 g759217 ( .a(n_20947), .b(n_20712), .o(n_20983) );
ao22s80 FE_RC_1344_0 ( .a(n_43613), .b(n_43832), .c(n_43614), .d(n_43831), .o(n_43861) );
in01f80 g750590 ( .a(n_31172), .o(n_30474) );
na02f80 g736880 ( .a(n_43523), .b(n_43500), .o(n_43601) );
oa22f80 FE_RC_537_0 ( .a(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .b(n_25825), .c(n_23254), .d(n_25826), .o(n_25920) );
na02f80 g758695 ( .a(n_22363), .b(n_21725), .o(n_22397) );
na02f80 g776598 ( .a(n_4218), .b(n_4092), .o(n_4385) );
in01f80 g740956 ( .a(n_39213), .o(n_39214) );
in01f80 g736443 ( .a(n_43777), .o(n_43778) );
no02f80 g750047 ( .a(n_29846), .b(n_28891), .o(n_29899) );
no02f80 g751475 ( .a(n_28568), .b(n_28577), .o(n_28601) );
in01f80 g757600 ( .a(n_22816), .o(n_22817) );
in01f80 g780305 ( .a(n_954), .o(n_1001) );
in01f80 g757971 ( .a(n_22049), .o(n_22086) );
na02f80 g771776 ( .a(FE_OCP_RBN3549_n_44575), .b(n_9157), .o(n_9158) );
no02f80 g775910 ( .a(n_5235), .b(n_4603), .o(n_5364) );
in01f80 g753650 ( .a(n_27283), .o(n_27319) );
ao12f80 g746390 ( .a(n_32947), .b(n_33458), .c(n_33021), .o(n_33506) );
no02f80 g753986 ( .a(n_26155), .b(n_23353), .o(n_26302) );
in01f80 g768177 ( .a(n_13514), .o(n_13515) );
na02f80 g746036 ( .a(n_33833), .b(n_34504), .o(n_33835) );
in01f80 g780548 ( .a(n_1111), .o(n_795) );
no02f80 g774301 ( .a(n_6806), .b(delay_xor_ln22_unr6_stage3_stallmux_q_15_), .o(n_7033) );
na02f80 g762182 ( .a(n_18153), .b(n_18152), .o(n_18202) );
oa12f80 g770384 ( .a(n_10489), .b(n_10575), .c(n_10417), .o(n_10650) );
na02f80 g740573 ( .a(n_39680), .b(n_39679), .o(n_39681) );
no02f80 g769042 ( .a(FE_OCP_RBN2119_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_9_), .o(n_11885) );
in01f80 newInst_104 ( .a(newNet_103), .o(newNet_104) );
in01f80 g750304 ( .a(n_29775), .o(n_29776) );
ms00f80 delay_xor_ln21_unr21_stage8_stallmux_q_reg_8_ ( .ck(newNet_873), .d(n_32370), .o(delay_xor_ln21_unr21_stage8_stallmux_q_8_) );
no02f80 g774083 ( .a(n_6833), .b(delay_add_ln22_unr5_stage3_stallmux_q_1_), .o(n_6834) );
in01f80 g760223 ( .a(n_20289), .o(n_20305) );
in01f80 g763931 ( .a(n_17207), .o(n_17463) );
na02f80 g756198 ( .a(n_24743), .b(n_24192), .o(n_24864) );
na02f80 g766651 ( .a(n_13860), .b(FE_OCP_RBN2249_n_13017), .o(n_13888) );
na02f80 g784416 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .o(n_46228) );
na02f80 g777996 ( .a(n_3128), .b(n_3127), .o(n_3200) );
oa12f80 g771251 ( .a(n_9783), .b(n_9782), .c(n_9781), .o(n_9878) );
in01f80 g749704 ( .a(n_31191), .o(n_31192) );
ao12f80 g780774 ( .a(n_541), .b(n_540), .c(n_539), .o(n_672) );
no02f80 g771235 ( .a(n_9686), .b(n_9615), .o(n_9817) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_19_ ( .ck(newNet_1121), .d(n_10868), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_19_) );
in01f80 g746702 ( .a(n_34774), .o(n_34299) );
na02f80 g751563 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_26_), .o(n_28722) );
oa12f80 g759663 ( .a(n_21879), .b(n_21878), .c(n_21877), .o(n_21929) );
no02f80 g751781 ( .a(n_28269), .b(n_28287), .o(n_28347) );
no02f80 g776139 ( .a(n_4611), .b(n_4639), .o(n_4784) );
na02f80 g764105 ( .a(n_16500), .b(n_16370), .o(n_16537) );
na02f80 g756741 ( .a(n_23541), .b(n_23497), .o(n_23719) );
no02f80 g746479 ( .a(n_34812), .b(n_34809), .o(n_34843) );
ao12f80 g743633 ( .a(n_37478), .b(n_37477), .c(n_46239), .o(n_37538) );
na02f80 g761909 ( .a(n_18268), .b(n_18291), .o(n_18345) );
no02f80 g775931 ( .a(n_5086), .b(n_3845), .o(n_5248) );
no02f80 FE_RC_3190_0 ( .a(FE_RN_1417_0), .b(n_17923), .o(n_18022) );
na02f80 g743523 ( .a(n_37613), .b(n_37538), .o(n_37632) );
na02f80 g737643 ( .a(n_42520), .b(n_42485), .o(n_42521) );
na02f80 g769938 ( .a(n_11003), .b(n_11013), .o(n_11091) );
no02f80 g753224 ( .a(n_27204), .b(FE_OCP_RBN2833_n_26081), .o(n_27384) );
in01f80 g773545 ( .a(n_7445), .o(n_7446) );
na02f80 g758269 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_22_), .o(n_22879) );
no02f80 g746973 ( .a(FE_OCP_RBN2167_n_32892), .b(n_32540), .o(n_33063) );
na02f80 g775283 ( .a(FE_OCP_RBN2980_n_5656), .b(n_4759), .o(n_5713) );
na02f80 g775579 ( .a(n_5309), .b(n_4759), .o(n_5581) );
na02f80 g746597 ( .a(n_34612), .b(n_34667), .o(n_34740) );
oa22f80 g766146 ( .a(n_14590), .b(FE_OCP_RBN2505_n_13896), .c(FE_OCP_RBN2627_n_14590), .d(FE_OCP_RBN2503_n_13896), .o(n_14704) );
no02f80 g768076 ( .a(n_12790), .b(n_12134), .o(n_12855) );
in01f80 g736833 ( .a(n_43064), .o(n_43065) );
in01f80 g743430 ( .a(n_36657), .o(n_36631) );
in01f80 FE_OCP_RBC2320_n_2382 ( .a(n_2382), .o(FE_OCP_RBN2320_n_2382) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_19_ ( .ck(newNet_2199), .d(n_1132), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_13_ ( .ck(newNet_3075), .d(n_1169), .o(delay_add_ln22_unr2_stage2_stallmux_q_13_) );
no02f80 g773502 ( .a(n_7488), .b(n_7295), .o(n_7497) );
in01f80 g746535 ( .a(n_34806), .o(n_34807) );
oa22f80 g776542 ( .a(n_47012), .b(n_4182), .c(n_4289), .d(n_4046), .o(n_4378) );
no02f80 g767500 ( .a(n_13265), .b(FE_OCP_DRV_N3152_n_13264), .o(n_13357) );
in01f80 g741928 ( .a(n_38820), .o(n_38144) );
in01f80 FE_OCP_DRV_C3152_n_13264 ( .a(FE_OCP_DRV_N3151_n_13264), .o(FE_OCP_DRV_N3152_n_13264) );
no02f80 FE_RC_2158_0 ( .a(n_14452), .b(FE_OCP_RBN3657_n_15314), .o(FE_RN_764_0) );
in01f80 g751768 ( .a(n_28329), .o(n_28330) );
in01f80 g748938 ( .a(n_31035), .o(n_31036) );
na02f80 g769561 ( .a(n_11416), .b(n_11374), .o(n_11503) );
na02f80 g771627 ( .a(n_9027), .b(n_8862), .o(n_9076) );
in01f80 FE_RC_1518_0 ( .a(FE_RN_428_0), .o(n_32224) );
oa12f80 g754205 ( .a(n_26910), .b(n_26909), .c(n_26908), .o(n_26973) );
in01f80 g740049 ( .a(n_40078), .o(n_40079) );
in01f80 FE_OCP_RBC2328_n_29378 ( .a(FE_OCP_RBN2327_n_29378), .o(FE_OCP_RBN2328_n_29378) );
in01f80 FE_OCP_RBC3595_n_14785 ( .a(n_14785), .o(FE_OCP_RBN3595_n_14785) );
in01f80 g773358 ( .a(n_7743), .o(n_7886) );
no02f80 FE_RC_1737_0 ( .a(FE_RN_484_0), .b(n_37245), .o(n_37291) );
na02f80 g754921 ( .a(n_25327), .b(n_25386), .o(n_25760) );
no02f80 g755163 ( .a(n_25373), .b(n_24570), .o(n_25647) );
in01f80 g747342 ( .a(n_32682), .o(n_32683) );
no02f80 g740760 ( .a(n_39532), .b(n_39072), .o(n_39533) );
oa12f80 g779107 ( .a(n_1794), .b(n_1958), .c(n_1619), .o(n_1974) );
in01f80 newInst_3102 ( .a(newNet_3101), .o(newNet_3102) );
in01f80 FE_RC_4072_0 ( .a(FE_RN_1774_0), .o(FE_RN_1773_0) );
ao12f80 g767094 ( .a(n_13412), .b(n_13413), .c(FE_OCP_DRV_N1536_n_12633), .o(n_13460) );
oa12f80 g737294 ( .a(n_42512), .b(n_42860), .c(n_42462), .o(n_42886) );
na02f80 g773247 ( .a(n_7624), .b(n_7623), .o(n_7625) );
in01f80 FE_OCP_RBC1909_n_20545 ( .a(n_20545), .o(FE_OCP_RBN1909_n_20545) );
in01f80 newInst_2060 ( .a(newNet_935), .o(newNet_2060) );
na02f80 g773522 ( .a(n_7468), .b(n_7467), .o(n_8302) );
na02f80 g758074 ( .a(n_22466), .b(n_22465), .o(n_22504) );
oa12f80 g736366 ( .a(n_43521), .b(n_43772), .c(n_43255), .o(n_43807) );
in01f80 g771717 ( .a(n_8865), .o(n_8908) );
in01f80 g753420 ( .a(n_27021), .o(n_27022) );
oa12f80 g755385 ( .a(n_25495), .b(n_25494), .c(n_25493), .o(n_25683) );
na02f80 g759639 ( .a(n_20723), .b(n_44160), .o(n_20724) );
no02f80 g780695 ( .a(n_647), .b(n_643), .o(n_644) );
in01f80 FE_OCP_RBC1346_n_19270 ( .a(n_19270), .o(FE_OCP_RBN1346_n_19270) );
oa22f80 g776149 ( .a(n_4782), .b(n_3993), .c(n_4783), .d(n_4017), .o(n_4989) );
na02f80 g775513 ( .a(n_5759), .b(FE_OCP_RBN2817_n_4458), .o(n_5842) );
na02f80 g760399 ( .a(n_20141), .b(FE_OCP_RBN1331_n_18866), .o(n_20190) );
na02f80 g742417 ( .a(FE_OCP_RBN2210_n_37694), .b(n_37054), .o(n_37722) );
in01f80 g771916 ( .a(n_9035), .o(n_9064) );
no02f80 FE_RC_3513_0 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_8_), .b(n_28273), .o(FE_RN_1517_0) );
in01f80 FE_RC_1931_0 ( .a(n_18741), .o(FE_RN_613_0) );
in01f80 newInst_2234 ( .a(newNet_2233), .o(newNet_2234) );
no02f80 g738364 ( .a(n_41549), .b(n_41514), .o(n_41594) );
no02f80 FE_RC_1935_0 ( .a(FE_RN_615_0), .b(n_19246), .o(FE_RN_616_0) );
in01f80 g745177 ( .a(n_34706), .o(n_36091) );
na02f80 g771283 ( .a(n_9447), .b(n_9464), .o(n_9615) );
na02f80 g750610 ( .a(n_29421), .b(FE_OCPN1752_n_29420), .o(n_29444) );
no02f80 g739320 ( .a(n_40670), .b(n_40699), .o(n_40740) );
oa22f80 g778967 ( .a(n_2103), .b(n_1901), .c(FE_OCP_RBN2196_n_2103), .d(n_1902), .o(n_2929) );
in01f80 g752290 ( .a(n_27895), .o(n_27896) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_11_ ( .ck(newNet_2977), .d(n_5645), .o(delay_add_ln22_unr5_stage3_stallmux_q_11_) );
no02f80 g754086 ( .a(n_25972), .b(n_26057), .o(n_26102) );
in01f80 newInst_3540 ( .a(newNet_3539), .o(newNet_3540) );
oa12f80 g759018 ( .a(n_21355), .b(n_21354), .c(n_21353), .o(n_21426) );
na02f80 g769728 ( .a(n_11254), .b(n_11253), .o(n_11345) );
na02f80 g737761 ( .a(n_42307), .b(n_42323), .o(n_42308) );
no02f80 g771549 ( .a(n_8881), .b(n_8913), .o(n_8977) );
na02f80 g738374 ( .a(n_41697), .b(FE_OCP_RBN2311_n_41420), .o(n_41746) );
oa22f80 g747676 ( .a(n_32061), .b(n_31894), .c(n_32062), .d(n_31893), .o(n_32147) );
na02f80 g745605 ( .a(n_34315), .b(FE_OCP_RBN1684_n_33491), .o(n_34381) );
no02f80 g741814 ( .a(n_38391), .b(n_38390), .o(n_38392) );
na02f80 g753229 ( .a(n_27204), .b(n_26146), .o(n_27338) );
in01f80 g754430 ( .a(n_25729), .o(n_25728) );
in01f80 newInst_2598 ( .a(newNet_2597), .o(newNet_2598) );
in01f80 FE_RC_1979_0 ( .a(n_19799), .o(FE_RN_643_0) );
no02f80 g761722 ( .a(n_18439), .b(n_18311), .o(n_18602) );
na02f80 g777853 ( .a(n_3356), .b(n_3310), .o(n_3363) );
na02f80 g752583 ( .a(n_45766), .b(n_27433), .o(n_27634) );
in01f80 newInst_1936 ( .a(newNet_927), .o(newNet_1936) );
na02f80 FE_RC_2671_0 ( .a(FE_RN_1116_0), .b(FE_RN_1117_0), .o(n_3890) );
na02f80 g769132 ( .a(n_11678), .b(n_11624), .o(n_11799) );
in01f80 g766302 ( .a(n_45521), .o(n_14439) );
no02f80 g776291 ( .a(FE_OCP_RBN3665_n_4604), .b(n_5529), .o(n_4713) );
in01f80 g761297 ( .a(n_19033), .o(n_20307) );
no02f80 g767079 ( .a(n_13791), .b(n_13790), .o(n_13792) );
oa22f80 g784546 ( .a(n_11453), .b(FE_OFN801_n_46285), .c(n_11422), .d(FE_OCP_RBN3044_n_46337), .o(n_46367) );
in01f80 g759706 ( .a(n_20680), .o(n_20681) );
oa12f80 g778242 ( .a(n_2111), .b(n_2615), .c(n_2153), .o(n_2699) );
no02f80 g746254 ( .a(n_33592), .b(n_33618), .o(n_33711) );
na02f80 g744462 ( .a(n_35470), .b(n_35469), .o(n_35484) );
ms00f80 delay_sub_ln22_unr24_stage9_stallmux_q_reg_2_ ( .ck(newNet_1908), .d(n_36782), .o(delay_sub_ln22_unr24_stage9_stallmux_q_2_) );
in01f80 g759187 ( .a(n_21159), .o(n_21160) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_3_ ( .ck(newNet_2356), .d(n_35426), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_3_) );
in01f80 newInst_2217 ( .a(newNet_2216), .o(newNet_2217) );
na02f80 g737777 ( .a(n_42328), .b(n_42327), .o(n_42348) );
na02f80 g766378 ( .a(FE_OCP_RBN2455_n_14157), .b(n_14274), .o(n_14277) );
in01f80 g770412 ( .a(n_10535), .o(n_10536) );
no02f80 g748180 ( .a(n_31967), .b(n_32046), .o(n_32126) );
in01f80 g767537 ( .a(n_14742), .o(n_14869) );
na02f80 g766021 ( .a(FE_OCP_RBN1183_n_14638), .b(FE_OCP_RBN3535_n_13765), .o(n_14695) );
na02f80 g751358 ( .a(n_29432), .b(n_29431), .o(n_29433) );
in01f80 newInst_746 ( .a(newNet_745), .o(newNet_746) );
no02f80 g753537 ( .a(n_26759), .b(n_26730), .o(n_26851) );
na02f80 g775859 ( .a(n_5262), .b(n_5261), .o(n_5263) );
na02f80 g759926 ( .a(n_21051), .b(n_21244), .o(n_21335) );
no02f80 g747114 ( .a(n_32890), .b(n_32907), .o(n_32990) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_15_ ( .ck(newNet_841), .d(n_1332), .o(delay_xor_ln21_unr3_stage2_stallmux_q_15_) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_1_ ( .ck(newNet_2658), .d(n_20970), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_1_) );
oa12f80 g756424 ( .a(n_23588), .b(n_23615), .c(n_23587), .o(n_23668) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_8_ ( .ck(newNet_1677), .d(n_21994), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_8_) );
na02f80 g766257 ( .a(n_14247), .b(n_14288), .o(n_14412) );
no02f80 g754411 ( .a(FE_OCP_RBN3630_n_25656), .b(FE_OCP_DRV_N3743_n_25400), .o(n_25707) );
no02f80 g766062 ( .a(n_14629), .b(n_47256), .o(n_14801) );
na02f80 g762302 ( .a(n_18094), .b(n_18110), .o(n_18161) );
na02f80 g781244 ( .a(n_102), .b(n_101), .o(n_149) );
na02f80 g767834 ( .a(n_12999), .b(n_12919), .o(n_13208) );
na02f80 g762202 ( .a(n_18624), .b(n_18623), .o(n_18625) );
in01f80 FE_OCP_RBC2558_n_44576 ( .a(FE_OCP_RBN2557_n_44576), .o(FE_OCP_RBN2558_n_44576) );
in01f80 g764720 ( .a(n_15802), .o(n_15803) );
na02f80 g748040 ( .a(n_32107), .b(n_31969), .o(n_32106) );
in01f80 newInst_1477 ( .a(newNet_1476), .o(newNet_1477) );
na02f80 FE_RC_2232_0 ( .a(FE_RN_812_0), .b(n_17499), .o(FE_RN_813_0) );
no02f80 g750819 ( .a(n_29188), .b(n_29187), .o(n_29190) );
no02f80 g749960 ( .a(n_29810), .b(n_29795), .o(n_29834) );
ao12f80 g780803 ( .a(n_491), .b(n_481), .c(n_509), .o(n_510) );
na02f80 g755629 ( .a(n_24614), .b(n_24613), .o(n_24713) );
na02f80 g754266 ( .a(n_25847), .b(n_23254), .o(n_25881) );
na02f80 g760171 ( .a(n_20334), .b(n_20399), .o(n_20460) );
na02f80 g742848 ( .a(n_37270), .b(n_37252), .o(n_37276) );
na02f80 g745613 ( .a(n_34369), .b(FE_OCP_RBN3433_n_33664), .o(n_34509) );
no02f80 g759201 ( .a(n_21309), .b(n_21268), .o(n_21461) );
na02f80 g737490 ( .a(n_42555), .b(n_42215), .o(n_42603) );
no02f80 g776036 ( .a(n_5077), .b(n_4428), .o(n_5181) );
na02f80 g772732 ( .a(n_8227), .b(n_8226), .o(n_8263) );
no02f80 g748217 ( .a(n_32780), .b(n_32501), .o(n_32778) );
in01f80 g742579 ( .a(n_37493), .o(n_38290) );
in01f80 FE_OCP_RBC2697_n_14814 ( .a(FE_OCP_RBN2696_n_14814), .o(FE_OCP_RBN2697_n_14814) );
in01f80 g778699 ( .a(n_2652), .o(n_2589) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_10_ ( .ck(newNet_3087), .d(n_1134), .o(delay_add_ln22_unr2_stage2_stallmux_q_10_) );
oa22f80 g744106 ( .a(n_36870), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_1_), .c(n_36871), .d(n_36898), .o(n_36915) );
na02f80 g776850 ( .a(n_4172), .b(n_4171), .o(n_4267) );
no02f80 g768736 ( .a(n_45659), .b(delay_xor_ln21_unr9_stage4_stallmux_q_14_), .o(n_12148) );
in01f80 g739889 ( .a(n_40400), .o(n_40401) );
no02f80 g760056 ( .a(n_20409), .b(n_20406), .o(n_20465) );
no02f80 g739282 ( .a(n_40775), .b(n_40774), .o(n_40776) );
in01f80 FE_RC_520_0 ( .a(n_23772), .o(FE_RN_163_0) );
na02f80 g753079 ( .a(n_27506), .b(n_27421), .o(n_27528) );
no02f80 g763942 ( .a(n_16570), .b(n_16533), .o(n_16611) );
in01f80 newInst_3379 ( .a(newNet_272), .o(newNet_3379) );
in01f80 FE_RC_2830_0 ( .a(n_23761), .o(FE_RN_1216_0) );
no02f80 g756812 ( .a(n_23377), .b(n_23376), .o(n_23394) );
oa22f80 g784532 ( .a(n_12145), .b(FE_OFN803_n_46285), .c(n_12102), .d(FE_OFN771_n_46337), .o(n_46353) );
in01f80 g751724 ( .a(n_30038), .o(n_30104) );
no02f80 g743350 ( .a(n_36660), .b(n_36635), .o(n_36693) );
in01f80 FE_OCP_RBC1987_delay_xor_ln23_unr6_stage3_stallmux_q ( .a(delay_xor_ln23_unr6_stage3_stallmux_q), .o(FE_OCP_RBN1987_delay_xor_ln23_unr6_stage3_stallmux_q) );
oa12f80 g746528 ( .a(FE_OCP_RBN2601_n_34388), .b(n_34615), .c(n_34614), .o(n_34642) );
na02f80 g739666 ( .a(n_40535), .b(n_40224), .o(n_40556) );
na02f80 g738291 ( .a(n_41888), .b(n_41550), .o(n_41776) );
in01f80 g759626 ( .a(n_20690), .o(n_20647) );
na02f80 g755492 ( .a(n_24777), .b(n_24822), .o(n_24883) );
in01f80 FE_RC_2064_0 ( .a(n_35078), .o(FE_RN_701_0) );
in01f80 g767300 ( .a(n_13714), .o(n_13715) );
na02f80 g752795 ( .a(n_27813), .b(n_27453), .o(n_27814) );
oa12f80 g781133 ( .a(n_116), .b(n_215), .c(n_82), .o(n_219) );
in01f80 g774421 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_0_), .o(n_6510) );
ao12f80 g761514 ( .a(n_19000), .b(n_18999), .c(n_18998), .o(n_20852) );
in01f80 g775432 ( .a(n_5436), .o(n_5437) );
na02f80 g736724 ( .a(n_43138), .b(n_43228), .o(n_43229) );
in01f80 g748527 ( .a(n_31713), .o(n_31714) );
no02f80 g763601 ( .a(n_16713), .b(n_16735), .o(n_16764) );
na02f80 g769774 ( .a(n_11144), .b(n_11134), .o(n_11198) );
in01f80 g780915 ( .a(n_411), .o(n_434) );
na02f80 FE_RC_2067_0 ( .a(n_30504), .b(FE_RN_702_0), .o(FE_RN_703_0) );
no02f80 g749957 ( .a(n_30443), .b(n_30422), .o(n_30482) );
in01f80 newInst_1705 ( .a(newNet_265), .o(newNet_1705) );
in01f80 newInst_1519 ( .a(newNet_1518), .o(newNet_1519) );
no02f80 g758169 ( .a(n_44268), .b(FE_OCP_RBN1915_n_20965), .o(n_22308) );
no02f80 g761480 ( .a(n_19649), .b(n_19825), .o(n_20178) );
na02f80 g760242 ( .a(FE_OCP_RBN3617_n_20249), .b(n_19340), .o(n_20458) );
ao12f80 g747704 ( .a(n_33571), .b(n_33653), .c(n_33720), .o(n_33654) );
ao12f80 g764593 ( .a(n_16025), .b(n_16448), .c(n_15821), .o(n_16573) );
na02f80 g746548 ( .a(n_34420), .b(n_34419), .o(n_34421) );
in01f80 FE_OCPC1406_n_25859 ( .a(FE_OCPN1405_n_25859), .o(FE_OCPN1406_n_25859) );
na02f80 g761205 ( .a(n_19080), .b(n_18596), .o(n_19105) );
no03m80 g738974 ( .a(n_41206), .b(n_41193), .c(n_40812), .o(n_41280) );
na02f80 FE_RC_2625_0 ( .a(n_28342), .b(n_28343), .o(FE_RN_1093_0) );
in01f80 g754353 ( .a(n_25874), .o(n_25890) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_0_ ( .ck(newNet_1267), .d(n_151), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_) );
in01f80 g753181 ( .a(n_27124), .o(n_27232) );
in01f80 g762211 ( .a(n_18771), .o(n_18772) );
in01f80 g745598 ( .a(n_34374), .o(n_34852) );
na02f80 g760573 ( .a(n_19862), .b(n_19839), .o(n_19863) );
in01f80 g763310 ( .a(n_17005), .o(n_17006) );
in01f80 g743401 ( .a(n_36730), .o(n_36731) );
oa12f80 g763222 ( .a(n_16869), .b(n_17001), .c(n_16951), .o(n_17091) );
in01f80 g753247 ( .a(n_27454), .o(n_27455) );
no02f80 g769371 ( .a(n_45685), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .o(n_12079) );
in01f80 g737954 ( .a(n_42339), .o(n_42340) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_17_ ( .ck(newNet_1126), .d(n_10815), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_17_) );
no02f80 g755622 ( .a(n_24518), .b(FE_OCPN1474_n_24624), .o(n_24564) );
in01f80 newInst_1552 ( .a(newNet_1551), .o(newNet_1552) );
ao22s80 g774235 ( .a(n_6580), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .d(delay_xor_ln22_unr6_stage3_stallmux_q_6_), .o(n_6609) );
in01f80 g745192 ( .a(n_34493), .o(n_34542) );
no02f80 g740166 ( .a(n_39816), .b(n_39917), .o(n_40042) );
na02f80 FE_RC_1898_0 ( .a(FE_RN_593_0), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24359) );
na02f80 g743675 ( .a(n_36411), .b(n_36013), .o(n_36427) );
no02f80 FE_RC_2411_0 ( .a(FE_RN_950_0), .b(n_2318), .o(FE_RN_951_0) );
na02f80 g768260 ( .a(n_12591), .b(n_12587), .o(n_12588) );
oa22f80 FE_RC_1624_0 ( .a(n_32187), .b(n_32211), .c(n_32210), .d(n_32186), .o(n_32259) );
in01f80 newInst_2053 ( .a(newNet_2052), .o(newNet_2053) );
oa12f80 g745694 ( .a(n_35436), .b(n_35435), .c(n_35434), .o(n_35840) );
oa22f80 g763434 ( .a(n_46975), .b(FE_OFN767_n_15670), .c(n_16895), .d(n_17753), .o(n_17029) );
no02f80 g766065 ( .a(n_14704), .b(FE_OCP_RBN2506_n_13896), .o(n_14782) );
na02f80 g749294 ( .a(n_30611), .b(n_30537), .o(n_30630) );
in01f80 g756491 ( .a(n_23716), .o(n_23717) );
no02f80 g780811 ( .a(n_504), .b(n_420), .o(n_536) );
in01f80 g777877 ( .a(n_3228), .o(n_3186) );
oa22f80 g779898 ( .a(n_44652), .b(n_1099), .c(n_44661), .d(n_1098), .o(n_1294) );
no02f80 g770697 ( .a(n_9861), .b(n_9111), .o(n_9946) );
na02f80 g745737 ( .a(n_34177), .b(n_34203), .o(n_34204) );
no02f80 g750173 ( .a(n_30898), .b(n_30897), .o(n_30899) );
ao12f80 g759690 ( .a(n_20309), .b(n_20476), .c(n_20311), .o(n_20616) );
oa12f80 g760059 ( .a(FE_OCP_RBN3845_FE_RN_1242_0), .b(FE_OCP_RBN3850_n_20290), .c(n_20125), .o(n_20344) );
in01f80 FE_RC_2253_0 ( .a(FE_RN_831_0), .o(n_18104) );
na02f80 g780392 ( .a(n_785), .b(n_745), .o(n_848) );
na02f80 g738432 ( .a(n_41506), .b(n_41541), .o(n_41593) );
in01f80 newInst_3633 ( .a(newNet_3632), .o(newNet_3633) );
na02f80 g745389 ( .a(n_36049), .b(n_35629), .o(n_36117) );
na02f80 g736780 ( .a(n_43305), .b(n_43350), .o(n_43396) );
na02f80 g766031 ( .a(n_14664), .b(n_14639), .o(n_14665) );
ao22s80 FE_RC_419_0 ( .a(FE_OCP_RBN3535_n_13765), .b(FE_OCP_RBN2590_n_14460), .c(n_14460), .d(FE_OCP_RBN3528_n_13765), .o(n_14591) );
in01f80 g775592 ( .a(n_5725), .o(n_5726) );
in01f80 g775088 ( .a(n_6086), .o(n_6094) );
na02f80 g751181 ( .a(n_29944), .b(n_29940), .o(n_30028) );
na02f80 g770032 ( .a(n_10852), .b(n_44464), .o(n_10877) );
no02f80 g740851 ( .a(n_39348), .b(n_39255), .o(n_39493) );
no02f80 FE_RC_3534_0 ( .a(FE_OCP_RBN3212_n_44365), .b(FE_RN_1528_0), .o(FE_RN_1529_0) );
na02f80 g762309 ( .a(n_18074), .b(n_17945), .o(n_18110) );
no02f80 g767377 ( .a(n_13398), .b(n_12436), .o(n_13480) );
ao12f80 g784695 ( .a(n_2605), .b(n_2604), .c(n_3039), .o(n_47025) );
in01f80 g751262 ( .a(FE_OCP_DRV_N1576_n_28829), .o(n_29866) );
ao12f80 g749614 ( .a(n_30383), .b(FE_OCP_RBN1357_n_30298), .c(n_30423), .o(n_30448) );
in01f80 g756759 ( .a(n_23539), .o(n_23540) );
no02f80 FE_RC_712_0 ( .a(FE_RN_227_0), .b(n_23194), .o(n_47337) );
in01f80 g737410 ( .a(n_43129), .o(n_42804) );
no02f80 g741947 ( .a(n_37991), .b(n_37989), .o(n_37990) );
na02f80 g762272 ( .a(n_18727), .b(n_18665), .o(n_19523) );
ao12f80 g746019 ( .a(n_33879), .b(n_33878), .c(n_33877), .o(n_35382) );
in01f80 g774812 ( .a(n_6368), .o(n_6369) );
in01f80 FE_RC_2691_0 ( .a(n_3862), .o(FE_RN_1127_0) );
oa22f80 g777217 ( .a(n_3637), .b(n_5109), .c(n_3690), .d(n_3381), .o(n_3929) );
ao12f80 g768816 ( .a(n_11685), .b(n_11850), .c(n_11597), .o(n_11952) );
in01f80 g755523 ( .a(n_25224), .o(n_25261) );
na02f80 g740833 ( .a(n_39239), .b(n_39058), .o(n_39292) );
in01f80 FE_OCPC1001_n_45660 ( .a(FE_OCPN1000_n_45660), .o(FE_OCPN1001_n_45660) );
in01f80 g753494 ( .a(n_26954), .o(n_26955) );
na02f80 g776327 ( .a(n_4762), .b(n_4761), .o(n_4823) );
in01f80 FE_OCP_RBC1726_n_20924 ( .a(n_20924), .o(FE_OCP_RBN1726_n_20924) );
na02f80 g769417 ( .a(n_11354), .b(n_11393), .o(n_11453) );
no02f80 g740642 ( .a(n_39526), .b(n_39498), .o(n_39577) );
in01f80 g757799 ( .a(n_22622), .o(n_22701) );
in01f80 g776750 ( .a(n_4009), .o(n_4069) );
no02f80 g775716 ( .a(FE_OCP_RBN2929_n_5221), .b(FE_OCPN846_n_4046), .o(n_5306) );
na02f80 g771607 ( .a(n_10210), .b(n_10209), .o(n_10211) );
no02f80 g751062 ( .a(n_30303), .b(n_30165), .o(n_30438) );
in01f80 g752100 ( .a(n_28793), .o(n_28897) );
no02f80 g754684 ( .a(FE_OCP_RBN2966_n_26231), .b(n_26680), .o(n_26860) );
in01f80 FE_RC_1423_0 ( .a(n_22351), .o(FE_RN_414_0) );
in01f80 g756592 ( .a(n_23874), .o(n_23875) );
no02f80 g781312 ( .a(beta_31), .b(beta_10), .o(n_60) );
na02f80 g770769 ( .a(n_10115), .b(n_10093), .o(n_10355) );
oa22f80 g741759 ( .a(n_38425), .b(n_38036), .c(FE_OCP_RBN3445_n_37945), .d(n_37639), .o(n_38478) );
no03m80 g738316 ( .a(n_41574), .b(n_41757), .c(n_41440), .o(n_41836) );
no02f80 FE_RC_2354_0 ( .a(FE_RN_904_0), .b(FE_RN_906_0), .o(FE_RN_907_0) );
in01f80 g749849 ( .a(n_31114), .o(n_31115) );
no02f80 g742836 ( .a(n_37200), .b(n_36989), .o(n_37223) );
no02f80 g771521 ( .a(n_8985), .b(FE_OCP_RBN2468_n_8767), .o(n_8986) );
no02f80 g778002 ( .a(n_3103), .b(n_3140), .o(n_3172) );
in01f80 g751891 ( .a(n_28838), .o(n_28839) );
in01f80 g746803 ( .a(n_33404), .o(n_33405) );
na02f80 g755038 ( .a(n_25323), .b(n_25206), .o(n_25628) );
no02f80 g769620 ( .a(n_11302), .b(n_11315), .o(n_11370) );
in01f80 g745209 ( .a(n_35521), .o(n_34628) );
no02f80 g766731 ( .a(n_13750), .b(FE_OCP_RBN2243_n_13017), .o(n_13808) );
in01f80 g765609 ( .a(n_15156), .o(n_15135) );
in01f80 newInst_3513 ( .a(newNet_3512), .o(newNet_3513) );
no02f80 g766073 ( .a(n_14641), .b(n_13487), .o(n_14662) );
no02f80 g742916 ( .a(n_36976), .b(n_37012), .o(n_37402) );
oa22f80 g744557 ( .a(n_36639), .b(n_36213), .c(n_36638), .d(n_36214), .o(n_36699) );
no02f80 g771985 ( .a(FE_OFN754_n_44461), .b(n_9369), .o(n_9596) );
na02f80 g760695 ( .a(n_19601), .b(n_19645), .o(n_19646) );
oa12f80 g768275 ( .a(n_12562), .b(n_12561), .c(n_12560), .o(n_12605) );
in01f80 g754344 ( .a(n_25893), .o(n_25909) );
no02f80 g758891 ( .a(n_21362), .b(n_45073), .o(n_21507) );
in01f80 newInst_508 ( .a(newNet_306), .o(newNet_508) );
oa22f80 FE_RC_1392_0 ( .a(n_11743), .b(n_11980), .c(n_11744), .d(n_44857), .o(n_12162) );
in01f80 FE_OCP_RBC2937_n_16113 ( .a(n_16113), .o(FE_OCP_RBN2937_n_16113) );
na02f80 g750637 ( .a(FE_OCP_RBN2331_n_29353), .b(n_28850), .o(n_29352) );
na02f80 g749644 ( .a(FE_OCP_RBN3708_n_31396), .b(n_31640), .o(n_31642) );
na02f80 g744241 ( .a(n_46228), .b(n_36855), .o(n_37958) );
no02f80 g769210 ( .a(n_11607), .b(n_11606), .o(n_11680) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_4_ ( .ck(newNet_3110), .d(n_39986), .o(delay_add_ln22_unr27_stage10_stallmux_q_4_) );
na02f80 g770418 ( .a(n_10369), .b(FE_OCP_RBN3637_n_44490), .o(n_10408) );
na02f80 g740116 ( .a(n_40188), .b(n_40106), .o(n_40223) );
no02f80 g778371 ( .a(n_2685), .b(n_1031), .o(n_2797) );
no02f80 g738741 ( .a(n_41483), .b(n_41481), .o(n_41527) );
in01f80 g741616 ( .a(n_38615), .o(n_38627) );
in01f80 g775999 ( .a(n_4959), .o(n_4960) );
oa12f80 g775598 ( .a(n_4788), .b(n_5552), .c(n_5548), .o(n_5553) );
in01f80 g766078 ( .a(n_14611), .o(n_14639) );
na02f80 g764482 ( .a(FE_OCP_RBN2937_n_16113), .b(n_16036), .o(n_16189) );
in01f80 newInst_1086 ( .a(newNet_1085), .o(newNet_1086) );
oa12f80 g773750 ( .a(n_7223), .b(n_7222), .c(n_7221), .o(n_7321) );
ao12f80 g765028 ( .a(n_14987), .b(n_15084), .c(n_14986), .o(n_15242) );
no02f80 g775441 ( .a(FE_OCP_RBN2973_n_5531), .b(n_4875), .o(n_5576) );
no02f80 g773679 ( .a(n_7269), .b(n_7291), .o(n_7318) );
oa22f80 FE_RC_1211_0 ( .a(n_12936), .b(n_13758), .c(n_12935), .d(n_13757), .o(n_13858) );
oa22f80 g764138 ( .a(n_16817), .b(n_16304), .c(n_16816), .d(n_16305), .o(n_16925) );
in01f80 newInst_1776 ( .a(newNet_1775), .o(newNet_1776) );
in01f80 g749677 ( .a(n_30149), .o(n_30150) );
na02f80 g762396 ( .a(n_45118), .b(n_17882), .o(n_18620) );
ao12f80 g780189 ( .a(n_796), .b(n_1069), .c(n_762), .o(n_1090) );
oa12f80 g742618 ( .a(n_37404), .b(n_37403), .c(n_37402), .o(n_37929) );
no02f80 g775169 ( .a(n_5881), .b(n_4556), .o(n_5943) );
no02f80 g745715 ( .a(n_34129), .b(n_44100), .o(n_34166) );
na02f80 g753174 ( .a(n_27070), .b(n_25595), .o(n_27126) );
in01f80 FE_OCP_RBC2954_n_26231 ( .a(n_26231), .o(FE_OCP_RBN2954_n_26231) );
in01f80 g766137 ( .a(n_14736), .o(n_14737) );
in01f80 g743960 ( .a(n_35828), .o(n_35829) );
in01f80 g748778 ( .a(n_32539), .o(n_32460) );
na02f80 g771567 ( .a(n_9079), .b(n_9115), .o(n_9305) );
na02f80 FE_RC_3929_0 ( .a(FE_RN_1699_0), .b(n_32578), .o(n_32520) );
ao12f80 g748511 ( .a(n_31332), .b(n_31426), .c(n_31382), .o(n_31447) );
in01f80 g766699 ( .a(n_46984), .o(n_14013) );
in01f80 newInst_2895 ( .a(newNet_2894), .o(newNet_2895) );
no02f80 g780026 ( .a(n_1255), .b(n_978), .o(n_1258) );
no03m80 g742466 ( .a(n_37602), .b(FE_OCP_RBN2183_FE_RN_464_0), .c(n_37567), .o(n_37666) );
ao12f80 g752523 ( .a(n_27388), .b(n_27634), .c(n_27425), .o(n_27703) );
no02f80 g763239 ( .a(FE_OCP_RBN3214_n_44365), .b(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .o(n_17339) );
no04s80 g743590 ( .a(n_46217), .b(n_46200), .c(n_37586), .d(n_46218), .o(n_37611) );
no02f80 g738732 ( .a(n_41483), .b(n_41482), .o(n_41532) );
in01f80 FE_RC_3015_0 ( .a(n_35057), .o(FE_RN_1322_0) );
in01f80 g781080 ( .a(n_262), .o(n_273) );
na02f80 g760998 ( .a(n_19321), .b(n_19351), .o(n_19445) );
in01f80 g745723 ( .a(n_35842), .o(n_35476) );
in01f80 FE_OFC349_n_8981 ( .a(FE_OFN790_n_8981), .o(FE_OFN349_n_8981) );
na02f80 g769639 ( .a(n_11294), .b(n_11260), .o(n_11346) );
in01f80 g770686 ( .a(n_10020), .o(n_10065) );
oa22f80 g752640 ( .a(n_27533), .b(n_27529), .c(n_27532), .d(n_27528), .o(n_27580) );
na02f80 g760154 ( .a(n_20537), .b(FE_OCP_RBN3521_n_19663), .o(n_20752) );
na02f80 g747279 ( .a(n_45753), .b(n_33885), .o(n_33887) );
ao22s80 FE_RC_3726_0 ( .a(n_14464), .b(FE_OCP_RBN2630_n_14912), .c(n_14465), .d(n_14912), .o(n_15021) );
na02f80 g771289 ( .a(n_9785), .b(n_9784), .o(n_9836) );
no02f80 FE_RC_1426_0 ( .a(FE_RN_415_0), .b(FE_RN_414_0), .o(FE_RN_416_0) );
in01f80 g775020 ( .a(n_6154), .o(n_6124) );
oa12f80 g738128 ( .a(n_42080), .b(n_42079), .c(n_42078), .o(n_42421) );
in01f80 newInst_2470 ( .a(newNet_1969), .o(newNet_2470) );
oa12f80 g748738 ( .a(n_31355), .b(n_31354), .c(n_31353), .o(n_31397) );
in01f80 FE_RC_1553_0 ( .a(FE_OCP_RBN2301_n_7817), .o(FE_RN_438_0) );
no02f80 g749025 ( .a(n_30961), .b(n_31025), .o(n_31032) );
in01f80 g754119 ( .a(n_26112), .o(n_26142) );
oa12f80 g781004 ( .a(n_87), .b(n_273), .c(n_100), .o(n_279) );
ao12f80 g755313 ( .a(n_24882), .b(n_24920), .c(n_24919), .o(n_24976) );
na02f80 g738468 ( .a(n_41387), .b(n_41153), .o(n_41470) );
na02f80 FE_RC_143_0 ( .a(n_18006), .b(FE_RN_40_0), .o(FE_RN_41_0) );
in01f80 g750511 ( .a(n_29525), .o(n_29526) );
in01f80 g766178 ( .a(n_14545), .o(n_14546) );
in01f80 FE_OFC747_n_13889 ( .a(FE_OCP_RBN2200_n_13889), .o(FE_OFN747_n_13889) );
oa22f80 g768103 ( .a(n_12602), .b(n_12494), .c(n_12603), .d(n_12493), .o(n_13163) );
na02f80 g759589 ( .a(n_20422), .b(n_20413), .o(n_20447) );
in01f80 g760597 ( .a(n_19817), .o(n_19895) );
no02f80 g744801 ( .a(n_35192), .b(n_30587), .o(n_35284) );
no02f80 g750395 ( .a(FE_OCP_RBN3525_n_29624), .b(n_29626), .o(n_29662) );
in01f80 newInst_1855 ( .a(newNet_1854), .o(newNet_1855) );
in01f80 newInst_2005 ( .a(newNet_2004), .o(newNet_2005) );
na02f80 FE_RC_2485_0 ( .a(n_9730), .b(FE_RN_1003_0), .o(FE_RN_1004_0) );
na02f80 g760833 ( .a(n_19585), .b(n_18119), .o(n_19615) );
no02f80 g737341 ( .a(n_42834), .b(n_42594), .o(n_42843) );
in01f80 g779508 ( .a(n_1446), .o(n_1447) );
no02f80 g767272 ( .a(n_13413), .b(n_13412), .o(n_13414) );
ao22s80 FE_RC_824_0 ( .a(n_28822), .b(n_29384), .c(n_28823), .d(n_29383), .o(n_29479) );
no02f80 FE_RC_633_0 ( .a(FE_RN_197_0), .b(n_17798), .o(n_17887) );
in01f80 g754041 ( .a(n_26221), .o(n_26306) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_0_ ( .ck(newNet_2601), .d(n_26111), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_) );
in01f80 FE_OCP_RBC1103_n_45224 ( .a(FE_OCP_RBN3267_n_45224), .o(FE_OCP_RBN1103_n_45224) );
no02f80 g755589 ( .a(n_24715), .b(n_24714), .o(n_24716) );
oa12f80 g742870 ( .a(n_37229), .b(n_37228), .c(n_37227), .o(n_37847) );
na02f80 g779171 ( .a(n_1890), .b(n_1857), .o(n_1901) );
na02f80 g769618 ( .a(n_11277), .b(n_11251), .o(n_11327) );
no02f80 g744525 ( .a(n_35370), .b(n_35256), .o(n_35401) );
no02f80 FE_RC_3110_0 ( .a(FE_RN_1375_0), .b(FE_RN_1376_0), .o(n_27028) );
in01f80 FE_RC_2518_0 ( .a(n_37109), .o(FE_RN_1025_0) );
na02f80 g740975 ( .a(n_39109), .b(n_38900), .o(n_39143) );
oa12f80 g759253 ( .a(n_21258), .b(n_21263), .c(n_21257), .o(n_21341) );
na02f80 g775190 ( .a(n_46996), .b(n_6030), .o(n_6066) );
no02f80 g772428 ( .a(n_8503), .b(n_7952), .o(n_8518) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_14_ ( .ck(newNet_3253), .d(n_36310), .o(delay_add_ln22_unr23_stage9_stallmux_q_14_) );
oa22f80 FE_RC_948_0 ( .a(n_22907), .b(n_22806), .c(n_20252), .d(n_22776), .o(n_22872) );
no02f80 g766958 ( .a(n_13670), .b(n_13643), .o(n_13740) );
in01f80 newInst_1412 ( .a(newNet_1411), .o(newNet_1412) );
na02f80 g776675 ( .a(n_4301), .b(n_4329), .o(n_4553) );
no02f80 g737444 ( .a(n_42703), .b(n_42357), .o(n_42718) );
in01f80 FE_OCP_RBC3269_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3269_n_45224) );
oa22f80 g752718 ( .a(n_27161), .b(n_27082), .c(n_27128), .d(n_27081), .o(n_27279) );
na02f80 g741578 ( .a(n_38657), .b(n_38685), .o(n_38755) );
in01f80 g750559 ( .a(n_29494), .o(n_29520) );
in01f80 newInst_1542 ( .a(newNet_1541), .o(newNet_1542) );
na02f80 g778479 ( .a(n_2340), .b(FE_OCPN3759_n_2346), .o(n_2347) );
oa12f80 g740517 ( .a(n_39689), .b(n_39676), .c(n_39675), .o(n_39716) );
in01f80 g771080 ( .a(n_9959), .o(n_9960) );
na02f80 g775163 ( .a(n_6015), .b(n_5822), .o(n_6016) );
na02f80 g764418 ( .a(n_16013), .b(n_14588), .o(n_16206) );
na02f80 g779207 ( .a(n_1905), .b(n_944), .o(n_1969) );
ao22s80 g736404 ( .a(n_43780), .b(n_43580), .c(n_43779), .d(n_43579), .o(n_43835) );
na02f80 g744674 ( .a(n_35184), .b(n_35119), .o(n_35186) );
in01f80 newInst_1450 ( .a(newNet_1449), .o(newNet_1450) );
in01f80 g778232 ( .a(n_2749), .o(n_2750) );
no02f80 g758220 ( .a(n_22725), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_26_), .o(n_23006) );
in01f80 newInst_668 ( .a(newNet_667), .o(newNet_668) );
no02f80 g773783 ( .a(n_7188), .b(n_7187), .o(n_7189) );
in01f80 newInst_2744 ( .a(newNet_2556), .o(newNet_2744) );
na02f80 g773715 ( .a(n_7327), .b(n_7364), .o(n_7933) );
na02f80 g740374 ( .a(n_39803), .b(n_39832), .o(n_39854) );
oa22f80 FE_RC_47_0 ( .a(n_4671), .b(n_4736), .c(FE_OCP_RBN2538_n_3645), .d(n_4730), .o(n_4916) );
na02f80 FE_RC_851_0 ( .a(FE_RN_252_0), .b(FE_RN_253_0), .o(FE_RN_254_0) );
no02f80 g747980 ( .a(n_33048), .b(n_33146), .o(n_33092) );
na02f80 g750479 ( .a(n_29570), .b(n_29526), .o(n_29607) );
no02f80 g759069 ( .a(FE_OCP_RBN1712_n_21087), .b(n_21011), .o(n_21166) );
oa12f80 g749114 ( .a(n_31394), .b(n_32158), .c(n_31220), .o(n_32232) );
in01f80 g774461 ( .a(n_6626), .o(n_6684) );
oa22f80 FE_RC_1133_0 ( .a(n_7712), .b(FE_OCP_RBN2330_n_9003), .c(n_9003), .d(FE_OCPN1241_n_7721), .o(n_8077) );
in01f80 newInst_2353 ( .a(newNet_2352), .o(newNet_2353) );
in01f80 fopt783568 ( .a(n_39648), .o(n_45188) );
in01f80 newInst_1296 ( .a(newNet_267), .o(newNet_1296) );
in01f80 g759724 ( .a(n_21827), .o(n_21828) );
no02f80 FE_RC_4194_0 ( .a(n_18594), .b(n_19034), .o(FE_RN_1838_0) );
in01f80 FE_OCP_RBC2300_n_7817 ( .a(n_7817), .o(FE_OCP_RBN2300_n_7817) );
no02f80 g764390 ( .a(n_16161), .b(n_16193), .o(n_16319) );
in01f80 g764489 ( .a(n_16157), .o(n_16188) );
no02f80 g771935 ( .a(n_8747), .b(n_7600), .o(n_8741) );
ao12f80 g757276 ( .a(n_23308), .b(n_44066), .c(delay_xor_ln22_unr15_stage6_stallmux_q_10_), .o(n_23074) );
in01f80 g736612 ( .a(n_43626), .o(n_43636) );
no02f80 g741285 ( .a(n_44955), .b(n_38573), .o(n_38998) );
ao12f80 g765368 ( .a(n_15715), .b(n_15874), .c(n_14652), .o(n_16546) );
no02f80 g773809 ( .a(n_7180), .b(n_6687), .o(n_7206) );
na02f80 g741994 ( .a(n_38089), .b(n_37984), .o(n_38085) );
no02f80 g740550 ( .a(n_39692), .b(n_45739), .o(n_39713) );
na02f80 g765879 ( .a(n_14880), .b(n_14808), .o(n_14903) );
in01f80 newInst_1618 ( .a(newNet_1593), .o(newNet_1618) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_21_ ( .ck(newNet_338), .d(n_1297), .o(delay_xor_ln22_unr3_stage2_stallmux_q_21_) );
in01f80 g741969 ( .a(n_38114), .o(n_38115) );
na02f80 g763365 ( .a(n_16905), .b(n_16998), .o(n_17039) );
in01f80 g772441 ( .a(n_8496), .o(n_8497) );
no02f80 g760380 ( .a(n_20740), .b(n_20042), .o(n_20834) );
na02f80 g748223 ( .a(FE_OCP_RBN3732_n_31819), .b(n_31740), .o(n_32139) );
ao12f80 g758137 ( .a(n_22877), .b(n_23115), .c(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_), .o(n_23201) );
in01f80 FE_OCP_RBC2733_n_4219 ( .a(FE_OCP_RBN2732_n_4219), .o(FE_OCP_RBN2733_n_4219) );
in01f80 newInst_1445 ( .a(newNet_590), .o(newNet_1445) );
ao12f80 g780729 ( .a(n_448), .b(n_608), .c(n_460), .o(n_612) );
no02f80 g764572 ( .a(n_15948), .b(n_14524), .o(n_16004) );
in01f80 FE_OCP_RBC2829_n_30731 ( .a(n_30731), .o(FE_OCP_RBN2829_n_30731) );
no02f80 g777202 ( .a(n_3534), .b(n_2731), .o(n_3582) );
in01f80 newInst_2933 ( .a(newNet_2932), .o(newNet_2933) );
no02f80 g753842 ( .a(n_26300), .b(FE_OCP_RBN2883_n_26292), .o(n_26399) );
oa22f80 FE_RC_3790_0 ( .a(n_22961), .b(FE_OCP_RBN3119_n_22755), .c(n_22833), .d(n_22755), .o(n_22834) );
na02f80 g740010 ( .a(n_39823), .b(n_39816), .o(n_39876) );
na02f80 g738083 ( .a(n_42041), .b(n_41905), .o(n_42060) );
no02f80 g763517 ( .a(n_17576), .b(n_17429), .o(n_17632) );
no02f80 g759980 ( .a(FE_OCP_RBN1358_FE_RN_677_0), .b(n_20407), .o(n_20468) );
na02f80 g780163 ( .a(n_1139), .b(n_1122), .o(n_1123) );
ao12f80 g745121 ( .a(FE_OCPN3779_n_36126), .b(n_36127), .c(n_35724), .o(n_36232) );
no02f80 g748162 ( .a(n_31947), .b(n_31863), .o(n_32057) );
in01f80 g750883 ( .a(n_29110), .o(n_29136) );
in01f80 g743992 ( .a(n_36365), .o(n_36366) );
in01f80 g752483 ( .a(n_27771), .o(n_27744) );
no02f80 g751716 ( .a(n_28385), .b(n_28381), .o(n_28382) );
in01f80 g756546 ( .a(n_23767), .o(n_23713) );
in01f80 newInst_620 ( .a(newNet_619), .o(newNet_620) );
in01f80 FE_OCPC1243_n_44460 ( .a(FE_OCPN997_n_44460), .o(FE_OCPN1243_n_44460) );
in01f80 newInst_3414 ( .a(newNet_3413), .o(newNet_3414) );
no02f80 g761461 ( .a(n_19647), .b(n_19735), .o(n_19830) );
no02f80 g776707 ( .a(n_47013), .b(n_3951), .o(n_4053) );
no02f80 g747734 ( .a(n_33239), .b(n_33372), .o(n_33812) );
oa22f80 g754607 ( .a(n_26133), .b(n_25740), .c(n_26132), .d(n_25739), .o(n_26740) );
in01f80 g761455 ( .a(n_19710), .o(n_19711) );
in01f80 g779749 ( .a(n_1673), .o(n_1674) );
in01f80 newInst_3268 ( .a(newNet_2037), .o(newNet_3268) );
oa12f80 g755422 ( .a(n_25348), .b(n_25347), .c(n_25346), .o(n_25440) );
in01f80 newInst_140 ( .a(newNet_139), .o(newNet_140) );
in01f80 g780786 ( .a(n_429), .o(n_430) );
no02f80 g763333 ( .a(n_17132), .b(n_17033), .o(n_17233) );
oa12f80 g748958 ( .a(n_31150), .b(n_31149), .c(n_31148), .o(n_31193) );
no02f80 g754539 ( .a(n_26311), .b(n_26271), .o(n_26312) );
no02f80 g743507 ( .a(n_37699), .b(n_37631), .o(n_37728) );
na02f80 g744059 ( .a(n_44221), .b(n_35742), .o(n_35784) );
na02f80 g737880 ( .a(n_42202), .b(n_42103), .o(n_42310) );
no02f80 g753107 ( .a(n_27250), .b(n_27173), .o(n_27301) );
in01f80 g757855 ( .a(n_23121), .o(n_23183) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_13_ ( .ck(newNet_2680), .d(n_22112), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_13_) );
na02f80 g777343 ( .a(n_4556), .b(n_4797), .o(n_5005) );
in01f80 g771797 ( .a(n_8906), .o(n_8907) );
oa12f80 g747772 ( .a(n_33357), .b(n_33571), .c(n_33314), .o(n_33892) );
in01f80 g743292 ( .a(n_38019), .o(n_38020) );
na02f80 g759304 ( .a(n_20889), .b(FE_RN_1585_0), .o(n_20922) );
na02f80 FE_RC_1952_0 ( .a(FE_RN_626_0), .b(FE_RN_627_0), .o(FE_RN_628_0) );
na02f80 g739140 ( .a(n_40943), .b(n_40885), .o(n_40944) );
na02f80 g780419 ( .a(n_815), .b(n_1098), .o(n_823) );
no02f80 FE_RC_1759_0 ( .a(FE_RN_499_0), .b(FE_RN_500_0), .o(FE_RN_501_0) );
na02f80 FE_RC_2677_0 ( .a(n_4083), .b(n_4134), .o(FE_RN_1120_0) );
no02f80 g751938 ( .a(n_28102), .b(n_28041), .o(n_28126) );
in01f80 FE_OCP_RBC3540_n_8784 ( .a(n_8784), .o(FE_OCP_RBN3540_n_8784) );
no02f80 g749417 ( .a(n_30603), .b(n_30246), .o(n_30604) );
na02f80 g770958 ( .a(n_10042), .b(n_8426), .o(n_10129) );
in01f80 g772708 ( .a(n_8163), .o(n_8185) );
in01f80 g774958 ( .a(n_6225), .o(n_6226) );
na02f80 g742414 ( .a(n_37737), .b(n_37764), .o(n_37759) );
in01f80 newInst_1917 ( .a(newNet_1916), .o(newNet_1917) );
na02f80 g765082 ( .a(FE_OCP_RBN2762_n_15200), .b(FE_OCPN1007_n_13962), .o(n_15283) );
in01f80 g747862 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_13_), .o(n_32083) );
no02f80 g766217 ( .a(n_14731), .b(n_14205), .o(n_14836) );
na02f80 g769342 ( .a(n_10035), .b(FE_OCP_RBN2104_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11634) );
in01f80 g777644 ( .a(n_3418), .o(n_3419) );
ao12f80 g741917 ( .a(n_37954), .b(n_38074), .c(n_38073), .o(n_38075) );
ao12f80 g759390 ( .a(n_21144), .b(n_21054), .c(n_21055), .o(n_21263) );
ao12f80 g756384 ( .a(n_23937), .b(n_24330), .c(n_23952), .o(n_24415) );
no02f80 g770188 ( .a(n_10785), .b(FE_OFN345_n_9247), .o(n_10903) );
in01f80 newInst_1151 ( .a(newNet_1150), .o(newNet_1151) );
no02f80 g757048 ( .a(n_23646), .b(n_22883), .o(n_23702) );
no02f80 g745843 ( .a(n_44104), .b(n_33975), .o(n_34302) );
na02f80 g748949 ( .a(n_32313), .b(n_46107), .o(n_32455) );
na02f80 g759566 ( .a(n_20689), .b(n_20594), .o(n_20730) );
no02f80 g745859 ( .a(n_34124), .b(n_34038), .o(n_34164) );
no02f80 g776268 ( .a(n_4752), .b(n_4798), .o(n_4954) );
in01f80 FE_OCP_RBC3097_n_6313 ( .a(n_6313), .o(FE_OCP_RBN3097_n_6313) );
in01f80 newInst_3176 ( .a(newNet_2546), .o(newNet_3176) );
no02f80 g744094 ( .a(n_44222), .b(n_34713), .o(n_35752) );
ao12f80 g738154 ( .a(n_42034), .b(n_42033), .c(n_42032), .o(n_42076) );
no02f80 g751339 ( .a(n_29463), .b(n_29462), .o(n_29464) );
in01f80 FE_OCP_RBC2592_n_25181 ( .a(n_25181), .o(FE_OCP_RBN2592_n_25181) );
in01f80 g754745 ( .a(n_26741), .o(n_26633) );
no02f80 g759174 ( .a(n_21264), .b(n_45026), .o(n_21314) );
in01f80 newInst_1209 ( .a(newNet_470), .o(newNet_1209) );
oa12f80 g736483 ( .a(n_43373), .b(n_43711), .c(n_43366), .o(n_43739) );
in01f80 FE_RC_2731_0 ( .a(n_22748), .o(FE_RN_1156_0) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_21_ ( .ck(newNet_2751), .d(n_17459), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_) );
no02f80 g772963 ( .a(n_7820), .b(n_7819), .o(n_7865) );
na02f80 g744899 ( .a(n_35075), .b(FE_OCPN1794_n_30612), .o(n_35094) );
no02f80 g742147 ( .a(FE_OCP_RBN2256_n_37844), .b(n_37555), .o(n_38038) );
na02f80 g747806 ( .a(n_33571), .b(n_33651), .o(n_33740) );
ao12f80 g741076 ( .a(n_38952), .b(FE_OCPN957_n_39096), .c(n_38930), .o(n_39366) );
in01f80 g749815 ( .a(n_31617), .o(n_31618) );
in01f80 newInst_154 ( .a(newNet_91), .o(newNet_154) );
in01f80 g739749 ( .a(n_40475), .o(n_40476) );
in01f80 newInst_2719 ( .a(newNet_2718), .o(newNet_2719) );
in01f80 newInst_1697 ( .a(newNet_1696), .o(newNet_1697) );
na02f80 g747046 ( .a(n_32795), .b(delay_xor_ln21_unr21_stage8_stallmux_q_10_), .o(n_32863) );
no02f80 g748272 ( .a(FE_OCP_RBN3084_n_31819), .b(n_46959), .o(n_31947) );
in01f80 g757367 ( .a(n_23038), .o(n_23039) );
oa12f80 g764800 ( .a(n_15599), .b(n_16177), .c(n_16244), .o(n_16265) );
no02f80 g766947 ( .a(n_13937), .b(n_13904), .o(n_14260) );
na02f80 FE_RC_2522_0 ( .a(FE_RN_1026_0), .b(n_40809), .o(FE_RN_1027_0) );
no02f80 g777621 ( .a(n_3482), .b(n_2913), .o(n_3573) );
na02f80 g749909 ( .a(n_29925), .b(n_29901), .o(n_29902) );
in01f80 g750956 ( .a(n_28968), .o(n_28969) );
oa12f80 g754978 ( .a(n_24983), .b(n_25118), .c(n_25035), .o(n_25128) );
na02f80 g759550 ( .a(n_20820), .b(n_20797), .o(n_20798) );
no02f80 g775904 ( .a(n_5193), .b(n_4503), .o(n_5262) );
oa22f80 FE_RC_1138_0 ( .a(n_1534), .b(FE_OCP_RBN3381_n_1732), .c(n_1535), .d(n_1732), .o(n_1827) );
no02f80 g764437 ( .a(n_16011), .b(FE_OCPN3775_n_14730), .o(n_16057) );
in01f80 FE_RC_4018_0 ( .a(n_45008), .o(FE_RN_1745_0) );
in01f80 FE_RC_1040_0 ( .a(n_32621), .o(FE_RN_301_0) );
no02f80 g751825 ( .a(n_28230), .b(n_28014), .o(n_28254) );
oa12f80 g759483 ( .a(n_20962), .b(n_20961), .c(n_20960), .o(n_21027) );
in01f80 FE_OCPC1863_n_26171 ( .a(n_26171), .o(FE_OCPN1863_n_26171) );
na02f80 g766915 ( .a(n_14258), .b(n_14296), .o(n_14947) );
na02f80 g779231 ( .a(n_1900), .b(n_1899), .o(n_2040) );
na02f80 g744657 ( .a(n_35186), .b(FE_OCP_RBN2656_FE_RN_1288_0), .o(n_35275) );
oa12f80 g756393 ( .a(n_24241), .b(n_24259), .c(n_24240), .o(n_25000) );
no02f80 g779058 ( .a(n_2105), .b(n_1881), .o(n_2118) );
na02f80 g743462 ( .a(n_37728), .b(n_37727), .o(n_37729) );
oa12f80 g743227 ( .a(n_36864), .b(n_36903), .c(n_36883), .o(n_36908) );
no02f80 g745632 ( .a(n_34248), .b(n_34250), .o(n_34249) );
in01f80 g753352 ( .a(n_27120), .o(n_27207) );
oa12f80 g744998 ( .a(n_34931), .b(n_34930), .c(n_34929), .o(n_35659) );
no02f80 g741973 ( .a(n_37953), .b(n_37945), .o(n_38015) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_11_ ( .ck(newNet_2685), .d(n_21969), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_) );
in01f80 FE_RC_183_0 ( .a(n_50), .o(FE_RN_61_0) );
in01f80 g758775 ( .a(n_21656), .o(n_21657) );
in01f80 g747296 ( .a(n_32752), .o(n_32753) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_22_ ( .ck(newNet_235), .d(n_46190), .o(delay_xor_ln22_unr6_stage3_stallmux_q_22_) );
in01f80 g758224 ( .a(n_22732), .o(n_22688) );
in01f80 g764503 ( .a(n_16267), .o(n_16422) );
in01f80 g755673 ( .a(FE_OCP_RBN2423_n_24501), .o(n_24555) );
oa22f80 FE_RC_1482_0 ( .a(n_32287), .b(n_32512), .c(n_28336), .d(n_32427), .o(n_32541) );
in01f80 FE_RC_2348_0 ( .a(n_1669), .o(FE_RN_901_0) );
in01f80 g748746 ( .a(n_32505), .o(n_32506) );
na02f80 g775241 ( .a(n_5902), .b(n_5761), .o(n_5928) );
na02f80 g757662 ( .a(n_22615), .b(n_22708), .o(n_22746) );
in01f80 g780236 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_18_), .o(n_1037) );
no02f80 g744115 ( .a(n_35729), .b(n_35690), .o(n_35782) );
no02f80 g776449 ( .a(n_4178), .b(n_4202), .o(n_4324) );
in01f80 g769592 ( .a(n_11425), .o(n_11581) );
no02f80 g768411 ( .a(n_12492), .b(n_12477), .o(n_12478) );
no02f80 g749146 ( .a(n_32205), .b(n_31453), .o(n_32230) );
na02f80 g738463 ( .a(n_41759), .b(n_41762), .o(n_41763) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_19_ ( .ck(newNet_3325), .d(n_32147), .o(delay_add_ln22_unr20_stage8_stallmux_q_19_) );
no02f80 g767025 ( .a(n_14758), .b(n_14256), .o(n_14347) );
in01f80 g771455 ( .a(n_9560), .o(n_9561) );
na02f80 g738516 ( .a(n_41420), .b(n_41634), .o(n_41676) );
in01f80 g748254 ( .a(n_32055), .o(n_32070) );
na02f80 g760814 ( .a(n_19366), .b(n_18787), .o(n_19476) );
no02f80 g773217 ( .a(n_7674), .b(n_7673), .o(n_7727) );
in01f80 FE_OCPC1027_n_4182 ( .a(n_4182), .o(FE_OCPN1027_n_4182) );
in01f80 g766010 ( .a(n_14669), .o(n_14670) );
in01f80 g740145 ( .a(n_39843), .o(n_40047) );
ao22s80 g780857 ( .a(n_457), .b(n_368), .c(n_420), .d(n_372), .o(n_533) );
no02f80 g756087 ( .a(n_24223), .b(n_24199), .o(n_24263) );
in01f80 newInst_2911 ( .a(newNet_2910), .o(newNet_2911) );
na02f80 g778056 ( .a(n_2914), .b(n_2264), .o(n_2944) );
ao22s80 g781135 ( .a(n_215), .b(n_134), .c(n_214), .d(n_133), .o(n_398) );
oa12f80 g744663 ( .a(n_36125), .b(n_36513), .c(n_35960), .o(n_36598) );
na02f80 g737064 ( .a(n_43230), .b(n_43243), .o(n_43483) );
in01f80 g770575 ( .a(n_10197), .o(n_10230) );
in01f80 newInst_967 ( .a(newNet_610), .o(newNet_967) );
na02f80 g760453 ( .a(n_20624), .b(n_20599), .o(n_20600) );
na02f80 g780630 ( .a(n_779), .b(n_859), .o(n_951) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_3_ ( .ck(newNet_790), .d(n_1291), .o(delay_xor_ln21_unr3_stage2_stallmux_q_3_) );
in01f80 g766759 ( .a(n_13732), .o(n_13778) );
oa12f80 g766987 ( .a(n_13738), .b(n_13737), .c(n_13736), .o(n_14216) );
oa12f80 g767081 ( .a(n_13578), .b(n_13612), .c(n_13517), .o(n_13684) );
in01f80 g766984 ( .a(n_13877), .o(n_13878) );
no02f80 g742070 ( .a(FE_OCP_RBN3446_n_37945), .b(FE_OCP_RBN2175_n_37559), .o(n_38087) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_28_ ( .ck(newNet_797), .d(n_1289), .o(delay_xor_ln21_unr3_stage2_stallmux_q_28_) );
oa12f80 g749804 ( .a(n_31460), .b(n_31311), .c(n_31145), .o(n_31643) );
na02f80 g768384 ( .a(n_12504), .b(n_12149), .o(n_12542) );
na02f80 g751495 ( .a(n_28600), .b(n_28545), .o(n_28624) );
ao12f80 g756370 ( .a(n_24381), .b(n_24380), .c(n_24379), .o(n_24980) );
no02f80 g758517 ( .a(n_21953), .b(FE_OCP_RBN1364_n_20412), .o(n_22003) );
in01f80 g769452 ( .a(n_11480), .o(n_11456) );
ao22s80 FE_RC_1608_0 ( .a(n_25722), .b(n_26324), .c(n_26376), .d(n_25721), .o(n_26464) );
na02f80 g758296 ( .a(n_22288), .b(n_21087), .o(n_22407) );
no02f80 g754013 ( .a(n_26156), .b(n_26038), .o(n_26157) );
na02f80 g755446 ( .a(n_24821), .b(n_24612), .o(n_24867) );
in01f80 g752518 ( .a(n_27726), .o(n_27704) );
in01f80 newInst_186 ( .a(newNet_185), .o(newNet_186) );
in01f80 FE_RC_2469_0 ( .a(n_14035), .o(FE_RN_994_0) );
no02f80 g770069 ( .a(n_10823), .b(n_10875), .o(n_10957) );
oa12f80 g744939 ( .a(n_34651), .b(n_34994), .c(n_34993), .o(n_35026) );
in01f80 g752732 ( .a(n_27237), .o(n_27238) );
no02f80 g777165 ( .a(n_4216), .b(n_4292), .o(n_4910) );
na02f80 g742672 ( .a(n_37399), .b(n_37278), .o(n_37416) );
oa12f80 g739197 ( .a(n_45149), .b(n_40763), .c(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n_40865) );
no02f80 g752333 ( .a(n_44723), .b(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .o(n_27864) );
na02f80 g775024 ( .a(n_6155), .b(n_6136), .o(n_6248) );
no02f80 g747333 ( .a(n_32637), .b(n_44962), .o(n_32666) );
na02f80 g750384 ( .a(n_29635), .b(n_29647), .o(n_29716) );
na02f80 g754915 ( .a(n_25327), .b(n_25390), .o(n_25424) );
na02f80 FE_RC_3722_0 ( .a(n_14871), .b(n_14959), .o(FE_RN_1637_0) );
oa12f80 g772469 ( .a(n_8470), .b(n_8469), .c(n_8468), .o(n_9544) );
oa12f80 g745353 ( .a(n_35962), .b(FE_OCP_RBN2995_n_35539), .c(n_35884), .o(n_36155) );
oa22f80 FE_RC_4030_0 ( .a(n_26061), .b(n_26068), .c(n_26028), .d(n_26062), .o(n_26184) );
oa22f80 FE_RC_3773_0 ( .a(n_18538), .b(n_19281), .c(n_18537), .d(n_19280), .o(n_19390) );
no02f80 g756585 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_), .o(n_23850) );
no02f80 g745036 ( .a(n_34771), .b(n_34256), .o(n_34829) );
na02f80 g740527 ( .a(n_39722), .b(n_39695), .o(n_39732) );
no02f80 g743783 ( .a(n_35989), .b(n_36151), .o(n_36152) );
no02f80 g755632 ( .a(n_24593), .b(n_24554), .o(n_24715) );
oa12f80 g776952 ( .a(n_3768), .b(n_3985), .c(n_3883), .o(n_4139) );
no02f80 g748425 ( .a(FE_OCP_RBN3713_n_31466), .b(n_31655), .o(n_32197) );
in01f80 g777968 ( .a(n_3210), .o(n_3211) );
in01f80 newInst_1763 ( .a(newNet_1762), .o(newNet_1763) );
oa12f80 g745873 ( .a(n_35339), .b(n_35338), .c(n_35337), .o(n_35388) );
no02f80 g743114 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_), .o(n_37092) );
in01f80 FE_RC_3194_0 ( .a(n_7246), .o(FE_RN_1419_0) );
in01f80 newInst_1283 ( .a(newNet_1282), .o(newNet_1283) );
ms00f80 delay_xor_ln21_unr6_stage3_stallmux_q_reg_21_ ( .ck(newNet_718), .d(n_46184), .o(delay_xor_ln21_unr6_stage3_stallmux_q_21_) );
in01f80 FE_RC_2578_0 ( .a(n_2913), .o(FE_RN_1062_0) );
in01f80 newInst_3740 ( .a(newNet_3739), .o(newNet_3740) );
na02f80 g780296 ( .a(n_786), .b(n_765), .o(n_766) );
na02f80 g762683 ( .a(n_17850), .b(n_17896), .o(n_17924) );
na02f80 g776464 ( .a(n_4509), .b(n_4571), .o(n_4720) );
in01f80 newInst_3435 ( .a(newNet_3434), .o(newNet_3435) );
ao12f80 g764941 ( .a(FE_OCP_RBN2681_n_15048), .b(FE_OCPN1257_n_13831), .c(n_15286), .o(n_15356) );
in01f80 g767661 ( .a(FE_OCP_RBN2223_n_12902), .o(n_12877) );
in01f80 g781140 ( .a(n_214), .o(n_215) );
in01f80 g739311 ( .a(n_40885), .o(n_40700) );
na02f80 g780702 ( .a(n_636), .b(n_509), .o(n_646) );
in01f80 g750013 ( .a(n_31040), .o(n_31064) );
no02f80 g772959 ( .a(n_7784), .b(n_8453), .o(n_7793) );
in01f80 g752814 ( .a(n_27851), .o(n_27852) );
in01f80 g737382 ( .a(n_42821), .o(n_42822) );
no02f80 FE_RC_3699_0 ( .a(n_17133), .b(FE_RN_1627_0), .o(n_17188) );
no02f80 g757215 ( .a(n_23491), .b(n_23181), .o(n_23546) );
in01f80 g754271 ( .a(n_25940), .o(n_25918) );
in01f80 FE_OCP_RBC2826_FE_RN_1573_0 ( .a(FE_RN_1573_0), .o(FE_OCP_RBN2826_FE_RN_1573_0) );
no02f80 g741989 ( .a(n_37980), .b(n_37406), .o(n_37953) );
na02f80 g739185 ( .a(n_40866), .b(n_40778), .o(n_41084) );
ao12f80 g764354 ( .a(n_16203), .b(n_16288), .c(n_16224), .o(n_16371) );
in01f80 g769952 ( .a(n_11212), .o(n_11184) );
oa12f80 g747851 ( .a(n_32104), .b(FE_OCP_RBN1212_n_32142), .c(n_31903), .o(n_32236) );
in01f80 g739417 ( .a(n_40725), .o(n_40810) );
in01f80 newInst_3723 ( .a(newNet_3722), .o(newNet_3723) );
na02f80 g744495 ( .a(n_35444), .b(n_35343), .o(n_35445) );
in01f80 g756849 ( .a(n_23369), .o(n_23370) );
na02f80 g740034 ( .a(n_39866), .b(n_39846), .o(n_39984) );
no02f80 g763304 ( .a(n_17076), .b(n_17120), .o(n_17190) );
in01f80 newInst_1823 ( .a(newNet_1822), .o(newNet_1823) );
in01f80 newInst_259 ( .a(newNet_49), .o(newNet_259) );
in01f80 g750715 ( .a(FE_OCP_RBN2310_n_29298), .o(n_30191) );
na02f80 g762044 ( .a(n_18910), .b(n_18738), .o(n_18964) );
no02f80 g745637 ( .a(n_34286), .b(n_33617), .o(n_34490) );
na02f80 g738876 ( .a(n_41307), .b(n_41306), .o(n_41308) );
na02f80 g753666 ( .a(n_26540), .b(n_44325), .o(n_26564) );
no02f80 FE_RC_2477_0 ( .a(n_40060), .b(n_40057), .o(FE_RN_999_0) );
na02f80 g764222 ( .a(n_16513), .b(n_16512), .o(n_16601) );
in01f80 g753326 ( .a(n_27151), .o(n_27113) );
no02f80 g740267 ( .a(n_40131), .b(n_40130), .o(n_40171) );
no02f80 g739209 ( .a(n_40859), .b(n_40843), .o(n_40860) );
in01f80 g753379 ( .a(n_27110), .o(n_27167) );
na02f80 g760736 ( .a(n_19560), .b(n_18117), .o(n_19604) );
in01f80 FE_OCP_RBC2233_n_13141 ( .a(FE_OCP_RBN2232_n_13141), .o(FE_OCP_RBN2233_n_13141) );
na02f80 FE_RC_1124_0 ( .a(FE_RN_339_0), .b(FE_RN_340_0), .o(FE_RN_341_0) );
na02f80 g767506 ( .a(n_13057), .b(n_13146), .o(n_13229) );
na02f80 g737765 ( .a(n_42215), .b(n_42232), .o(n_42233) );
no02f80 g771092 ( .a(n_9515), .b(n_8452), .o(n_9726) );
in01f80 newInst_1986 ( .a(newNet_1985), .o(newNet_1986) );
in01f80 FE_OCPC3181_FE_OCP_RBN2831_n_10198 ( .a(FE_OCP_RBN2831_n_10198), .o(FE_OCPN3181_FE_OCP_RBN2831_n_10198) );
in01f80 newInst_598 ( .a(newNet_41), .o(newNet_598) );
in01f80 newInst_484 ( .a(newNet_483), .o(newNet_484) );
no02f80 g753828 ( .a(n_26429), .b(n_26428), .o(n_26462) );
in01f80 FE_OCP_RBC1202_n_25898 ( .a(n_25898), .o(FE_OCP_RBN1202_n_25898) );
in01f80 FE_OCP_RBC3615_n_20249 ( .a(FE_OCP_RBN2670_n_20249), .o(FE_OCP_RBN3615_n_20249) );
in01f80 g769582 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_17_), .o(n_11391) );
in01f80 g774240 ( .a(n_6637), .o(n_6638) );
na02f80 g781111 ( .a(n_233), .b(n_232), .o(n_234) );
na02f80 g779155 ( .a(n_1915), .b(delay_add_ln22_unr2_stage2_stallmux_q_11_), .o(n_1979) );
na02f80 g740348 ( .a(n_40204), .b(n_40166), .o(n_40304) );
ao12f80 g784650 ( .a(n_15738), .b(n_15649), .c(n_15696), .o(n_46980) );
in01f80 g747051 ( .a(n_33015), .o(n_33035) );
in01f80 g769022 ( .a(n_11760), .o(n_11845) );
na02f80 g745710 ( .a(n_34337), .b(n_44102), .o(n_34452) );
ao22s80 g736324 ( .a(n_43810), .b(n_43398), .c(n_43809), .d(n_43399), .o(n_43856) );
in01f80 g762354 ( .a(n_18495), .o(n_18496) );
na02f80 g743927 ( .a(n_35748), .b(n_44222), .o(n_35830) );
no02f80 g780880 ( .a(n_403), .b(n_424), .o(n_441) );
no02f80 g737908 ( .a(n_42202), .b(n_41910), .o(n_42213) );
na02f80 g767287 ( .a(n_13511), .b(FE_OCPN1428_n_13510), .o(n_13578) );
na02f80 g747280 ( .a(n_32691), .b(n_32623), .o(n_32732) );
in01f80 FE_RC_2293_0 ( .a(n_28128), .o(FE_RN_862_0) );
oa22f80 g759798 ( .a(n_21714), .b(n_20809), .c(n_21691), .d(n_21591), .o(n_21857) );
no02f80 g748391 ( .a(FE_OCP_RBN3714_n_31466), .b(n_30507), .o(n_31735) );
ao12f80 g754737 ( .a(n_25771), .b(n_26161), .c(n_25736), .o(n_26235) );
no02f80 g737066 ( .a(n_43230), .b(n_43243), .o(n_43292) );
oa12f80 g749598 ( .a(n_30421), .b(n_30483), .c(n_30443), .o(n_30486) );
in01f80 FE_OCP_RBC2674_n_14991 ( .a(FE_OCP_RBN2673_n_14991), .o(FE_OCP_RBN2674_n_14991) );
in01f80 newInst_1372 ( .a(newNet_1340), .o(newNet_1372) );
in01f80 g771757 ( .a(n_10381), .o(n_10382) );
no02f80 FE_RC_2912_0 ( .a(FE_RN_1266_0), .b(n_12980), .o(FE_RN_1267_0) );
no02f80 g745648 ( .a(n_34272), .b(n_34246), .o(n_34385) );
in01f80 FE_OCPC1797_n_20333 ( .a(n_20333), .o(FE_OCPN1797_n_20333) );
na02f80 g744791 ( .a(FE_OCP_RBN2657_FE_RN_1288_0), .b(n_35119), .o(n_35146) );
na02f80 g738023 ( .a(n_42153), .b(n_42146), .o(n_42169) );
na02f80 g769913 ( .a(n_10991), .b(n_44463), .o(n_11033) );
na02f80 g778714 ( .a(n_2365), .b(n_2357), .o(n_2452) );
na02f80 g776345 ( .a(n_4399), .b(n_4495), .o(n_4580) );
in01f80 g745345 ( .a(n_36113), .o(n_36114) );
ao12f80 g770871 ( .a(FE_OCP_RBN2759_n_9843), .b(n_10171), .c(n_9999), .o(n_10212) );
no02f80 g737692 ( .a(n_42285), .b(n_42312), .o(n_42334) );
in01f80 FE_OCP_RBC2722_n_4219 ( .a(n_4219), .o(FE_OCP_RBN2722_n_4219) );
na02f80 g756432 ( .a(n_24114), .b(n_24113), .o(n_24115) );
no02f80 g784780 ( .a(n_44222), .b(n_35906), .o(n_47266) );
oa22f80 g774029 ( .a(n_6823), .b(n_6601), .c(n_6760), .d(n_6602), .o(n_6874) );
in01f80 FE_OCP_RBC2886_n_10570 ( .a(n_10570), .o(FE_OCP_RBN2886_n_10570) );
na02f80 g753765 ( .a(FE_OCP_RBN2969_n_26398), .b(n_23509), .o(n_26472) );
no02f80 g743862 ( .a(n_37814), .b(n_36863), .o(n_37898) );
oa12f80 g767264 ( .a(n_13202), .b(n_13716), .c(n_13088), .o(n_13762) );
oa12f80 g768811 ( .a(n_11753), .b(n_11823), .c(n_11676), .o(n_11922) );
no02f80 g776833 ( .a(n_3851), .b(n_3754), .o(n_3954) );
in01f80 FE_OCP_RBC2564_FE_RN_1125_0 ( .a(FE_RN_1125_0), .o(FE_OCP_RBN2564_FE_RN_1125_0) );
in01f80 FE_OCPC1257_n_13831 ( .a(FE_OCPN1256_n_13831), .o(FE_OCPN1257_n_13831) );
no02f80 g753675 ( .a(n_27203), .b(n_26738), .o(n_27284) );
no02f80 g774100 ( .a(n_6759), .b(n_6691), .o(n_6797) );
in01f80 FE_OCP_RBC2814_n_25817 ( .a(n_25817), .o(FE_OCP_RBN2814_n_25817) );
in01f80 g779598 ( .a(n_1882), .o(n_1883) );
in01f80 FE_OCP_RBC2524_n_8951 ( .a(FE_OCP_RBN2523_n_8951), .o(FE_OCP_RBN2524_n_8951) );
no02f80 g760753 ( .a(n_19596), .b(n_19564), .o(n_19688) );
in01f80 g759028 ( .a(n_21281), .o(n_21282) );
na02f80 FE_RC_4247_0 ( .a(n_26842), .b(FE_RN_1867_0), .o(FE_RN_1868_0) );
in01f80 g754858 ( .a(n_25724), .o(n_25725) );
na02f80 g762977 ( .a(n_17959), .b(n_17958), .o(n_17960) );
no02f80 g744268 ( .a(n_44174), .b(n_34919), .o(n_35620) );
ao12f80 g784682 ( .a(n_3942), .b(n_3894), .c(n_3792), .o(n_47012) );
in01f80 g772350 ( .a(n_8504), .o(n_8546) );
in01f80 newInst_2872 ( .a(newNet_2871), .o(newNet_2872) );
na02f80 g757691 ( .a(FE_OCP_RBN3818_n_44061), .b(n_45204), .o(n_22582) );
no02f80 g737187 ( .a(n_42978), .b(n_42965), .o(n_42998) );
oa12f80 g766244 ( .a(n_14400), .b(n_14365), .c(n_14318), .o(n_14508) );
no02f80 g776711 ( .a(n_3731), .b(n_3728), .o(n_3838) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_6_ ( .ck(newNet_3279), .d(n_31363), .o(delay_add_ln22_unr20_stage8_stallmux_q_6_) );
na02f80 FE_RC_1917_0 ( .a(n_18331), .b(FE_OCP_RBN2205_n_18242), .o(FE_RN_604_0) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_28_ ( .ck(newNet_3399), .d(n_27771), .o(delay_add_ln22_unr17_stage7_stallmux_q_28_) );
ao12f80 g768098 ( .a(n_12220), .b(n_12663), .c(n_12046), .o(n_12711) );
oa12f80 g769103 ( .a(FE_OCPN858_n_45697), .b(n_11889), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n_12013) );
na02f80 g775315 ( .a(n_5933), .b(n_4784), .o(n_6011) );
oa12f80 g751377 ( .a(FE_OCPN987_n_28402), .b(n_28535), .c(FE_OCPN989_n_28353), .o(n_28611) );
na02f80 g748264 ( .a(FE_OCP_RBN3730_n_31819), .b(n_30608), .o(n_32019) );
in01f80 newInst_222 ( .a(newNet_221), .o(newNet_222) );
in01f80 g763443 ( .a(n_17120), .o(n_17174) );
na02f80 g775481 ( .a(n_5505), .b(n_5496), .o(n_5614) );
ao12f80 g755769 ( .a(n_24442), .b(n_24393), .c(n_24336), .o(n_24549) );
in01f80 g772823 ( .a(n_7943), .o(n_7944) );
na02f80 g740909 ( .a(n_39340), .b(n_39370), .o(n_39864) );
oa22f80 g739842 ( .a(n_40234), .b(n_39984), .c(n_40235), .d(n_39985), .o(n_40350) );
in01f80 g736771 ( .a(n_43318), .o(n_43319) );
na02f80 g748375 ( .a(n_31476), .b(n_30323), .o(n_31501) );
no02f80 g765342 ( .a(n_15112), .b(n_15049), .o(n_15153) );
oa12f80 g770378 ( .a(n_10145), .b(n_10404), .c(n_10116), .o(n_10541) );
no02f80 g776084 ( .a(n_4840), .b(n_4804), .o(n_4841) );
in01f80 g777406 ( .a(n_3485), .o(n_3533) );
na02f80 g770993 ( .a(n_9666), .b(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .o(n_9806) );
in01f80 g773960 ( .a(n_7002), .o(n_7003) );
na02f80 g766316 ( .a(n_14271), .b(FE_OCP_RBN2250_n_13017), .o(n_14332) );
no02f80 g743845 ( .a(n_35674), .b(n_35553), .o(n_35835) );
in01f80 FE_OCPC1734_n_16143 ( .a(FE_OCPN1733_n_16143), .o(FE_OCPN1734_n_16143) );
in01f80 newInst_3450 ( .a(newNet_430), .o(newNet_3450) );
in01f80 g739170 ( .a(n_40914), .o(n_40895) );
no02f80 g776929 ( .a(n_4014), .b(n_3938), .o(n_4072) );
in01f80 g758647 ( .a(n_21849), .o(n_21847) );
oa22f80 FE_RC_3936_0 ( .a(n_22769), .b(n_22672), .c(n_22575), .d(n_22673), .o(n_22827) );
in01f80 g770845 ( .a(n_10015), .o(n_11253) );
in01f80 g739866 ( .a(n_40261), .o(n_40262) );
na02f80 FE_RC_1055_0 ( .a(FE_OFN783_delay_sub_ln23_0_unr15_stage6_stallmux_q), .b(n_24181), .o(FE_RN_309_0) );
in01f80 g781087 ( .a(n_476), .o(n_261) );
in01f80 newInst_3390 ( .a(newNet_2174), .o(newNet_3390) );
in01f80 g741850 ( .a(n_38484), .o(n_38508) );
no02f80 g784775 ( .a(n_15103), .b(n_14169), .o(n_47261) );
no02f80 g767244 ( .a(n_13537), .b(n_13552), .o(n_13597) );
no02f80 g762442 ( .a(n_18049), .b(n_18048), .o(n_18071) );
oa12f80 g766847 ( .a(n_47253), .b(n_13689), .c(n_13017), .o(n_13702) );
in01f80 FE_RC_2274_0 ( .a(n_17609), .o(FE_RN_847_0) );
in01f80 g773930 ( .a(n_7055), .o(n_7004) );
na02f80 g747383 ( .a(n_33574), .b(n_33576), .o(n_33577) );
in01f80 FE_RC_631_0 ( .a(n_17797), .o(FE_RN_196_0) );
na02f80 g744103 ( .a(n_35898), .b(FE_OCP_RBN2902_n_44174), .o(n_35976) );
in01f80 newInst_1740 ( .a(newNet_1739), .o(newNet_1740) );
no02f80 g780454 ( .a(n_1203), .b(n_1099), .o(n_878) );
na02f80 g749869 ( .a(FE_OCP_RBN3011_n_31117), .b(n_31277), .o(n_31344) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_25_ ( .ck(newNet_1833), .d(n_16967), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_25_) );
no02f80 g765001 ( .a(n_15429), .b(n_14419), .o(n_15430) );
in01f80 newInst_3286 ( .a(newNet_2234), .o(newNet_3286) );
in01f80 g745225 ( .a(n_34415), .o(n_34358) );
no02f80 g741597 ( .a(FE_OCP_RBN2484_n_38601), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38631) );
in01f80 FE_RC_3409_0 ( .a(n_21090), .o(FE_RN_1476_0) );
no02f80 g738228 ( .a(n_41949), .b(n_41947), .o(n_41948) );
oa12f80 g776379 ( .a(n_4106), .b(n_4608), .c(n_4170), .o(n_4697) );
in01f80 newInst_3711 ( .a(newNet_2977), .o(newNet_3711) );
in01f80 g755946 ( .a(n_24267), .o(n_25316) );
na02f80 g762080 ( .a(FE_OCP_RBN2205_n_18242), .b(n_17692), .o(n_18394) );
na02f80 g751284 ( .a(n_29742), .b(n_29741), .o(n_29743) );
na02f80 g760584 ( .a(n_19886), .b(FE_OFN816_n_19885), .o(n_19968) );
ao12f80 g763760 ( .a(n_17308), .b(n_17207), .c(n_17152), .o(n_17469) );
ao22s80 FE_RC_2941_0 ( .a(n_5832), .b(n_5854), .c(n_5816), .d(n_5833), .o(n_5989) );
in01f80 newInst_2232 ( .a(newNet_2231), .o(newNet_2232) );
in01f80 g754611 ( .a(FE_OCPN1410_n_27014), .o(n_27062) );
no02f80 g772808 ( .a(n_8115), .b(n_8114), .o(n_8159) );
in01f80 g747358 ( .a(n_32549), .o(n_32550) );
na02f80 g751044 ( .a(n_30126), .b(n_30099), .o(n_30785) );
no02f80 g737571 ( .a(n_42377), .b(n_42287), .o(n_42316) );
ao12f80 g769125 ( .a(n_11372), .b(n_11480), .c(n_11479), .o(n_11523) );
in01f80 g750053 ( .a(n_29960), .o(n_29982) );
in01f80 g773472 ( .a(n_7558), .o(n_7553) );
in01f80 newInst_1358 ( .a(newNet_32), .o(newNet_1358) );
ao12f80 g745119 ( .a(n_34684), .b(n_34683), .c(n_34682), .o(n_34751) );
ao12f80 g780796 ( .a(n_360), .b(n_386), .c(n_367), .o(n_528) );
in01f80 FE_RC_1950_0 ( .a(n_25418), .o(FE_RN_626_0) );
na02f80 g746602 ( .a(FE_OCP_RBN2598_n_34388), .b(n_34547), .o(n_34644) );
in01f80 g741192 ( .a(n_39421), .o(n_39422) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_26_ ( .ck(newNet_2374), .d(n_36569), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_) );
in01f80 FE_OCP_RBC3643_n_44490 ( .a(FE_OCP_RBN3639_n_44490), .o(FE_OCP_RBN3643_n_44490) );
in01f80 g760782 ( .a(n_20155), .o(n_20201) );
in01f80 FE_RC_4142_0 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(FE_RN_1799_0) );
no02f80 g753636 ( .a(n_26659), .b(n_26658), .o(n_26660) );
oa12f80 g753468 ( .a(n_26763), .b(FE_OCP_RBN2983_n_26767), .c(n_26762), .o(n_26807) );
in01f80 g739220 ( .a(n_40783), .o(n_40784) );
in01f80 g774210 ( .a(n_7024), .o(n_7025) );
in01f80 g752035 ( .a(n_28123), .o(n_28145) );
in01f80 g737171 ( .a(n_43032), .o(n_43030) );
na02f80 g751753 ( .a(n_28272), .b(n_28062), .o(n_28307) );
na02f80 g769827 ( .a(n_46987), .b(n_9682), .o(n_11235) );
ao12f80 g773991 ( .a(n_6950), .b(n_6949), .c(n_6948), .o(n_7788) );
na02f80 g742971 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n_36975) );
in01f80 g765769 ( .a(FE_OCP_RBN2715_n_14982), .o(n_15105) );
in01f80 g764170 ( .a(n_16600), .o(n_16620) );
in01f80 newInst_3224 ( .a(newNet_3223), .o(newNet_3224) );
no02f80 g771418 ( .a(n_9118), .b(n_9095), .o(n_9313) );
in01f80 fopt783049 ( .a(n_44498), .o(n_44511) );
oa12f80 g750286 ( .a(n_29698), .b(n_29735), .c(n_29660), .o(n_29755) );
in01f80 g754123 ( .a(n_26140), .o(n_26141) );
na02f80 g783834 ( .a(n_14586), .b(n_14612), .o(n_45520) );
no02f80 g745188 ( .a(FE_OCP_DRV_N1594_n_34494), .b(n_34466), .o(n_34467) );
in01f80 g767491 ( .a(n_13151), .o(n_13152) );
oa12f80 g738895 ( .a(n_41203), .b(n_41202), .c(n_41201), .o(n_41254) );
in01f80 g769598 ( .a(n_11318), .o(n_11335) );
no02f80 g743193 ( .a(n_36918), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_), .o(n_37030) );
no03m80 FE_RC_374_0 ( .a(n_11882), .b(FE_OCP_RBN2136_n_11907), .c(n_11991), .o(n_11992) );
in01f80 FE_OCP_DRV_C3153_n_24425 ( .a(n_24425), .o(FE_OCP_DRV_N3153_n_24425) );
in01f80 newInst_1094 ( .a(newNet_1093), .o(newNet_1094) );
na02f80 g750990 ( .a(n_28871), .b(n_28581), .o(n_28935) );
in01f80 g755397 ( .a(n_24784), .o(n_24785) );
in01f80 g770786 ( .a(n_9860), .o(n_9861) );
ao12f80 g779476 ( .a(n_1703), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_14_), .o(n_1824) );
no02f80 g762369 ( .a(n_45002), .b(n_18689), .o(n_18769) );
in01f80 g746849 ( .a(n_33260), .o(n_33261) );
na02f80 g777906 ( .a(n_3189), .b(n_2759), .o(n_3243) );
no02f80 g760484 ( .a(n_19950), .b(n_19948), .o(n_19949) );
in01f80 g765921 ( .a(n_14775), .o(n_14802) );
na02f80 g777086 ( .a(n_3881), .b(n_3690), .o(n_4036) );
no02f80 g742101 ( .a(n_37876), .b(n_37910), .o(n_37911) );
in01f80 newInst_3181 ( .a(newNet_3180), .o(newNet_3181) );
in01f80 g767062 ( .a(n_14205), .o(n_14206) );
in01f80 g769643 ( .a(n_11383), .o(n_11400) );
in01f80 newInst_2322 ( .a(newNet_2234), .o(newNet_2322) );
no02f80 g748079 ( .a(n_31746), .b(n_31687), .o(n_31810) );
in01f80 newInst_1271 ( .a(newNet_1270), .o(newNet_1271) );
in01f80 g747641 ( .a(n_32255), .o(n_32240) );
in01f80 g770004 ( .a(n_10915), .o(n_10916) );
ao12f80 g768297 ( .a(n_12546), .b(n_12545), .c(n_12544), .o(n_12985) );
in01f80 newInst_2151 ( .a(newNet_2150), .o(newNet_2151) );
in01f80 g773128 ( .a(n_7698), .o(n_7699) );
ao12f80 g761512 ( .a(n_19647), .b(n_19051), .c(n_19733), .o(n_20058) );
na02f80 g777173 ( .a(n_4361), .b(n_4426), .o(n_4460) );
in01f80 newInst_3562 ( .a(newNet_3561), .o(newNet_3562) );
in01f80 g774319 ( .a(n_6870), .o(n_6871) );
in01f80 g757539 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_7_), .o(n_22935) );
in01f80 newInst_547 ( .a(newNet_546), .o(newNet_547) );
na02f80 g748435 ( .a(FE_OCPN1052_n_31674), .b(FE_OCP_RBN2921_n_31107), .o(n_31757) );
ao12f80 g759828 ( .a(n_21247), .b(n_21691), .c(n_21294), .o(n_22008) );
oa12f80 g744008 ( .a(n_35536), .b(n_35537), .c(n_35535), .o(n_35578) );
na02f80 g771203 ( .a(n_9450), .b(n_8362), .o(n_9594) );
oa22f80 g743664 ( .a(n_36373), .b(n_36366), .c(n_36374), .d(n_36365), .o(n_36430) );
in01f80 fopt783793 ( .a(n_17723), .o(n_45472) );
no02f80 g745320 ( .a(n_35850), .b(n_35796), .o(n_35851) );
in01f80 FE_OCP_RBC3249_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_ ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(FE_OCP_RBN3249_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_) );
oa12f80 g749082 ( .a(n_31569), .b(n_32205), .c(n_31409), .o(n_32249) );
no02f80 g750277 ( .a(n_29751), .b(n_28582), .o(n_29810) );
na02f80 g760065 ( .a(n_20752), .b(n_20705), .o(n_20812) );
no02f80 g738704 ( .a(n_41491), .b(n_41490), .o(n_41533) );
no02f80 g761286 ( .a(n_19034), .b(n_18546), .o(n_19036) );
na02f80 g769890 ( .a(n_11108), .b(n_11159), .o(n_11178) );
in01f80 g743775 ( .a(n_37292), .o(n_37293) );
no02f80 g750641 ( .a(n_30419), .b(n_30418), .o(n_30420) );
na02f80 g778959 ( .a(n_2129), .b(n_2128), .o(n_2130) );
oa22f80 g757625 ( .a(n_22564), .b(n_22167), .c(n_45721), .d(n_22165), .o(n_22718) );
oa22f80 g781146 ( .a(n_203), .b(n_96), .c(n_202), .d(n_97), .o(n_385) );
na02f80 g767626 ( .a(n_12866), .b(n_12829), .o(n_12980) );
no02f80 g779429 ( .a(n_1397), .b(n_1399), .o(n_1460) );
no02f80 g770824 ( .a(n_9809), .b(n_8538), .o(n_9862) );
oa22f80 g749169 ( .a(n_32153), .b(n_31623), .c(n_32152), .d(n_31624), .o(n_32229) );
oa22f80 g784351 ( .a(FE_OFN774_n_46137), .b(FE_OCP_RBN3097_n_6313), .c(n_46195), .d(n_6313), .o(n_46157) );
na02f80 g778687 ( .a(n_2277), .b(n_2276), .o(n_2308) );
no02f80 g746728 ( .a(n_34231), .b(n_34230), .o(n_34232) );
oa22f80 g780223 ( .a(n_1008), .b(n_1099), .c(n_1056), .d(n_1098), .o(n_1134) );
oa12f80 g741891 ( .a(n_38250), .b(n_38242), .c(n_38310), .o(n_38383) );
ao12f80 g767624 ( .a(n_13253), .b(n_13346), .c(n_13315), .o(n_13347) );
no02f80 g747425 ( .a(n_32613), .b(n_44962), .o(n_32631) );
in01f80 g768565 ( .a(n_12342), .o(n_12343) );
in01f80 g746856 ( .a(n_33140), .o(n_33141) );
no02f80 g758730 ( .a(n_21662), .b(n_21577), .o(n_21710) );
in01f80 g761839 ( .a(n_18475), .o(n_18476) );
in01f80 newInst_2377 ( .a(newNet_2376), .o(newNet_2377) );
ao12f80 g742157 ( .a(n_37865), .b(n_37864), .c(n_37863), .o(n_38764) );
in01f80 FE_RC_4232_0 ( .a(n_25916), .o(FE_RN_1858_0) );
in01f80 g778639 ( .a(n_2299), .o(n_2278) );
no02f80 g755076 ( .a(n_25693), .b(n_25644), .o(n_25719) );
no02f80 g748334 ( .a(FE_OCP_RBN3084_n_31819), .b(n_30654), .o(n_31993) );
ao12f80 g768380 ( .a(n_12417), .b(n_12362), .c(n_12416), .o(n_12469) );
no02f80 g750891 ( .a(n_30106), .b(n_29818), .o(n_30168) );
in01f80 FE_RC_3610_0 ( .a(FE_RN_1579_0), .o(n_26842) );
oa12f80 g767999 ( .a(n_12667), .b(n_12616), .c(n_12666), .o(n_12728) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_4_ ( .ck(newNet_3002), .d(n_958), .o(delay_add_ln22_unr2_stage2_stallmux_q_4_) );
na02f80 g770573 ( .a(n_10021), .b(n_9974), .o(n_10101) );
na02f80 g737024 ( .a(n_43097), .b(n_42773), .o(n_43217) );
oa22f80 FE_RC_3391_0 ( .a(n_36268), .b(FE_OCP_RBN3066_n_36547), .c(n_36269), .d(n_36547), .o(n_36651) );
in01f80 g765244 ( .a(n_15635), .o(n_15636) );
no02f80 g774311 ( .a(n_6863), .b(n_6862), .o(n_7428) );
in01f80 g768536 ( .a(n_12370), .o(n_12349) );
in01f80 g768840 ( .a(n_12402), .o(n_12059) );
in01f80 g766113 ( .a(n_14632), .o(n_14633) );
oa12f80 g746775 ( .a(n_32892), .b(n_33063), .c(delay_sub_ln21_0_unr20_stage8_stallmux_q_27_), .o(n_33065) );
in01f80 newInst_1852 ( .a(newNet_1851), .o(newNet_1852) );
in01f80 g741300 ( .a(n_38876), .o(n_38877) );
no02f80 g763412 ( .a(n_16876), .b(n_16837), .o(n_16995) );
na02f80 g772864 ( .a(n_8017), .b(n_8016), .o(n_8122) );
ao12f80 g747315 ( .a(n_33843), .b(n_33842), .c(n_33841), .o(n_33910) );
na02f80 g751826 ( .a(n_28228), .b(n_28227), .o(n_28284) );
na02f80 g764370 ( .a(n_16285), .b(n_14730), .o(n_16286) );
in01f80 g758746 ( .a(n_21665), .o(n_21711) );
in01f80 g776295 ( .a(n_4630), .o(n_4706) );
in01f80 g757584 ( .a(delay_add_ln22_unr14_stage6_stallmux_q_19_), .o(n_23611) );
na02f80 g739476 ( .a(FE_OCPN897_n_44776), .b(n_40737), .o(n_41006) );
no02f80 g758843 ( .a(n_21476), .b(n_45026), .o(n_21509) );
na02f80 g762717 ( .a(n_17828), .b(n_17804), .o(n_17932) );
no02f80 g738675 ( .a(n_41564), .b(n_41563), .o(n_41607) );
in01f80 newInst_1753 ( .a(newNet_1752), .o(newNet_1753) );
na02f80 g769872 ( .a(n_11000), .b(n_10998), .o(n_11056) );
in01f80 g749769 ( .a(n_31631), .o(n_31632) );
no02f80 g776796 ( .a(n_4212), .b(n_4211), .o(n_4248) );
na02f80 g769299 ( .a(n_11407), .b(n_11379), .o(n_11482) );
na02f80 g780463 ( .a(n_1203), .b(FE_OFN50_n_1045), .o(n_872) );
na02f80 g769906 ( .a(n_10915), .b(n_44498), .o(n_10939) );
in01f80 newInst_806 ( .a(newNet_805), .o(newNet_806) );
no02f80 g742072 ( .a(FE_OCP_RBN3444_n_37945), .b(n_38032), .o(n_38112) );
no02f80 g758085 ( .a(n_44268), .b(n_44160), .o(n_22481) );
no02f80 g755090 ( .a(n_24972), .b(n_25024), .o(n_25025) );
oa12f80 g754958 ( .a(n_25288), .b(n_25868), .c(FE_RN_871_0), .o(n_25923) );
in01f80 g756012 ( .a(n_25735), .o(n_25736) );
in01f80 newInst_3559 ( .a(newNet_3558), .o(newNet_3559) );
in01f80 newInst_2718 ( .a(newNet_2717), .o(newNet_2718) );
in01f80 g774563 ( .a(n_6521), .o(n_6585) );
na02f80 g746079 ( .a(n_33735), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33785) );
in01f80 g750567 ( .a(n_29485), .o(n_29507) );
oa12f80 g743638 ( .a(n_36012), .b(n_36352), .c(n_35821), .o(n_36398) );
na02f80 g772658 ( .a(n_8275), .b(n_8273), .o(n_8274) );
in01f80 FE_OCP_RBC3109_n_43711 ( .a(n_43711), .o(FE_OCP_RBN3109_n_43711) );
no02f80 g745363 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35258), .o(n_35805) );
in01f80 g737427 ( .a(n_42772), .o(n_42773) );
na02f80 g755357 ( .a(n_24963), .b(FE_OCPN1744_n_24962), .o(n_24983) );
in01f80 g754499 ( .a(n_25595), .o(n_25596) );
in01f80 newInst_2200 ( .a(newNet_257), .o(newNet_2200) );
na02f80 g748832 ( .a(n_31265), .b(n_31264), .o(n_31352) );
in01f80 g768313 ( .a(n_12638), .o(n_12639) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_17_ ( .ck(newNet_353), .d(n_1338), .o(delay_xor_ln22_unr3_stage2_stallmux_q_17_) );
na02f80 g768336 ( .a(n_12484), .b(n_12512), .o(n_12533) );
in01f80 newInst_1141 ( .a(newNet_362), .o(newNet_1141) );
in01f80 g749425 ( .a(n_30542), .o(n_30543) );
no02f80 g757992 ( .a(n_47278), .b(n_22194), .o(n_22230) );
in01f80 g737590 ( .a(n_42788), .o(n_42789) );
na02f80 g768020 ( .a(n_12703), .b(n_12702), .o(n_12704) );
in01f80 newInst_903 ( .a(newNet_902), .o(newNet_903) );
in01f80 g759246 ( .a(n_21264), .o(n_21265) );
na02f80 g766932 ( .a(n_14041), .b(n_14138), .o(n_14700) );
in01f80 newInst_3271 ( .a(newNet_3270), .o(newNet_3271) );
no02f80 g749037 ( .a(n_31093), .b(n_31148), .o(n_31095) );
na02f80 g751597 ( .a(n_28447), .b(n_28541), .o(n_28542) );
na02f80 g770114 ( .a(n_10700), .b(n_10280), .o(n_10764) );
oa22f80 FE_RC_4273_0 ( .a(n_17377), .b(n_17660), .c(n_17376), .d(n_17695), .o(n_17835) );
ao12f80 g748100 ( .a(n_32808), .b(n_32807), .c(n_32806), .o(n_33310) );
na02f80 g781018 ( .a(sin_out_6), .b(FE_OFN3_n_43918), .o(n_326) );
ao12f80 g749977 ( .a(n_30318), .b(n_29869), .c(n_29530), .o(n_30319) );
in01f80 FE_OCP_RBC3074_n_43230 ( .a(FE_OCP_RBN3069_n_43230), .o(FE_OCP_RBN3074_n_43230) );
in01f80 newInst_1189 ( .a(newNet_736), .o(newNet_1189) );
no02f80 g746640 ( .a(n_34359), .b(n_34332), .o(n_34333) );
in01f80 FE_OCP_RBC2723_n_4219 ( .a(n_4219), .o(FE_OCP_RBN2723_n_4219) );
no02f80 g775300 ( .a(n_5644), .b(n_4556), .o(n_5672) );
in01f80 g761306 ( .a(n_19098), .o(n_19099) );
in01f80 newInst_431 ( .a(newNet_430), .o(newNet_431) );
in01f80 g772445 ( .a(n_8651), .o(n_8686) );
in01f80 newInst_1202 ( .a(newNet_1201), .o(newNet_1202) );
na02f80 g775814 ( .a(n_5359), .b(n_5013), .o(n_5420) );
oa22f80 FE_RC_1129_0 ( .a(n_12500), .b(n_12690), .c(n_12501), .d(n_12691), .o(n_12771) );
in01f80 FE_OCP_RBC1912_n_20965 ( .a(n_20965), .o(FE_OCP_RBN1912_n_20965) );
na02f80 g772848 ( .a(n_7969), .b(n_7331), .o(n_8011) );
na02f80 g781163 ( .a(state_cordic_1_), .b(mux_while_ln12_psv_q_3_), .o(n_198) );
in01f80 g777182 ( .a(n_5174), .o(n_5175) );
na02f80 g759426 ( .a(n_21059), .b(FE_OCPUNCON3146_n_21058), .o(n_21114) );
no02f80 g759668 ( .a(n_20508), .b(n_20294), .o(n_20553) );
no02f80 g749223 ( .a(n_30821), .b(n_30846), .o(n_30958) );
na02f80 g754922 ( .a(n_25327), .b(n_24419), .o(n_25385) );
na02f80 g762022 ( .a(n_18394), .b(n_18393), .o(n_18427) );
in01f80 newInst_260 ( .a(newNet_259), .o(newNet_260) );
no02f80 g757301 ( .a(n_44066), .b(delay_xor_ln22_unr15_stage6_stallmux_q_13_), .o(n_23022) );
no02f80 g781332 ( .a(n_7), .b(beta_23), .o(n_140) );
no02f80 g739363 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_30_), .o(n_40932) );
na02f80 g771030 ( .a(n_9644), .b(n_9717), .o(n_9895) );
na02f80 g743889 ( .a(n_35954), .b(n_35822), .o(n_36011) );
na02f80 g748189 ( .a(n_31705), .b(n_31730), .o(n_31776) );
oa22f80 FE_RC_48_0 ( .a(n_5066), .b(n_5347), .c(n_5065), .d(n_5346), .o(n_5490) );
na02f80 g778531 ( .a(n_2550), .b(n_1197), .o(n_2658) );
na02f80 g761435 ( .a(n_18868), .b(n_18371), .o(n_18900) );
no02f80 g767544 ( .a(n_13007), .b(n_12984), .o(n_13141) );
na02f80 g740189 ( .a(n_39798), .b(n_39797), .o(n_39799) );
na02f80 g743623 ( .a(n_36416), .b(n_36041), .o(n_36445) );
in01f80 g777091 ( .a(n_3926), .o(n_4121) );
in01f80 g766643 ( .a(n_13948), .o(n_14019) );
in01f80 g770144 ( .a(n_10672), .o(n_10673) );
in01f80 FE_OCP_RBC3408_n_28597 ( .a(FE_OCP_RBN3406_n_28597), .o(FE_OCP_RBN3408_n_28597) );
na02f80 g745714 ( .a(n_34120), .b(n_44101), .o(n_34150) );
oa22f80 g739591 ( .a(FE_OCP_RBN3338_n_44610), .b(delay_xor_ln21_unr28_stage10_stallmux_q_3_), .c(n_40624), .d(n_44610), .o(n_40643) );
in01f80 g764040 ( .a(n_17900), .o(n_19170) );
na02f80 g760506 ( .a(n_19970), .b(n_19803), .o(n_20001) );
na02f80 g744909 ( .a(n_34959), .b(n_34936), .o(n_35029) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_14_ ( .ck(newNet_2312), .d(n_40385), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_14_) );
in01f80 FE_OCP_DRV_C3167_FE_RN_1789_0 ( .a(FE_RN_1789_0), .o(FE_OCP_DRV_N3167_FE_RN_1789_0) );
na02f80 g767788 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_24_), .o(n_12867) );
na02f80 g752354 ( .a(n_27884), .b(n_27821), .o(n_27934) );
na02f80 g777694 ( .a(n_3365), .b(n_2880), .o(n_3423) );
in01f80 g776629 ( .a(n_4302), .o(n_4303) );
no02f80 g760610 ( .a(n_19747), .b(n_18230), .o(n_19859) );
in01f80 fopt782907 ( .a(n_44355), .o(n_44354) );
in01f80 g742038 ( .a(n_38258), .o(n_38259) );
in01f80 g753205 ( .a(n_27426), .o(n_27388) );
no02f80 g740758 ( .a(n_39535), .b(n_40183), .o(n_39536) );
na02f80 g779008 ( .a(n_2106), .b(n_1953), .o(n_2107) );
no02f80 g746928 ( .a(n_32860), .b(n_32329), .o(n_32897) );
in01f80 FE_RC_1794_0 ( .a(n_28083), .o(FE_RN_529_0) );
no03m80 g746344 ( .a(n_33411), .b(n_33163), .c(n_33020), .o(n_33494) );
in01f80 FE_OCPC3752_n_1448 ( .a(n_1448), .o(FE_OCPN3752_n_1448) );
no02f80 g748642 ( .a(n_32609), .b(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_32629) );
in01f80 newInst_2334 ( .a(newNet_553), .o(newNet_2334) );
na02f80 g749462 ( .a(n_31888), .b(n_31323), .o(n_31981) );
in01f80 newInst_3278 ( .a(newNet_3277), .o(newNet_3278) );
na03f80 FE_RC_1212_0 ( .a(n_41348), .b(n_41332), .c(n_44428), .o(n_41362) );
na02f80 FE_RC_678_0 ( .a(n_17583), .b(FE_RN_218_0), .o(n_17667) );
oa22f80 FE_RC_4024_0 ( .a(n_35347), .b(n_35225), .c(n_35346), .d(n_35226), .o(n_35421) );
in01f80 g760995 ( .a(n_19377), .o(n_19378) );
oa22f80 FE_RC_3348_0 ( .a(n_17136), .b(n_17626), .c(n_17191), .d(n_17600), .o(n_17782) );
oa22f80 FE_RC_3298_0 ( .a(n_34558), .b(n_34876), .c(n_34877), .d(n_34559), .o(n_34980) );
in01f80 g748815 ( .a(n_32530), .o(n_32531) );
oa22f80 g752706 ( .a(n_27238), .b(n_27043), .c(n_27237), .d(n_27042), .o(n_27360) );
no02f80 g754316 ( .a(n_25763), .b(n_25831), .o(n_25793) );
in01f80 g773051 ( .a(n_7752), .o(n_7724) );
in01f80 newInst_1835 ( .a(newNet_1834), .o(newNet_1835) );
na02f80 g762748 ( .a(n_18015), .b(n_17965), .o(n_18036) );
no02f80 g740415 ( .a(FE_OCP_RBN3022_n_39942), .b(n_39495), .o(n_40131) );
na02f80 g738405 ( .a(n_41701), .b(n_41300), .o(n_41702) );
in01f80 newInst_986 ( .a(newNet_985), .o(newNet_986) );
no02f80 g773183 ( .a(FE_OCP_RBN2228_n_7598), .b(n_8568), .o(n_7680) );
in01f80 FE_OCPC854_n_45450 ( .a(FE_OCPN853_n_45450), .o(FE_OCPN854_n_45450) );
ao12f80 g755322 ( .a(n_25223), .b(n_25410), .c(n_25084), .o(n_25470) );
in01f80 g779877 ( .a(n_1356), .o(n_1360) );
ao12f80 g773444 ( .a(n_6904), .b(n_7516), .c(n_6817), .o(n_7528) );
in01f80 newInst_1884 ( .a(newNet_1470), .o(newNet_1884) );
in01f80 g766790 ( .a(n_13690), .o(n_13707) );
na02f80 g769087 ( .a(n_11752), .b(n_11580), .o(n_11808) );
in01f80 newInst_867 ( .a(newNet_866), .o(newNet_867) );
na02f80 g766167 ( .a(n_14592), .b(FE_OCP_RBN2506_n_13896), .o(n_14655) );
in01f80 FE_OCP_RBC3435_n_29163 ( .a(n_29163), .o(FE_OCP_RBN3435_n_29163) );
na02f80 FE_RC_2341_0 ( .a(FE_RN_896_0), .b(n_47211), .o(n_12296) );
no02f80 g750480 ( .a(n_29483), .b(n_29407), .o(n_29529) );
oa12f80 g773805 ( .a(n_7139), .b(n_7144), .c(n_7138), .o(n_8099) );
na02f80 g746833 ( .a(n_33053), .b(n_33099), .o(n_33423) );
ms00f80 delay_xor_ln22_unr21_stage8_stallmux_q_reg_2_ ( .ck(newNet_414), .d(n_32545), .o(delay_xor_ln22_unr21_stage8_stallmux_q_2_) );
na02f80 g745270 ( .a(n_35933), .b(n_35956), .o(n_35995) );
in01f80 FE_RC_1203_0 ( .a(n_17488), .o(FE_RN_363_0) );
in01f80 g763654 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_15_), .o(n_18159) );
oa12f80 g743136 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_17_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_16_), .o(n_37210) );
no02f80 g774352 ( .a(FE_OCP_RBN1982_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_7_), .o(n_6651) );
no02f80 g739332 ( .a(n_45144), .b(n_40696), .o(n_40734) );
in01f80 newInst_64 ( .a(newNet_63), .o(newNet_64) );
no02f80 g770948 ( .a(n_9682), .b(FE_OFN755_n_44461), .o(n_9753) );
in01f80 g739734 ( .a(n_40524), .o(n_40501) );
in01f80 g738475 ( .a(n_41426), .o(n_41427) );
in01f80 newInst_3326 ( .a(newNet_1280), .o(newNet_3326) );
oa12f80 g765116 ( .a(n_15264), .b(n_15415), .c(n_15339), .o(n_15532) );
in01f80 g767042 ( .a(n_13973), .o(n_14039) );
in01f80 FE_OCP_RBC2904_n_10474 ( .a(n_10474), .o(FE_OCP_RBN2904_n_10474) );
in01f80 newInst_1329 ( .a(newNet_1328), .o(newNet_1329) );
in01f80 g743453 ( .a(n_36612), .o(n_36613) );
na02f80 g738595 ( .a(n_41502), .b(n_41501), .o(n_41503) );
oa12f80 g784336 ( .a(n_5384), .b(n_6315), .c(n_6304), .o(n_46137) );
na02f80 FE_RC_2342_0 ( .a(n_18659), .b(n_18658), .o(FE_RN_897_0) );
no02f80 g765143 ( .a(n_15638), .b(n_15788), .o(n_15721) );
in01f80 g768409 ( .a(n_12523), .o(n_12524) );
in01f80 g740062 ( .a(n_40143), .o(n_40144) );
na02f80 g749360 ( .a(n_30723), .b(FE_OCPN1410_n_27014), .o(n_30817) );
na03f80 FE_RC_3808_0 ( .a(n_22231), .b(n_22153), .c(n_22232), .o(n_22273) );
na03f80 FE_RC_3216_0 ( .a(n_8584), .b(n_8595), .c(n_8663), .o(n_8729) );
no02f80 g755682 ( .a(n_25438), .b(n_25437), .o(n_25439) );
no02f80 g763895 ( .a(n_17498), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_17_), .o(n_17308) );
in01f80 g758101 ( .a(n_22047), .o(n_22078) );
in01f80 newInst_2188 ( .a(newNet_2187), .o(newNet_2188) );
in01f80 g737339 ( .a(n_42889), .o(n_42855) );
na02f80 FE_RC_510_0 ( .a(FE_RN_156_0), .b(FE_RN_157_0), .o(FE_RN_158_0) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_27_ ( .ck(newNet_1299), .d(n_1274), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_27_) );
no02f80 g740686 ( .a(n_39474), .b(n_39500), .o(n_39540) );
no02f80 g759960 ( .a(n_20416), .b(n_20381), .o(n_20501) );
ao12f80 g755027 ( .a(n_22484), .b(n_25048), .c(n_24829), .o(n_25117) );
in01f80 newInst_2637 ( .a(newNet_2296), .o(newNet_2637) );
na02f80 g754851 ( .a(n_25399), .b(n_25275), .o(n_25400) );
oa22f80 g750874 ( .a(FE_OCP_RBN1905_n_29080), .b(n_29109), .c(FE_OCP_RBN1906_n_29080), .d(n_27914), .o(n_30671) );
in01f80 newInst_50 ( .a(newNet_32), .o(newNet_50) );
na02f80 g758791 ( .a(n_21587), .b(n_45081), .o(n_21684) );
na02f80 FE_RC_2050_0 ( .a(n_25966), .b(FE_RN_691_0), .o(FE_RN_692_0) );
na02f80 g780583 ( .a(n_666), .b(n_672), .o(n_669) );
na02f80 g777082 ( .a(n_3677), .b(n_3705), .o(n_3743) );
in01f80 g772265 ( .a(n_8692), .o(n_8709) );
in01f80 drc784124 ( .a(n_45872), .o(n_45873) );
ao12f80 g765866 ( .a(n_15211), .b(n_15210), .c(n_15209), .o(n_15957) );
na02f80 g773534 ( .a(n_7477), .b(n_7276), .o(n_7488) );
in01f80 g750954 ( .a(n_28950), .o(n_28951) );
in01f80 g760503 ( .a(n_20002), .o(n_20024) );
no02f80 g779147 ( .a(n_1928), .b(n_1927), .o(n_1929) );
na02f80 g754803 ( .a(n_25458), .b(n_25455), .o(n_25459) );
in01f80 g744327 ( .a(n_35683), .o(n_35729) );
in01f80 FE_OCP_RBC1905_n_29080 ( .a(n_29080), .o(FE_OCP_RBN1905_n_29080) );
in01f80 fopt783135 ( .a(n_24862), .o(n_44621) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_15_ ( .ck(newNet_1025), .d(n_17855), .o(delay_xor_ln21_unr12_stage5_stallmux_q_15_) );
in01f80 FE_OCP_RBC2136_n_11907 ( .a(n_11907), .o(FE_OCP_RBN2136_n_11907) );
ao12f80 g756755 ( .a(n_23459), .b(n_23458), .c(n_23457), .o(n_24919) );
na02f80 g775676 ( .a(n_5565), .b(n_5589), .o(n_5620) );
no02f80 g773661 ( .a(n_7267), .b(n_7265), .o(n_7266) );
in01f80 newInst_2469 ( .a(newNet_2468), .o(newNet_2469) );
in01f80 newInst_1948 ( .a(newNet_1947), .o(newNet_1948) );
na02f80 g770952 ( .a(n_10027), .b(n_10164), .o(n_10288) );
ao22s80 FE_RC_3906_0 ( .a(n_20527), .b(FE_RN_422_0), .c(n_20526), .d(FE_OCP_RBN1725_FE_RN_422_0), .o(n_21004) );
ao12f80 g773844 ( .a(n_7128), .b(n_7127), .c(n_7126), .o(n_8050) );
in01f80 newInst_2811 ( .a(newNet_2412), .o(newNet_2811) );
na02f80 g767003 ( .a(n_14758), .b(n_14170), .o(n_14211) );
no02f80 g761142 ( .a(n_19797), .b(n_19714), .o(n_20115) );
na02f80 g754479 ( .a(n_26686), .b(n_26708), .o(n_26742) );
na02f80 g760068 ( .a(n_20482), .b(FE_OCP_RBN3617_n_20249), .o(n_20538) );
na02f80 g738588 ( .a(n_41400), .b(n_41449), .o(n_41520) );
na02f80 g765279 ( .a(n_15714), .b(n_15749), .o(n_15750) );
oa12f80 g770661 ( .a(n_9947), .b(n_10030), .c(n_9891), .o(n_10102) );
in01f80 newInst_656 ( .a(newNet_655), .o(newNet_656) );
in01f80 FE_OCP_RBC1709_n_22150 ( .a(FE_OCP_RBN1708_n_22150), .o(FE_OCP_RBN1709_n_22150) );
ao12f80 g778443 ( .a(n_2935), .b(n_2876), .c(n_3297), .o(n_3465) );
in01f80 FE_RC_4196_0 ( .a(FE_OCPUNCON3143_n_19138), .o(FE_RN_1839_0) );
oa12f80 g767248 ( .a(n_13525), .b(n_13568), .c(n_13608), .o(n_13623) );
na03f80 g778960 ( .a(n_1697), .b(n_2144), .c(n_1714), .o(n_2177) );
no02f80 g761649 ( .a(n_18601), .b(n_18316), .o(n_18683) );
no02f80 g742193 ( .a(n_44869), .b(n_37871), .o(n_37872) );
in01f80 g776117 ( .a(n_5150), .o(n_5224) );
na02f80 g765792 ( .a(n_14978), .b(n_14977), .o(n_15003) );
in01f80 newInst_939 ( .a(newNet_938), .o(newNet_939) );
in01f80 newInst_493 ( .a(newNet_492), .o(newNet_493) );
in01f80 g767891 ( .a(n_12925), .o(n_12926) );
na02f80 g749198 ( .a(n_30820), .b(n_27246), .o(n_30851) );
oa22f80 g778647 ( .a(FE_OCP_RBN2320_n_2382), .b(n_2070), .c(n_2382), .d(n_2071), .o(n_2484) );
in01f80 FE_OCPC1239_n_37945 ( .a(FE_OCP_RBN3443_n_37945), .o(FE_OCPN1239_n_37945) );
oa22f80 g748198 ( .a(FE_OCPN981_n_31961), .b(n_30299), .c(FE_OCPN880_n_31944), .d(n_30327), .o(n_32182) );
in01f80 newInst_704 ( .a(newNet_703), .o(newNet_704) );
no02f80 g751373 ( .a(n_29388), .b(n_28960), .o(n_29432) );
in01f80 g777158 ( .a(n_5258), .o(n_5259) );
in01f80 g769328 ( .a(n_11863), .o(n_11864) );
oa12f80 g764554 ( .a(n_16545), .b(n_16544), .c(n_16543), .o(n_16592) );
no02f80 g778524 ( .a(n_2546), .b(n_2521), .o(n_2566) );
na02f80 g740190 ( .a(FE_OCP_RBN3719_n_39913), .b(FE_OCP_RBN2834_n_39586), .o(n_40106) );
in01f80 FE_OCP_RBC2138_n_11909 ( .a(n_11909), .o(FE_OCP_RBN2138_n_11909) );
in01f80 g777898 ( .a(n_3176), .o(n_3135) );
no02f80 g754076 ( .a(n_26119), .b(n_26096), .o(n_26194) );
in01f80 newInst_201 ( .a(newNet_200), .o(newNet_201) );
ao22s80 FE_RC_476_0 ( .a(n_30466), .b(FE_OCP_RBN1296_n_30451), .c(n_27014), .d(n_30451), .o(n_30542) );
in01f80 newInst_2412 ( .a(newNet_2411), .o(newNet_2412) );
ao12f80 g752973 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_28109) );
ao12f80 g779811 ( .a(n_1632), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_11_), .o(n_1850) );
in01f80 g749746 ( .a(n_31573), .o(n_31574) );
ao12f80 g766296 ( .a(n_14702), .b(n_14701), .c(n_14700), .o(n_14779) );
in01f80 g768691 ( .a(n_12285), .o(n_12286) );
in01f80 drc784749 ( .a(n_30614), .o(n_30633) );
na02f80 g770671 ( .a(n_10373), .b(n_10351), .o(n_10352) );
na02f80 g769602 ( .a(n_11320), .b(FE_OCP_RBN2845_n_10326), .o(n_11392) );
no02f80 g738922 ( .a(n_41277), .b(n_41276), .o(n_41278) );
na02f80 FE_RC_2837_0 ( .a(FE_RN_1219_0), .b(FE_OCP_RBN3082_n_16977), .o(n_17130) );
in01f80 FE_OCP_RBC2770_n_9892 ( .a(n_9892), .o(FE_OCP_RBN2770_n_9892) );
in01f80 FE_RC_3101_0 ( .a(n_45073), .o(FE_RN_1371_0) );
in01f80 FE_OCP_RBC3470_n_7886 ( .a(FE_OCP_RBN3464_n_7886), .o(FE_OCP_RBN3470_n_7886) );
na02f80 g747431 ( .a(n_32368), .b(n_32433), .o(n_32472) );
na02f80 g772357 ( .a(n_8626), .b(n_8603), .o(n_8628) );
in01f80 g762939 ( .a(n_17523), .o(n_17595) );
no02f80 g776062 ( .a(n_4559), .b(n_4427), .o(n_4683) );
in01f80 newInst_1041 ( .a(newNet_1040), .o(newNet_1041) );
no02f80 g736584 ( .a(n_43657), .b(n_43464), .o(n_43658) );
na02f80 FE_RC_2312_0 ( .a(FE_RN_877_0), .b(n_34666), .o(FE_RN_878_0) );
ao12f80 g782651 ( .a(n_28836), .b(n_28883), .c(n_28690), .o(n_44045) );
no02f80 g750607 ( .a(FE_OCP_RBN2332_n_29380), .b(n_29328), .o(n_29422) );
in01f80 g780807 ( .a(n_1108), .o(n_419) );
in01f80 FE_OCPC3785_FE_OCP_RBN2831_n_10198 ( .a(FE_OCPN3784_FE_OCP_RBN2831_n_10198), .o(FE_OCPN3785_FE_OCP_RBN2831_n_10198) );
in01f80 g738467 ( .a(n_41470), .o(n_41471) );
no02f80 g759165 ( .a(n_21012), .b(n_20976), .o(n_21049) );
no02f80 g763824 ( .a(n_17355), .b(n_17263), .o(n_17818) );
in01f80 g768390 ( .a(n_12445), .o(n_12427) );
in01f80 g769422 ( .a(n_11440), .o(n_11627) );
no02f80 g747421 ( .a(n_32399), .b(n_44962), .o(n_32475) );
in01f80 g737035 ( .a(n_43048), .o(n_43067) );
no02f80 g751449 ( .a(n_28574), .b(delay_add_ln22_unr17_stage7_stallmux_q_23_), .o(n_28575) );
na02f80 g737387 ( .a(n_42775), .b(n_42628), .o(n_42795) );
no02f80 g777777 ( .a(n_3306), .b(n_3305), .o(n_3307) );
no02f80 g768285 ( .a(n_12644), .b(n_12372), .o(n_12675) );
no02f80 g773129 ( .a(n_7674), .b(n_7663), .o(n_7698) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_7_ ( .ck(newNet_289), .d(n_1285), .o(delay_xor_ln22_unr3_stage2_stallmux_q_7_) );
no02f80 g779628 ( .a(FE_OCP_RBN3246_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_4_), .o(n_1380) );
in01f80 newInst_203 ( .a(newNet_107), .o(newNet_203) );
no02f80 g778275 ( .a(n_47026), .b(n_2702), .o(n_2739) );
in01f80 fopt783239 ( .a(n_44798), .o(n_44797) );
in01f80 newInst_1172 ( .a(newNet_197), .o(newNet_1172) );
in01f80 FE_OCPC1474_n_24624 ( .a(FE_OCPN1473_n_24624), .o(FE_OCPN1474_n_24624) );
in01f80 FE_RC_639_0 ( .a(n_28460), .o(FE_RN_201_0) );
na02f80 g761734 ( .a(n_19339), .b(n_18965), .o(n_19338) );
na02f80 g740399 ( .a(FE_OCP_RBN3021_n_39942), .b(n_46949), .o(n_39995) );
no02f80 FE_RC_1041_0 ( .a(FE_RN_300_0), .b(FE_RN_301_0), .o(FE_RN_302_0) );
in01f80 newInst_2876 ( .a(newNet_2875), .o(newNet_2876) );
no02f80 g743100 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_26_), .o(n_37100) );
in01f80 g741562 ( .a(n_38676), .o(n_38677) );
no02f80 g756852 ( .a(n_23404), .b(n_23403), .o(n_23418) );
oa12f80 g762311 ( .a(n_18001), .b(n_17971), .c(n_18052), .o(n_18059) );
no02f80 g756194 ( .a(n_24164), .b(n_24162), .o(n_24163) );
in01f80 g769835 ( .a(n_11166), .o(n_11228) );
na02f80 g776245 ( .a(n_4319), .b(n_4263), .o(n_4338) );
in01f80 newInst_1090 ( .a(newNet_1089), .o(newNet_1090) );
no02f80 g744061 ( .a(n_44223), .b(n_35824), .o(n_36293) );
in01f80 FE_OCP_RBC3689_n_16146 ( .a(n_16146), .o(FE_OCP_RBN3689_n_16146) );
oa12f80 g759675 ( .a(n_21334), .b(n_21337), .c(n_21406), .o(n_21452) );
no02f80 g746005 ( .a(n_34010), .b(n_34009), .o(n_34030) );
na02f80 FE_RC_4017_0 ( .a(FE_RN_1744_0), .b(n_15427), .o(n_15468) );
in01f80 g756330 ( .a(n_24588), .o(n_24542) );
no02f80 g775673 ( .a(n_5455), .b(n_5405), .o(n_5406) );
in01f80 g772051 ( .a(n_47244), .o(n_8950) );
ao12f80 g741486 ( .a(n_38737), .b(n_38747), .c(n_38736), .o(n_38767) );
in01f80 FE_RC_3352_0 ( .a(n_21067), .o(FE_RN_1462_0) );
no02f80 g767552 ( .a(n_13306), .b(n_13305), .o(n_13307) );
in01f80 FE_OCPC1475_n_23708 ( .a(n_23708), .o(FE_OCPN1475_n_23708) );
in01f80 g755350 ( .a(n_24810), .o(n_24840) );
in01f80 g773223 ( .a(n_8676), .o(n_7635) );
in01f80 fopt783244 ( .a(n_44800), .o(n_44804) );
na02f80 FE_RC_2544_0 ( .a(n_38904), .b(n_38959), .o(FE_RN_1041_0) );
na02f80 g748431 ( .a(n_31466), .b(n_30954), .o(n_31682) );
in01f80 g768512 ( .a(n_12412), .o(n_12366) );
no02f80 FE_RC_1735_0 ( .a(n_37003), .b(n_37014), .o(FE_RN_483_0) );
na02f80 g762969 ( .a(n_17623), .b(n_17672), .o(n_17746) );
in01f80 newInst_1406 ( .a(newNet_735), .o(newNet_1406) );
na02f80 g773681 ( .a(n_7933), .b(n_7795), .o(n_7407) );
no02f80 g754090 ( .a(n_26097), .b(n_23466), .o(n_26156) );
ao12f80 g739026 ( .a(n_41136), .b(n_41135), .c(n_41134), .o(n_41473) );
na02f80 g745293 ( .a(n_35891), .b(n_35890), .o(n_35935) );
no02f80 g756732 ( .a(n_23426), .b(n_23142), .o(n_23478) );
na02f80 g772257 ( .a(n_8579), .b(n_8578), .o(n_8641) );
na02f80 g768925 ( .a(n_12213), .b(n_12168), .o(n_12214) );
in01f80 g763834 ( .a(n_16684), .o(n_16685) );
na02f80 g737731 ( .a(n_42392), .b(n_42117), .o(n_42522) );
no02f80 g755141 ( .a(n_25551), .b(n_25104), .o(n_25693) );
in01f80 FE_OFC790_n_8981 ( .a(n_8981), .o(FE_OFN790_n_8981) );
na02f80 g772235 ( .a(n_8727), .b(n_8104), .o(n_8761) );
no02f80 g743003 ( .a(n_37094), .b(n_37109), .o(n_37357) );
no02f80 g752801 ( .a(n_28076), .b(n_27853), .o(n_28585) );
in01f80 FE_OCP_RBC1181_n_19726 ( .a(n_19726), .o(FE_OCP_RBN1181_n_19726) );
na02f80 g778144 ( .a(n_2956), .b(n_2903), .o(n_2983) );
in01f80 FE_OCP_RBC3390_n_33108 ( .a(FE_OCP_RBN3388_n_33108), .o(FE_OCP_RBN3390_n_33108) );
in01f80 g776182 ( .a(n_4966), .o(n_5035) );
oa12f80 g749229 ( .a(n_31418), .b(n_32094), .c(n_31313), .o(n_32158) );
in01f80 newInst_2561 ( .a(newNet_2560), .o(newNet_2561) );
in01f80 newInst_1082 ( .a(newNet_734), .o(newNet_1082) );
in01f80 FE_OCP_RBC2374_n_8221 ( .a(FE_OCP_RBN2372_n_8221), .o(FE_OCP_RBN2374_n_8221) );
ao22s80 FE_RC_802_0 ( .a(FE_OCP_RBN2304_n_7817), .b(n_8637), .c(n_8612), .d(FE_OCP_RBN3474_n_7886), .o(n_8790) );
in01f80 g742106 ( .a(n_38010), .o(n_37907) );
no02f80 g758333 ( .a(n_22187), .b(n_22251), .o(n_22291) );
no02f80 g753096 ( .a(n_27119), .b(n_27117), .o(n_27154) );
no02f80 g747720 ( .a(n_32088), .b(n_32086), .o(n_32087) );
in01f80 g770091 ( .a(n_11015), .o(n_11016) );
in01f80 g768762 ( .a(n_12223), .o(n_12224) );
no02f80 g765501 ( .a(n_15599), .b(n_15712), .o(n_15928) );
no02f80 g738729 ( .a(n_41483), .b(n_41484), .o(n_41828) );
na02f80 g759899 ( .a(n_21374), .b(n_20895), .o(n_21598) );
in01f80 newInst_2789 ( .a(newNet_1167), .o(newNet_2789) );
na02f80 g747300 ( .a(n_33630), .b(n_33629), .o(n_33631) );
ms00f80 delay_sub_ln23_0_unr21_stage8_stallmux_q_reg ( .ck(newNet_1555), .d(n_28897), .o(delay_sub_ln23_0_unr21_stage8_stallmux_q) );
ao12f80 g738235 ( .a(n_41929), .b(n_41928), .c(n_41927), .o(n_41956) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_26_ ( .ck(newNet_3516), .d(n_22819), .o(delay_add_ln22_unr14_stage6_stallmux_q_26_) );
na02f80 g751585 ( .a(n_28440), .b(n_28465), .o(n_28486) );
oa12f80 g760585 ( .a(n_19531), .b(n_19860), .c(n_19451), .o(n_19861) );
in01f80 g766576 ( .a(n_13992), .o(n_14190) );
ao12f80 g763856 ( .a(n_17360), .b(n_17256), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_13_), .o(n_18033) );
in01f80 FE_OCP_DRV_C1608_n_31473 ( .a(FE_OCP_DRV_N1607_n_31473), .o(FE_OCP_DRV_N1608_n_31473) );
in01f80 g752164 ( .a(n_28664), .o(n_28665) );
in01f80 FE_RC_3184_0 ( .a(n_6715), .o(FE_RN_1413_0) );
na02f80 g753809 ( .a(n_26329), .b(n_26245), .o(n_26374) );
no02f80 g747336 ( .a(n_33863), .b(n_33862), .o(n_33864) );
in01f80 newInst_1303 ( .a(newNet_1302), .o(newNet_1303) );
in01f80 FE_RC_439_0 ( .a(FE_RN_125_0), .o(n_17601) );
in01f80 g765106 ( .a(n_16259), .o(n_16260) );
oa12f80 g770915 ( .a(n_10087), .b(n_10131), .c(n_10086), .o(n_10168) );
in01f80 FE_OFC821_n_4632 ( .a(FE_OFN838_n_4632), .o(FE_OFN821_n_4632) );
na02f80 g776259 ( .a(n_4547), .b(n_4638), .o(n_4782) );
in01f80 g765196 ( .a(n_16131), .o(n_16132) );
in01f80 newInst_1078 ( .a(newNet_1077), .o(newNet_1078) );
in01f80 g747234 ( .a(n_33588), .o(n_33689) );
na02f80 g778258 ( .a(n_2677), .b(n_2646), .o(n_2795) );
na02f80 g751014 ( .a(n_30159), .b(n_30093), .o(n_30160) );
in01f80 g758948 ( .a(n_21676), .o(n_21677) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_20_ ( .ck(newNet_2754), .d(n_17440), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_20_) );
no02f80 g738266 ( .a(n_41891), .b(n_41890), .o(n_41892) );
oa12f80 g742856 ( .a(n_37250), .b(n_37249), .c(n_37248), .o(n_37877) );
na02f80 g757254 ( .a(n_23136), .b(n_23135), .o(n_23214) );
no02f80 g744981 ( .a(n_34828), .b(n_30588), .o(n_34862) );
in01f80 FE_OCP_RBC2363_n_13785 ( .a(n_13785), .o(FE_OCP_RBN2363_n_13785) );
in01f80 newInst_2202 ( .a(newNet_2201), .o(newNet_2202) );
in01f80 g741680 ( .a(n_38568), .o(n_39025) );
no02f80 g773410 ( .a(n_7584), .b(n_7651), .o(n_7671) );
in01f80 g779776 ( .a(n_1396), .o(n_1443) );
in01f80 g778505 ( .a(n_2558), .o(n_2828) );
in01f80 newInst_3116 ( .a(newNet_710), .o(newNet_3116) );
in01f80 newInst_2373 ( .a(newNet_133), .o(newNet_2373) );
in01f80 g779114 ( .a(n_2066), .o(n_2523) );
oa12f80 g749001 ( .a(n_31005), .b(n_31004), .c(n_31003), .o(n_31051) );
in01f80 g780960 ( .a(n_420), .o(n_521) );
ao12f80 g780134 ( .a(n_711), .b(n_948), .c(n_727), .o(n_1029) );
in01f80 g747449 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_27_), .o(n_32355) );
no02f80 g780529 ( .a(n_682), .b(n_673), .o(n_686) );
no02f80 g744892 ( .a(n_35077), .b(n_30587), .o(n_35134) );
oa12f80 g761685 ( .a(n_18243), .b(n_18647), .c(n_18221), .o(n_18756) );
in01f80 FE_RC_2864_0 ( .a(n_34560), .o(FE_RN_1234_0) );
in01f80 FE_RC_3254_0 ( .a(n_11500), .o(FE_RN_1436_0) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_30_ ( .ck(newNet_2823), .d(n_12211), .o(delay_add_ln22_unr8_stage4_stallmux_q_30_) );
ao12f80 g774232 ( .a(n_6560), .b(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .c(delay_xor_ln21_unr6_stage3_stallmux_q_6_), .o(n_6596) );
na02f80 FE_RC_3013_0 ( .a(FE_RN_1320_0), .b(n_15768), .o(FE_RN_1321_0) );
na02f80 g752590 ( .a(n_27573), .b(n_27512), .o(n_27602) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_17_ ( .ck(newNet_2010), .d(n_11369), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_17_) );
in01f80 g765943 ( .a(n_14792), .o(n_14793) );
oa12f80 g768508 ( .a(n_12371), .b(n_12327), .c(FE_OCPN1002_n_45660), .o(n_12570) );
no02f80 g743435 ( .a(n_36552), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36587) );
in01f80 g739064 ( .a(n_41073), .o(n_41119) );
na02f80 g771006 ( .a(n_10070), .b(n_10204), .o(n_10302) );
in01f80 g749345 ( .a(n_30824), .o(n_30792) );
in01f80 g766465 ( .a(n_14176), .o(n_14225) );
in01f80 g749823 ( .a(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36750) );
ao22s80 g778306 ( .a(n_2558), .b(FE_OCPN1234_n_2414), .c(n_2664), .d(FE_OCPN1234_n_2414), .o(n_2673) );
na02f80 g780033 ( .a(n_1248), .b(n_1053), .o(n_1255) );
na02f80 g747577 ( .a(n_33361), .b(n_33362), .o(n_33363) );
na02f80 g766823 ( .a(n_14381), .b(n_14297), .o(n_14382) );
ao12f80 g769392 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_8_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_7_), .o(n_11890) );
ao12f80 g749092 ( .a(FE_OCPN1490_n_30823), .b(n_30910), .c(n_30824), .o(n_30961) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_27_ ( .ck(newNet_3608), .d(n_17811), .o(delay_add_ln22_unr11_stage5_stallmux_q_27_) );
no02f80 g741781 ( .a(n_38400), .b(n_38399), .o(n_38401) );
oa12f80 g746995 ( .a(n_34023), .b(n_34022), .c(n_34021), .o(n_34613) );
no02f80 g758748 ( .a(n_21615), .b(n_21505), .o(n_21664) );
in01f80 newInst_3193 ( .a(newNet_3192), .o(newNet_3193) );
na02f80 g767239 ( .a(n_13535), .b(n_13530), .o(n_13536) );
na02f80 g777717 ( .a(n_3337), .b(n_3358), .o(n_3645) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_25_ ( .ck(newNet_2175), .d(n_1048), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_25_) );
no02f80 g738822 ( .a(n_41324), .b(n_41343), .o(n_41430) );
in01f80 FE_OCP_RBC3043_n_46337 ( .a(FE_OCP_RBN3040_n_46337), .o(FE_OCP_RBN3043_n_46337) );
no02f80 g772500 ( .a(n_8374), .b(n_45827), .o(n_8443) );
oa22f80 g765403 ( .a(n_15874), .b(n_15482), .c(n_16245), .d(n_15513), .o(n_16342) );
oa12f80 g760810 ( .a(n_20122), .b(n_20121), .c(n_20120), .o(n_20180) );
in01f80 fopt783398 ( .a(n_23525), .o(n_44996) );
in01f80 newInst_770 ( .a(newNet_680), .o(newNet_770) );
oa12f80 g737630 ( .a(n_42540), .b(FE_OCPN887_n_42367), .c(n_41909), .o(n_42644) );
in01f80 newInst_1390 ( .a(newNet_1341), .o(newNet_1390) );
ao12f80 g746515 ( .a(n_34666), .b(n_34776), .c(n_34738), .o(n_34812) );
in01f80 FE_OCP_RBC2271_n_13489 ( .a(n_13489), .o(FE_OCP_RBN2271_n_13489) );
oa12f80 g782635 ( .a(n_44610), .b(FE_OCP_RBN3356_delay_xor_ln22_unr28_stage10_stallmux_q_0_), .c(n_40604), .o(n_44028) );
in01f80 FE_RC_2989_0 ( .a(n_9979), .o(FE_RN_1305_0) );
na02f80 FE_RC_2766_0 ( .a(FE_RN_1178_0), .b(n_33957), .o(n_33977) );
no02f80 g747815 ( .a(n_33226), .b(n_33240), .o(n_33241) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_8_ ( .ck(newNet_3094), .d(n_40428), .o(delay_add_ln22_unr27_stage10_stallmux_q_8_) );
in01f80 FE_RC_2506_0 ( .a(n_17845), .o(FE_RN_1018_0) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_11_ ( .ck(newNet_2026), .d(n_10848), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_11_) );
na02f80 g739298 ( .a(n_40766), .b(n_40508), .o(n_40767) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_28_ ( .ck(newNet_1973), .d(n_12114), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_28_) );
in01f80 FE_RC_2804_0 ( .a(n_25301), .o(FE_RN_1200_0) );
na02f80 g740862 ( .a(n_39377), .b(n_38978), .o(n_39436) );
na02f80 g756349 ( .a(n_24066), .b(n_23966), .o(n_24092) );
in01f80 g738800 ( .a(n_41456), .o(n_41491) );
in01f80 FE_OCP_RBC1338_n_20941 ( .a(FE_OCP_RBN1337_n_20941), .o(FE_OCP_RBN1338_n_20941) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_13_ ( .ck(newNet_2970), .d(n_5840), .o(delay_add_ln22_unr5_stage3_stallmux_q_13_) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_3_ ( .ck(newNet_3111), .d(n_39896), .o(delay_add_ln22_unr27_stage10_stallmux_q_3_) );
in01f80 g752337 ( .a(n_27911), .o(n_28095) );
no02f80 g767352 ( .a(n_13433), .b(n_13453), .o(n_13454) );
no02f80 FE_RC_472_0 ( .a(n_28568), .b(FE_RN_139_0), .o(FE_RN_140_0) );
ao12f80 g778453 ( .a(n_2398), .b(n_2397), .c(n_2396), .o(n_3771) );
ao12f80 g747168 ( .a(n_33894), .b(n_33893), .c(n_33892), .o(n_34580) );
in01f80 g778984 ( .a(n_2214), .o(n_2257) );
in01f80 g748442 ( .a(n_31784), .o(n_31785) );
na02f80 g776104 ( .a(n_4906), .b(n_4905), .o(n_5026) );
no02f80 g736713 ( .a(n_43267), .b(FE_OCP_RBN3067_n_43230), .o(n_43364) );
na02f80 g772529 ( .a(n_8569), .b(n_8568), .o(n_8590) );
na02f80 FE_RC_1851_0 ( .a(n_44962), .b(FE_RN_564_0), .o(n_32632) );
oa12f80 g778020 ( .a(n_2856), .b(n_3020), .c(n_3034), .o(n_3090) );
na02f80 g758317 ( .a(n_22288), .b(n_21282), .o(n_22399) );
oa22f80 g751524 ( .a(FE_OCP_RBN3407_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .c(FE_OCP_RBN2215_FE_OCPN950_n_28595), .d(n_27806), .o(n_28847) );
na02f80 g740107 ( .a(n_40074), .b(n_40180), .o(n_40281) );
in01f80 g753530 ( .a(n_26837), .o(n_26838) );
in01f80 newInst_3477 ( .a(newNet_3476), .o(newNet_3477) );
in01f80 fopt784710 ( .a(n_21558), .o(n_47187) );
no02f80 g761154 ( .a(n_19912), .b(n_19845), .o(n_20016) );
in01f80 newInst_2100 ( .a(newNet_2099), .o(newNet_2100) );
no02f80 g757264 ( .a(n_23450), .b(n_23058), .o(n_23490) );
na02f80 g775006 ( .a(n_6132), .b(n_6131), .o(n_6148) );
in01f80 g758282 ( .a(n_22018), .o(n_22019) );
na02f80 g766735 ( .a(n_13726), .b(FE_OCPN860_n_12880), .o(n_13727) );
in01f80 g747387 ( .a(n_32572), .o(n_32573) );
na02f80 g740038 ( .a(n_39846), .b(n_39844), .o(n_39871) );
in01f80 newInst_2079 ( .a(newNet_2078), .o(newNet_2079) );
na02f80 g772206 ( .a(n_8641), .b(n_8633), .o(n_8739) );
in01f80 newInst_2891 ( .a(newNet_2890), .o(newNet_2891) );
na02f80 g773029 ( .a(n_7692), .b(n_7728), .o(n_7729) );
ao12f80 g748755 ( .a(n_30708), .b(n_31241), .c(n_31027), .o(n_31243) );
ao12f80 g757870 ( .a(n_23026), .b(n_22841), .c(n_22725), .o(n_23085) );
na02f80 g779054 ( .a(n_2043), .b(n_1900), .o(n_2044) );
in01f80 g736475 ( .a(n_43750), .o(n_43751) );
in01f80 g761041 ( .a(n_19565), .o(n_19313) );
no02f80 g759947 ( .a(n_21374), .b(n_21593), .o(n_21748) );
no02f80 g757553 ( .a(FE_OCP_RBN3821_n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_3_), .o(n_22823) );
in01f80 newInst_1426 ( .a(newNet_673), .o(newNet_1426) );
na02f80 g756938 ( .a(n_23722), .b(n_23863), .o(n_23723) );
na02f80 g768942 ( .a(FE_OCPN3188_n_11012), .b(n_11698), .o(n_11699) );
in01f80 FE_RC_792_0 ( .a(n_41425), .o(FE_RN_240_0) );
in01f80 FE_OCP_RBC2264_n_29033 ( .a(FE_OCP_RBN2263_n_29033), .o(FE_OCP_RBN2264_n_29033) );
in01f80 FE_OCP_RBC2570_n_29922 ( .a(n_29857), .o(FE_OCP_RBN2570_n_29922) );
in01f80 FE_OCP_DRV_C3745_FE_OFN737_n_22641 ( .a(FE_OCP_DRV_N3744_FE_OFN737_n_22641), .o(FE_OCP_DRV_N3745_FE_OFN737_n_22641) );
na02f80 g763915 ( .a(n_17054), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_4_), .o(n_17159) );
no02f80 g740979 ( .a(n_38933), .b(n_38882), .o(n_39086) );
oa12f80 FE_RC_2536_0 ( .a(FE_RN_1034_0), .b(n_36490), .c(n_36234), .o(n_36567) );
no02f80 g779762 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_), .o(n_1749) );
oa12f80 g764901 ( .a(n_15754), .b(n_15753), .c(n_15752), .o(n_15842) );
in01f80 newInst_3580 ( .a(newNet_3579), .o(newNet_3580) );
oa22f80 g776075 ( .a(n_5048), .b(n_5422), .c(n_44862), .d(FE_OCP_RBN2700_n_4238), .o(n_5056) );
ao12f80 g773888 ( .a(n_7057), .b(n_7094), .c(n_7056), .o(n_7769) );
na02f80 g762790 ( .a(n_17942), .b(delay_add_ln22_unr11_stage5_stallmux_q_10_), .o(n_18015) );
no02f80 g781107 ( .a(n_257), .b(n_264), .o(n_265) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_23_ ( .ck(newNet_2092), .d(n_6476), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_) );
no02f80 g768427 ( .a(n_12453), .b(n_12452), .o(n_12475) );
in01f80 FE_OCP_RBC3404_n_28597 ( .a(FE_OCP_RBN2192_n_28597), .o(FE_OCP_RBN3404_n_28597) );
na02f80 g745153 ( .a(n_34604), .b(n_34603), .o(n_34605) );
in01f80 FE_OCP_RBC3221_n_22068 ( .a(FE_OCP_RBN1847_n_22068), .o(FE_OCP_RBN3221_n_22068) );
na03f80 FE_RC_1153_0 ( .a(n_37156), .b(n_37488), .c(n_37337), .o(n_37536) );
oa12f80 g777669 ( .a(n_3368), .b(n_3407), .c(n_2759), .o(n_3478) );
no02f80 g761451 ( .a(n_20086), .b(n_19873), .o(n_20084) );
na02f80 g774801 ( .a(n_45479), .b(n_6263), .o(n_6299) );
oa22f80 g752752 ( .a(n_27077), .b(n_27037), .c(n_27076), .d(n_27038), .o(n_27129) );
na02f80 g767990 ( .a(n_12813), .b(n_12841), .o(n_13215) );
in01f80 newInst_2164 ( .a(newNet_2163), .o(newNet_2164) );
in01f80 g761244 ( .a(n_19131), .o(n_19345) );
in01f80 g764271 ( .a(n_16434), .o(n_16435) );
no02f80 g765893 ( .a(n_15092), .b(n_14968), .o(n_14969) );
no02f80 g778273 ( .a(n_2642), .b(n_2294), .o(n_2704) );
na02f80 g743142 ( .a(n_37033), .b(n_37032), .o(n_37085) );
na02f80 g741297 ( .a(FE_OCP_RBN2549_n_44944), .b(n_38829), .o(n_38906) );
in01f80 FE_OCP_RBC3454_FE_OCPN1240_n_7721 ( .a(FE_OCP_RBN3453_FE_OCPN1240_n_7721), .o(FE_OCP_RBN3454_FE_OCPN1240_n_7721) );
na02f80 g736958 ( .a(FE_OCPN912_n_43022), .b(n_42922), .o(n_43254) );
na02f80 g778037 ( .a(n_2969), .b(n_3013), .o(n_2970) );
na02f80 g776905 ( .a(n_3811), .b(n_3843), .o(n_3847) );
ao12f80 g774097 ( .a(n_6967), .b(n_6966), .c(n_6965), .o(n_7663) );
na02f80 g775089 ( .a(n_6034), .b(n_4903), .o(n_6086) );
in01f80 g753464 ( .a(n_26808), .o(n_26809) );
na03f80 g750810 ( .a(n_29036), .b(n_29039), .c(n_28703), .o(n_29065) );
in01f80 g751056 ( .a(n_30061), .o(n_30164) );
no02f80 g761541 ( .a(n_19548), .b(n_19547), .o(n_19549) );
na02f80 g740174 ( .a(FE_OCP_RBN3719_n_39913), .b(n_40011), .o(n_40180) );
na02f80 g755183 ( .a(n_25145), .b(n_25144), .o(n_25146) );
in01f80 FE_OCP_RBC2920_n_31107 ( .a(n_31107), .o(FE_OCP_RBN2920_n_31107) );
in01f80 g755967 ( .a(n_29561), .o(n_29630) );
no02f80 g745527 ( .a(n_34377), .b(n_34319), .o(n_34709) );
na02f80 g754448 ( .a(n_25654), .b(n_25296), .o(n_25676) );
in01f80 FE_OCPC3169_n_23227 ( .a(n_23227), .o(FE_OCPN3169_n_23227) );
in01f80 g758255 ( .a(n_22647), .o(n_22648) );
in01f80 g768802 ( .a(n_12207), .o(n_12208) );
na02f80 g751834 ( .a(n_28255), .b(n_28224), .o(n_28225) );
no02f80 g776627 ( .a(n_3964), .b(n_3106), .o(n_4166) );
no02f80 g755573 ( .a(n_24646), .b(n_24645), .o(n_24647) );
na02f80 g775589 ( .a(n_5783), .b(n_5658), .o(n_5784) );
no02f80 g759634 ( .a(n_20727), .b(n_45067), .o(n_20756) );
in01f80 g744084 ( .a(n_35622), .o(n_35623) );
in01f80 g762087 ( .a(n_18541), .o(n_18455) );
in01f80 newInst_3122 ( .a(newNet_3121), .o(newNet_3122) );
no02f80 g769030 ( .a(n_45659), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_), .o(n_12278) );
in01f80 FE_OCP_RBC3342_delay_add_ln22_unr23_stage9_stallmux_q_24_ ( .a(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(FE_OCP_RBN3342_delay_add_ln22_unr23_stage9_stallmux_q_24_) );
no02f80 g746008 ( .a(n_33908), .b(n_33907), .o(n_33923) );
na02f80 g761027 ( .a(n_19244), .b(n_17837), .o(n_19348) );
in01f80 g738149 ( .a(n_42071), .o(n_42037) );
na02f80 g752233 ( .a(n_27869), .b(n_44735), .o(n_27971) );
in01f80 g774488 ( .a(n_6683), .o(n_6623) );
in01f80 g744216 ( .a(n_36186), .o(n_36187) );
no02f80 g742433 ( .a(n_37610), .b(n_37117), .o(n_37650) );
in01f80 FE_OCP_RBC2285_n_2433 ( .a(n_2433), .o(FE_OCP_RBN2285_n_2433) );
no02f80 g760363 ( .a(n_20160), .b(n_20170), .o(n_20171) );
in01f80 g742712 ( .a(n_37454), .o(n_37455) );
ao12f80 g763125 ( .a(n_17399), .b(n_17433), .c(n_17477), .o(n_17635) );
oa22f80 g747776 ( .a(n_33571), .b(n_33240), .c(n_33372), .d(n_33256), .o(n_34071) );
na02f80 g756446 ( .a(n_23686), .b(n_23599), .o(n_23737) );
na02f80 g744018 ( .a(n_36882), .b(n_36838), .o(n_36901) );
in01f80 newInst_192 ( .a(newNet_191), .o(newNet_192) );
na02f80 g780382 ( .a(n_715), .b(n_714), .o(n_716) );
in01f80 FE_OCP_RBC1986_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1986_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
na02f80 FE_RC_1676_0 ( .a(FE_RN_465_0), .b(FE_RN_466_0), .o(FE_RN_467_0) );
na02f80 g740789 ( .a(n_39431), .b(n_39391), .o(n_39472) );
in01f80 FE_RC_2984_0 ( .a(FE_RN_1303_0), .o(n_10953) );
in01f80 newInst_352 ( .a(newNet_351), .o(newNet_352) );
in01f80 g754688 ( .a(n_26486), .o(n_26862) );
in01f80 g765057 ( .a(n_15385), .o(n_15423) );
ao12f80 g751934 ( .a(n_28752), .b(n_28751), .c(n_28750), .o(n_29123) );
in01f80 g756304 ( .a(n_24606), .o(n_24607) );
in01f80 g750165 ( .a(n_29795), .o(n_29796) );
in01f80 g764804 ( .a(n_15700), .o(n_15708) );
na02f80 g746133 ( .a(n_33775), .b(n_33774), .o(n_33776) );
oa22f80 g743737 ( .a(n_36339), .b(n_36361), .c(n_36338), .d(n_36362), .o(n_36422) );
oa22f80 g737658 ( .a(FE_OCPN888_n_42367), .b(n_42066), .c(n_42392), .d(n_42048), .o(n_42756) );
in01f80 FE_OCPUNCOC1801_n_29375 ( .a(n_29375), .o(FE_OCPUNCON1801_n_29375) );
in01f80 g751548 ( .a(n_28468), .o(n_28469) );
na02f80 g760621 ( .a(n_19856), .b(FE_OCPN1436_n_19855), .o(n_19941) );
na02f80 g755414 ( .a(n_24755), .b(FE_OCPN1482_n_22207), .o(n_24829) );
na02f80 g745703 ( .a(n_35433), .b(n_34865), .o(n_35453) );
in01f80 g769745 ( .a(n_11209), .o(n_11247) );
in01f80 FE_OCP_RBC3826_n_18951 ( .a(n_18951), .o(FE_OCP_RBN3826_n_18951) );
oa22f80 g737648 ( .a(FE_OCPN888_n_42367), .b(n_41936), .c(n_42392), .d(n_42358), .o(n_42681) );
in01f80 newInst_1109 ( .a(newNet_1108), .o(newNet_1109) );
na02f80 g769649 ( .a(n_11317), .b(n_11345), .o(n_11366) );
ao12f80 g766688 ( .a(n_13124), .b(n_13778), .c(n_13777), .o(n_13812) );
na02f80 g780292 ( .a(n_1046), .b(n_1203), .o(n_1080) );
in01f80 g771982 ( .a(n_9649), .o(n_9650) );
no02f80 g749077 ( .a(n_30878), .b(n_30942), .o(n_31004) );
na02f80 g743513 ( .a(n_37699), .b(n_36826), .o(n_37711) );
in01f80 g751798 ( .a(n_28930), .o(n_28931) );
na02f80 g778555 ( .a(n_2335), .b(n_2238), .o(n_2392) );
no02f80 g765975 ( .a(n_13577), .b(n_14770), .o(n_14789) );
in01f80 newInst_1512 ( .a(newNet_177), .o(newNet_1512) );
no02f80 g738288 ( .a(n_41842), .b(n_41841), .o(n_41843) );
in01f80 FE_OCP_RBC2831_n_10198 ( .a(n_10198), .o(FE_OCP_RBN2831_n_10198) );
no02f80 g784405 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_17_), .o(n_46217) );
in01f80 newInst_1457 ( .a(newNet_889), .o(newNet_1457) );
na02f80 g737548 ( .a(n_42492), .b(n_42471), .o(n_42506) );
no02f80 g771763 ( .a(n_9110), .b(FE_OCP_RBN3552_n_44575), .o(n_9129) );
na02f80 g763868 ( .a(n_16642), .b(n_16663), .o(n_16757) );
no02f80 g770515 ( .a(n_10197), .b(n_10228), .o(n_10317) );
na02f80 g746697 ( .a(n_34330), .b(n_34329), .o(n_34331) );
na02f80 g771846 ( .a(n_44511), .b(n_10122), .o(n_10209) );
na02f80 g751490 ( .a(n_28508), .b(n_28495), .o(n_29011) );
na02f80 g751796 ( .a(n_28253), .b(n_28284), .o(n_28406) );
in01f80 g740332 ( .a(n_40392), .o(n_40393) );
no02f80 g736843 ( .a(n_43026), .b(n_43025), .o(n_43027) );
no02f80 g756824 ( .a(n_24029), .b(n_23987), .o(n_24030) );
na02f80 g764875 ( .a(n_16353), .b(n_16352), .o(n_16354) );
no02f80 g747797 ( .a(n_33226), .b(n_33281), .o(n_33317) );
no02f80 g751396 ( .a(n_29363), .b(n_28992), .o(n_29388) );
in01f80 g772587 ( .a(n_8511), .o(n_8512) );
in01f80 g764380 ( .a(n_16388), .o(n_16389) );
na02f80 g779357 ( .a(n_1592), .b(n_1560), .o(n_1638) );
no02f80 g740327 ( .a(n_40246), .b(n_39939), .o(n_40359) );
no02f80 g752186 ( .a(FE_OCP_RBN2126_n_44734), .b(delay_xor_ln21_unr18_stage7_stallmux_q_11_), .o(n_28039) );
in01f80 g765953 ( .a(n_14771), .o(n_14790) );
na02f80 g755821 ( .a(n_24396), .b(n_24017), .o(n_24423) );
na03f80 FE_RC_2995_0 ( .a(n_6412), .b(n_6535), .c(n_6447), .o(FE_RN_1309_0) );
in01f80 FE_OCPC1487_n_23447 ( .a(n_23447), .o(FE_OCPN1487_n_23447) );
na02f80 g773862 ( .a(n_7023), .b(delay_add_ln22_unr5_stage3_stallmux_q_10_), .o(n_7093) );
in01f80 g775479 ( .a(n_5614), .o(n_5640) );
na02f80 g750552 ( .a(n_29418), .b(n_29231), .o(n_29453) );
oa12f80 g743442 ( .a(n_37729), .b(n_37728), .c(n_37727), .o(n_37784) );
oa12f80 g780938 ( .a(n_374), .b(n_384), .c(n_516), .o(n_408) );
no02f80 g761210 ( .a(n_19015), .b(n_18280), .o(n_19059) );
in01f80 FE_OCP_RBC1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1983_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
no03m80 FE_RC_3741_0 ( .a(n_17036), .b(n_17137), .c(n_17027), .o(FE_RN_1400_0) );
na02f80 g749070 ( .a(n_30954), .b(n_27246), .o(n_30994) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_3_ ( .ck(newNet_449), .d(n_27700), .o(delay_xor_ln22_unr18_stage7_stallmux_q_3_) );
in01f80 g762101 ( .a(n_18195), .o(n_18226) );
na02f80 g762232 ( .a(n_18135), .b(n_17946), .o(n_18148) );
no02f80 g758885 ( .a(n_21365), .b(n_21397), .o(n_21438) );
no03m80 FE_RC_4214_0 ( .a(n_20125), .b(FE_OCP_RBN3844_FE_RN_1242_0), .c(n_20290), .o(n_20292) );
in01f80 FE_OCP_RBC2646_n_47015 ( .a(n_47015), .o(FE_OCP_RBN2646_n_47015) );
in01f80 newInst_483 ( .a(newNet_482), .o(newNet_483) );
na02f80 g741985 ( .a(n_37984), .b(n_37983), .o(n_37985) );
na02f80 g778652 ( .a(n_2380), .b(n_2379), .o(n_3317) );
ao22s80 FE_RC_3068_0 ( .a(n_45013), .b(FE_OCP_RBN1714_n_20734), .c(n_45050), .d(n_20734), .o(n_20857) );
no02f80 g777698 ( .a(n_3503), .b(FE_OCP_RBN2382_n_3502), .o(n_3535) );
in01f80 newInst_871 ( .a(newNet_745), .o(newNet_871) );
oa12f80 g759733 ( .a(FE_OCP_RBN3678_n_21051), .b(n_21482), .c(n_21481), .o(n_21483) );
in01f80 FE_OCP_RBC3476_n_7886 ( .a(FE_OCP_RBN3471_n_7886), .o(FE_OCP_RBN3476_n_7886) );
na02f80 g767965 ( .a(n_12832), .b(n_12815), .o(n_13018) );
in01f80 newInst_3497 ( .a(newNet_3496), .o(newNet_3497) );
in01f80 newInst_1979 ( .a(newNet_147), .o(newNet_1979) );
in01f80 g766309 ( .a(n_14370), .o(n_14371) );
in01f80 g780923 ( .a(n_530), .o(n_531) );
ao12f80 g773825 ( .a(n_7066), .b(n_7065), .c(n_7064), .o(n_7136) );
in01f80 FE_OCP_RBC2822_n_10023 ( .a(n_10023), .o(FE_OCP_RBN2822_n_10023) );
in01f80 newInst_2099 ( .a(newNet_1360), .o(newNet_2099) );
na02f80 g759993 ( .a(n_20291), .b(n_20267), .o(n_20379) );
in01f80 g757659 ( .a(n_22672), .o(n_22673) );
ao12f80 g760528 ( .a(n_20425), .b(n_20450), .c(n_20424), .o(n_21405) );
no02f80 g768683 ( .a(n_12108), .b(n_11711), .o(n_12104) );
na02f80 g739316 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_28_), .o(n_40888) );
na02f80 g736746 ( .a(n_43355), .b(n_43339), .o(n_43435) );
na02f80 g760200 ( .a(FE_OCP_RBN3615_n_20249), .b(n_20369), .o(n_20399) );
no02f80 g738298 ( .a(n_41865), .b(n_41578), .o(n_41823) );
na02f80 g746380 ( .a(n_33536), .b(n_33535), .o(n_33537) );
na02f80 FE_RC_2571_0 ( .a(n_43303), .b(n_43350), .o(FE_RN_1056_0) );
in01f80 g736817 ( .a(n_43263), .o(n_43264) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_14_ ( .ck(newNet_1133), .d(n_10652), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_14_) );
no02f80 g776501 ( .a(n_4479), .b(FE_OCP_RBN2490_n_3338), .o(n_4544) );
no02f80 g750852 ( .a(n_29136), .b(n_29053), .o(n_29159) );
in01f80 g754860 ( .a(n_25427), .o(n_25428) );
in01f80 newInst_252 ( .a(newNet_251), .o(newNet_252) );
no02f80 g777122 ( .a(n_3828), .b(n_47023), .o(n_3983) );
na02f80 g769217 ( .a(n_11439), .b(FE_OCP_RBN2916_n_10644), .o(n_11451) );
ao12f80 FE_RC_2764_0 ( .a(FE_RN_1175_0), .b(n_8998), .c(FE_RN_1176_0), .o(FE_RN_1177_0) );
oa12f80 g748610 ( .a(n_31109), .b(n_31273), .c(n_31136), .o(n_31336) );
no02f80 g771532 ( .a(n_9102), .b(FE_OCP_RBN3549_n_44575), .o(n_9317) );
na02f80 g736685 ( .a(n_43436), .b(n_43523), .o(n_43524) );
in01f80 g754292 ( .a(n_46962), .o(n_25957) );
na03f80 g747322 ( .a(n_32578), .b(n_32582), .c(n_32577), .o(n_32625) );
in01f80 FE_RC_1867_0 ( .a(FE_RN_575_0), .o(n_22769) );
in01f80 g770449 ( .a(n_10598), .o(n_10604) );
na02f80 g769677 ( .a(n_11271), .b(n_11263), .o(n_11281) );
no02f80 g743587 ( .a(n_36482), .b(n_36147), .o(n_36504) );
no02f80 g767304 ( .a(n_13678), .b(n_13671), .o(n_13672) );
in01f80 FE_OCP_RBC2202_n_12808 ( .a(n_12808), .o(FE_OCP_RBN2202_n_12808) );
na02f80 g770175 ( .a(n_10796), .b(n_10772), .o(n_10847) );
oa12f80 g773453 ( .a(n_7524), .b(n_7534), .c(n_7523), .o(n_7925) );
oa22f80 g740026 ( .a(n_39784), .b(n_39782), .c(n_39824), .d(n_39783), .o(n_39848) );
in01f80 newInst_3035 ( .a(newNet_3034), .o(newNet_3035) );
in01f80 g768229 ( .a(FE_OCP_RBN3415_n_12739), .o(n_12790) );
in01f80 g739563 ( .a(n_40651), .o(n_40652) );
oa12f80 g771158 ( .a(n_9882), .b(n_9881), .c(n_9880), .o(n_9957) );
in01f80 g739873 ( .a(n_40414), .o(n_40415) );
in01f80 FE_OCP_RBC3059_n_36515 ( .a(n_36515), .o(FE_OCP_RBN3059_n_36515) );
in01f80 g758442 ( .a(n_23317), .o(n_23339) );
na02f80 g772683 ( .a(n_8235), .b(n_7728), .o(n_8346) );
na02f80 g743506 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_0_), .b(delay_add_ln22_unr23_stage9_stallmux_q_24_), .o(n_36624) );
no02f80 g780686 ( .a(n_906), .b(n_905), .o(n_658) );
na02f80 g762389 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18416), .o(n_18658) );
no02f80 g746793 ( .a(n_33075), .b(n_33158), .o(n_33184) );
in01f80 FE_OCP_RBC3672_n_30820 ( .a(n_30820), .o(FE_OCP_RBN3672_n_30820) );
in01f80 newInst_1089 ( .a(newNet_1088), .o(newNet_1089) );
no02f80 g770731 ( .a(n_10141), .b(n_9966), .o(n_10152) );
no02f80 g750177 ( .a(n_29861), .b(FE_OCP_DRV_N1572_n_29860), .o(n_29888) );
in01f80 FE_OCP_RBC3098_n_17315 ( .a(n_17315), .o(FE_OCP_RBN3098_n_17315) );
no02f80 g763277 ( .a(n_17194), .b(n_17193), .o(n_17335) );
in01f80 g780280 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_7_), .o(n_1033) );
in01f80 g739766 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_15_), .o(n_40761) );
in01f80 FE_RC_4209_0 ( .a(FE_OCP_RBN3535_n_13765), .o(FE_RN_1843_0) );
no02f80 g742488 ( .a(n_37596), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37643) );
na02f80 g753417 ( .a(n_27006), .b(n_26456), .o(n_27023) );
na02f80 g771298 ( .a(n_9266), .b(n_9108), .o(n_9297) );
in01f80 newInst_527 ( .a(newNet_35), .o(newNet_527) );
no02f80 g774374 ( .a(n_6816), .b(n_6828), .o(n_7550) );
no02f80 g742209 ( .a(n_44920), .b(n_37852), .o(n_37892) );
no02f80 g775827 ( .a(n_5050), .b(n_5030), .o(n_5136) );
in01f80 g749185 ( .a(n_30750), .o(n_30776) );
no02f80 g759285 ( .a(n_20919), .b(n_20856), .o(n_20942) );
in01f80 newInst_1747 ( .a(newNet_1746), .o(newNet_1747) );
na02f80 g775776 ( .a(n_5584), .b(n_5583), .o(n_5606) );
no02f80 g751483 ( .a(n_28428), .b(n_28406), .o(n_28407) );
na02f80 g746905 ( .a(n_33035), .b(delay_add_ln22_unr20_stage8_stallmux_q_11_), .o(n_33055) );
in01f80 g746276 ( .a(n_33568), .o(n_33569) );
ao12f80 g749719 ( .a(n_31414), .b(n_31311), .c(n_31410), .o(n_31576) );
in01f80 g766392 ( .a(n_14286), .o(n_14186) );
oa22f80 FE_RC_3448_0 ( .a(n_18032), .b(FE_OCP_RBN2390_n_19434), .c(FE_OCPN1800_FE_OFN780_n_17093), .d(n_19434), .o(n_19561) );
no02f80 FE_RC_3202_0 ( .a(FE_RN_1421_0), .b(FE_RN_1422_0), .o(FE_RN_1423_0) );
in01f80 g760976 ( .a(n_19416), .o(n_19417) );
ao12f80 g747142 ( .a(n_33934), .b(n_33952), .c(n_33933), .o(n_34643) );
na02f80 g780892 ( .a(n_521), .b(n_549), .o(n_570) );
in01f80 newInst_3514 ( .a(newNet_3513), .o(newNet_3514) );
oa12f80 g746635 ( .a(n_34473), .b(n_34643), .c(n_33992), .o(n_34634) );
in01f80 g763028 ( .a(n_17678), .o(n_17621) );
in01f80 newInst_1992 ( .a(newNet_1991), .o(newNet_1992) );
in01f80 g744647 ( .a(n_36577), .o(n_36601) );
in01f80 FE_RC_1044_0 ( .a(FE_OCP_RBN3369_n_32436), .o(FE_RN_304_0) );
na02f80 g760227 ( .a(n_20285), .b(n_20262), .o(n_20286) );
no02f80 g764444 ( .a(n_16146), .b(n_14524), .o(n_16195) );
in01f80 newInst_1571 ( .a(newNet_1570), .o(newNet_1571) );
ao12f80 g757315 ( .a(n_22967), .b(n_23071), .c(n_23019), .o(n_23191) );
na02f80 g780486 ( .a(n_664), .b(n_670), .o(n_671) );
in01f80 newInst_134 ( .a(newNet_133), .o(newNet_134) );
na02f80 g754947 ( .a(n_25867), .b(n_26507), .o(n_25882) );
in01f80 g738905 ( .a(n_41316), .o(n_41317) );
na02f80 g766374 ( .a(FE_OCPN3765_FE_OCP_RBN2222_n_13010), .b(n_14278), .o(n_14400) );
na02f80 g756745 ( .a(n_23422), .b(delay_add_ln22_unr14_stage6_stallmux_q_13_), .o(n_23480) );
in01f80 FE_OCP_RBC1686_n_18986 ( .a(FE_OCP_RBN1685_n_18986), .o(FE_OCP_RBN1686_n_18986) );
in01f80 g740518 ( .a(n_39778), .o(n_39755) );
na02f80 g772856 ( .a(n_7968), .b(FE_OCPN915_n_7832), .o(n_8033) );
no02f80 g743026 ( .a(n_37097), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_21_), .o(n_37053) );
ao22s80 FE_RC_49_0 ( .a(n_5378), .b(n_5612), .c(n_5377), .d(n_5611), .o(n_5759) );
no02f80 g765549 ( .a(n_15105), .b(n_13992), .o(n_15144) );
no02f80 g744247 ( .a(n_35487), .b(n_35521), .o(n_35531) );
in01f80 FE_OCP_RBC2209_n_18280 ( .a(n_18280), .o(FE_OCP_RBN2209_n_18280) );
in01f80 g757925 ( .a(n_23055), .o(n_23117) );
oa12f80 g761249 ( .a(n_19682), .b(n_19681), .c(n_19680), .o(n_19912) );
in01f80 g778730 ( .a(n_2838), .o(n_2825) );
ms00f80 cos_out_reg_24_ ( .ck(newNet_3713), .d(n_43884), .o(cos_out_24) );
in01f80 g740098 ( .a(n_40287), .o(n_40288) );
no02f80 g778397 ( .a(n_2488), .b(n_2487), .o(n_2489) );
no02f80 g740900 ( .a(n_44312), .b(n_39134), .o(n_39377) );
no02f80 g755393 ( .a(n_24857), .b(n_22207), .o(n_24858) );
no02f80 g772665 ( .a(n_8272), .b(n_7725), .o(n_8392) );
no02f80 g744503 ( .a(n_35422), .b(n_35412), .o(n_35483) );
na02f80 g738396 ( .a(n_41677), .b(n_41676), .o(n_41678) );
na02f80 g753279 ( .a(FE_OCPN964_n_27287), .b(n_26323), .o(n_27413) );
ao12f80 g740728 ( .a(n_39358), .b(n_39448), .c(n_39425), .o(n_39473) );
na02f80 g769253 ( .a(n_11556), .b(n_11031), .o(n_11673) );
in01f80 newInst_2503 ( .a(newNet_2502), .o(newNet_2503) );
na02f80 g773555 ( .a(n_7439), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_21_), .o(n_7492) );
in01f80 g740011 ( .a(n_39874), .o(n_39875) );
in01f80 fopt782980 ( .a(n_44451), .o(n_44450) );
in01f80 g749152 ( .a(n_30888), .o(n_30943) );
in01f80 FE_OCP_RBC3722_n_39913 ( .a(FE_OCP_RBN3720_n_39913), .o(FE_OCP_RBN3722_n_39913) );
na02f80 g774013 ( .a(n_6889), .b(n_6876), .o(n_6937) );
in01f80 newInst_2484 ( .a(newNet_1527), .o(newNet_2484) );
in01f80 g745294 ( .a(n_35964), .o(n_35965) );
oa12f80 g776007 ( .a(n_4644), .b(n_4986), .c(n_4765), .o(n_5157) );
no02f80 g772661 ( .a(n_8271), .b(n_7726), .o(n_8293) );
na02f80 g745098 ( .a(n_34714), .b(n_34685), .o(n_34686) );
na02f80 g738952 ( .a(n_41241), .b(n_41240), .o(n_41242) );
in01f80 newInst_343 ( .a(newNet_342), .o(newNet_343) );
na02f80 g747247 ( .a(n_32667), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .o(n_32733) );
ao12f80 g754160 ( .a(n_25540), .b(n_25974), .c(n_25973), .o(n_26000) );
oa12f80 g742303 ( .a(n_37783), .b(FE_OCP_RBN3424_n_37794), .c(n_37838), .o(n_37844) );
na02f80 FE_RC_3100_0 ( .a(FE_RN_1370_0), .b(n_16442), .o(n_16466) );
in01f80 FE_OCPC1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(FE_OCPN1224_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCPN1225_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01f80 FE_OCP_RBC3364_n_44722 ( .a(FE_OCP_RBN3306_n_44722), .o(FE_OCP_RBN3364_n_44722) );
in01f80 FE_OCP_RBC2998_n_11004 ( .a(FE_OCP_RBN2997_n_11004), .o(FE_OCP_RBN2998_n_11004) );
oa22f80 g739827 ( .a(n_40381), .b(n_40396), .c(n_40382), .d(n_40397), .o(n_40452) );
ao22s80 FE_RC_1154_0 ( .a(n_10374), .b(n_44575), .c(n_46990), .d(n_44566), .o(n_9034) );
in01f80 newInst_53 ( .a(newNet_52), .o(newNet_53) );
in01f80 FE_OCP_RBC2691_FE_OCPN843_n_3912 ( .a(FE_OCPN843_n_3912), .o(FE_OCP_RBN2691_FE_OCPN843_n_3912) );
no02f80 FE_RC_2106_0 ( .a(FE_RN_727_0), .b(n_20441), .o(FE_RN_728_0) );
no02f80 g766692 ( .a(n_13854), .b(n_13853), .o(n_13855) );
in01f80 newInst_680 ( .a(newNet_679), .o(newNet_680) );
na02f80 g776634 ( .a(n_4300), .b(n_3951), .o(n_4387) );
oa22f80 FE_RC_3355_0 ( .a(n_35307), .b(n_35532), .c(n_35499), .d(n_35323), .o(n_35595) );
na02f80 g748570 ( .a(n_32746), .b(n_32558), .o(n_32776) );
in01f80 g760237 ( .a(n_20459), .o(n_20488) );
in01f80 g777925 ( .a(n_3214), .o(n_3215) );
no02f80 g779605 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .o(n_1685) );
in01f80 g764885 ( .a(n_16177), .o(n_16178) );
no02f80 g777119 ( .a(n_3784), .b(FE_OCPN966_n_47020), .o(n_3841) );
no02f80 g740889 ( .a(n_39368), .b(n_39298), .o(n_39397) );
na02f80 g740615 ( .a(n_39578), .b(n_39560), .o(n_39614) );
in01f80 FE_OCP_RBC2641_n_34921 ( .a(FE_OCP_RBN2640_n_34921), .o(FE_OCP_RBN2641_n_34921) );
in01f80 g765229 ( .a(n_15971), .o(n_16210) );
oa22f80 g768767 ( .a(n_45747), .b(n_11638), .c(n_45748), .d(n_11639), .o(n_12117) );
in01f80 newInst_2366 ( .a(newNet_2365), .o(newNet_2366) );
no02f80 g753905 ( .a(n_26354), .b(n_26353), .o(n_26456) );
in01f80 g746303 ( .a(n_33529), .o(n_33530) );
na02f80 g775742 ( .a(n_5089), .b(n_5045), .o(n_5215) );
na02f80 g773778 ( .a(n_7181), .b(n_6743), .o(n_7270) );
in01f80 g768164 ( .a(FE_OCP_RBN2250_n_13017), .o(n_13437) );
in01f80 newInst_1308 ( .a(newNet_1307), .o(newNet_1308) );
in01f80 g754880 ( .a(n_25775), .o(n_25776) );
no02f80 g773857 ( .a(n_7088), .b(n_7079), .o(n_7080) );
no02f80 g776305 ( .a(n_4568), .b(n_4475), .o(n_4609) );
in01f80 FE_OCPC1386_n_470 ( .a(FE_OCPN1385_n_470), .o(FE_OCPN1386_n_470) );
na02f80 g738055 ( .a(n_42099), .b(n_42196), .o(n_42135) );
in01f80 FE_OFC27_n_1142 ( .a(FE_OFN826_n_1142), .o(FE_OFN27_n_1142) );
na02f80 g763590 ( .a(FE_OCP_RBN3286_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_2_), .o(n_16835) );
na02f80 g772047 ( .a(n_8770), .b(n_8858), .o(n_8898) );
in01f80 g748965 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .o(n_32393) );
in01f80 FE_OCP_RBC1980_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(FE_OCP_RBN1981_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1980_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
no02f80 FE_RC_1601_0 ( .a(FE_RN_447_0), .b(FE_RN_448_0), .o(FE_RN_449_0) );
in01f80 g763889 ( .a(delay_sub_ln23_0_unr12_stage5_stallmux_q_19_), .o(n_17057) );
in01f80 g777972 ( .a(n_3190), .o(n_3191) );
in01f80 FE_RC_710_0 ( .a(n_23138), .o(FE_RN_226_0) );
no02f80 g750594 ( .a(n_29345), .b(n_28847), .o(n_29387) );
no02f80 g762406 ( .a(n_45002), .b(n_18531), .o(n_18655) );
in01f80 g756495 ( .a(n_23846), .o(n_23847) );
na02f80 g781248 ( .a(n_55), .b(n_116), .o(n_133) );
in01f80 g768051 ( .a(n_13111), .o(n_13112) );
na02f80 g770684 ( .a(n_9897), .b(n_9974), .o(n_9982) );
in01f80 FE_OCPC1439_n_23339 ( .a(n_23339), .o(FE_OCPN1439_n_23339) );
ao12f80 g757406 ( .a(n_23461), .b(n_44068), .c(delay_xor_ln21_unr15_stage6_stallmux_q_13_), .o(n_23097) );
na02f80 g765311 ( .a(n_15922), .b(n_15822), .o(n_15959) );
no02f80 g741474 ( .a(n_38759), .b(n_38778), .o(n_38779) );
no02f80 g758039 ( .a(n_22839), .b(n_22842), .o(n_22924) );
na02f80 g766998 ( .a(n_13497), .b(FE_OCPN860_n_12880), .o(n_13573) );
in01f80 newInst_929 ( .a(newNet_529), .o(newNet_929) );
na02f80 g738720 ( .a(n_41386), .b(n_41385), .o(n_41449) );
in01f80 FE_OCP_RBC3046_n_40231 ( .a(n_40231), .o(FE_OCP_RBN3046_n_40231) );
in01f80 FE_OCP_RBC3025_n_39942 ( .a(FE_OCP_RBN3022_n_39942), .o(FE_OCP_RBN3025_n_39942) );
ao12f80 g755910 ( .a(n_25053), .b(n_25188), .c(n_25028), .o(n_25606) );
no02f80 g759361 ( .a(n_21673), .b(n_21295), .o(n_21754) );
oa22f80 FE_RC_3780_0 ( .a(n_24684), .b(n_24870), .c(n_24850), .d(n_24717), .o(n_24934) );
no02f80 g748288 ( .a(n_31612), .b(n_31559), .o(n_31613) );
na02f80 g766383 ( .a(n_14126), .b(n_14063), .o(n_14189) );
in01f80 FE_OCPC1415_FE_OCP_RBN1362_n_20504 ( .a(FE_OCP_RBN1362_n_20504), .o(FE_OCPN1415_FE_OCP_RBN1362_n_20504) );
in01f80 FE_OCPC912_n_43022 ( .a(FE_OCPN911_n_43022), .o(FE_OCPN912_n_43022) );
in01f80 g762635 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_30_), .o(n_17856) );
in01f80 g780722 ( .a(n_809), .o(n_620) );
oa12f80 g743822 ( .a(n_35921), .b(n_35920), .c(n_35919), .o(n_35990) );
in01f80 FE_RC_3587_0 ( .a(n_34765), .o(FE_RN_1565_0) );
no02f80 g746434 ( .a(n_34892), .b(n_34913), .o(n_34943) );
no02f80 FE_RC_2038_0 ( .a(n_26785), .b(FE_RN_681_0), .o(n_26920) );
na02f80 g756027 ( .a(n_24953), .b(n_25000), .o(n_25031) );
na02f80 g763300 ( .a(n_17323), .b(n_17035), .o(n_17324) );
no02f80 g764484 ( .a(n_16010), .b(n_15954), .o(n_16123) );
na02f80 g770457 ( .a(n_10513), .b(n_44463), .o(n_10514) );
na02f80 g776940 ( .a(n_4118), .b(FE_OFN78_n_4117), .o(n_4119) );
no04s80 g768787 ( .a(n_11718), .b(n_11918), .c(n_11927), .d(n_11919), .o(n_11998) );
ao12f80 g751296 ( .a(n_29652), .b(n_29651), .c(n_29650), .o(n_29709) );
no02f80 g765054 ( .a(n_15490), .b(n_15530), .o(n_15640) );
na02f80 g771544 ( .a(n_9086), .b(FE_OCPN1251_n_8210), .o(n_9212) );
no02f80 g770962 ( .a(n_9507), .b(n_9582), .o(n_9630) );
in01f80 newInst_3211 ( .a(newNet_3210), .o(newNet_3211) );
no02f80 g760295 ( .a(FE_OCPN1261_n_20242), .b(n_19455), .o(n_20518) );
ao12f80 g741555 ( .a(n_38778), .b(n_38654), .c(n_38624), .o(n_38667) );
in01f80 newInst_1333 ( .a(newNet_1332), .o(newNet_1333) );
no02f80 FE_RC_3481_0 ( .a(FE_RN_1496_0), .b(n_40466), .o(n_40472) );
no02f80 g753629 ( .a(n_26630), .b(n_26277), .o(n_26697) );
in01f80 newInst_720 ( .a(newNet_719), .o(newNet_720) );
in01f80 g773143 ( .a(n_7768), .o(n_7740) );
na02f80 g756605 ( .a(FE_OFN745_n_23604), .b(n_23603), .o(n_23684) );
no02f80 g743729 ( .a(n_36309), .b(n_35752), .o(n_36343) );
no02f80 g756917 ( .a(n_23617), .b(n_22788), .o(n_23750) );
ao12f80 g737328 ( .a(n_42648), .b(n_42834), .c(n_42503), .o(n_42857) );
no02f80 g747393 ( .a(n_33574), .b(n_33416), .o(n_33575) );
in01f80 g759090 ( .a(n_21194), .o(n_21226) );
in01f80 newInst_2730 ( .a(newNet_2729), .o(newNet_2730) );
ao12f80 g746860 ( .a(n_33149), .b(FE_OCP_RBN3385_n_33108), .c(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n_33637) );
in01f80 g745819 ( .a(n_34184), .o(n_34161) );
oa22f80 FE_RC_3382_0 ( .a(n_37060), .b(n_37509), .c(n_37059), .d(n_37510), .o(n_37606) );
na02f80 g753940 ( .a(n_26167), .b(n_26120), .o(n_26224) );
in01f80 g737263 ( .a(n_42954), .o(n_42955) );
in01f80 g770083 ( .a(n_10827), .o(n_10855) );
na02f80 g752951 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_10_), .o(n_27848) );
in01f80 g751993 ( .a(n_28955), .o(n_28956) );
in01f80 newInst_1237 ( .a(newNet_1236), .o(newNet_1237) );
na02f80 g771063 ( .a(n_9621), .b(FE_OCP_RBN2619_n_44561), .o(n_9804) );
in01f80 g741790 ( .a(n_38448), .o(n_38449) );
no02f80 g751903 ( .a(n_28864), .b(n_28984), .o(n_28883) );
na02f80 g781027 ( .a(sin_out_2), .b(FE_OFN5_n_43918), .o(n_306) );
na02f80 g774928 ( .a(n_6197), .b(n_6148), .o(n_6191) );
in01f80 newInst_1924 ( .a(newNet_1923), .o(newNet_1924) );
ao12f80 g760628 ( .a(n_19438), .b(n_19707), .c(n_19505), .o(n_19781) );
oa22f80 FE_RC_726_0 ( .a(n_7430), .b(n_8211), .c(n_7431), .d(n_8212), .o(n_8321) );
in01f80 g777886 ( .a(n_3204), .o(n_3198) );
na02f80 g742223 ( .a(n_37598), .b(FE_OCP_RBN3425_n_44881), .o(n_37996) );
no02f80 g768917 ( .a(n_12053), .b(n_11895), .o(n_12054) );
oa12f80 g754600 ( .a(n_25203), .b(n_25403), .c(n_25268), .o(n_25515) );
na02f80 g759317 ( .a(n_21263), .b(n_21257), .o(n_21258) );
in01f80 newInst_1773 ( .a(newNet_1772), .o(newNet_1773) );
in01f80 g757492 ( .a(n_22933), .o(n_22934) );
no02f80 g772430 ( .a(n_8503), .b(n_8494), .o(n_8495) );
in01f80 FE_RC_2646_0 ( .a(FE_RN_1104_0), .o(n_32905) );
in01f80 g777313 ( .a(n_4215), .o(n_4292) );
in01f80 g754181 ( .a(n_25999), .o(n_27117) );
in01f80 g778357 ( .a(n_2531), .o(n_2532) );
no02f80 g777764 ( .a(n_3410), .b(n_3409), .o(n_3411) );
in01f80 g746158 ( .a(n_33717), .o(n_33733) );
no02f80 g774035 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_28_), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n_6784) );
oa22f80 g742425 ( .a(n_37689), .b(n_37574), .c(n_37755), .d(n_37556), .o(n_37771) );
na02f80 g747809 ( .a(n_33571), .b(n_33438), .o(n_33624) );
in01f80 FE_OCP_DRV_C1586_n_35594 ( .a(FE_OCP_DRV_N1585_n_35594), .o(FE_OCP_DRV_N1586_n_35594) );
oa12f80 g778077 ( .a(n_2724), .b(n_2891), .c(n_2669), .o(n_3013) );
na02f80 g756706 ( .a(n_23504), .b(n_23161), .o(n_23505) );
no02f80 g765347 ( .a(n_15180), .b(n_14169), .o(n_15228) );
na02f80 g766960 ( .a(n_13825), .b(n_13824), .o(n_13826) );
na02f80 g771408 ( .a(n_9523), .b(n_9440), .o(n_9549) );
no02f80 g742640 ( .a(n_37417), .b(n_37151), .o(n_37463) );
no02f80 g736411 ( .a(n_43800), .b(n_43657), .o(n_43820) );
no02f80 g765097 ( .a(n_15459), .b(n_15458), .o(n_15530) );
in01f80 g771648 ( .a(n_9010), .o(n_9011) );
ao12f80 g784619 ( .a(n_39533), .b(n_39532), .c(n_39072), .o(n_46948) );
in01f80 g773335 ( .a(n_8309), .o(n_8232) );
no02f80 g749621 ( .a(n_30458), .b(n_30457), .o(n_30459) );
in01f80 g760938 ( .a(n_19358), .o(n_19386) );
no03m80 FE_RC_1666_0 ( .a(FE_OCP_RBN2185_FE_RN_464_0), .b(n_37659), .c(n_37602), .o(n_37755) );
oa12f80 g752649 ( .a(n_27527), .b(n_27442), .c(n_27454), .o(n_27555) );
no02f80 g757297 ( .a(n_23064), .b(FE_OCPN3170_n_23227), .o(n_23173) );
no02f80 g746394 ( .a(n_33458), .b(n_32999), .o(n_33486) );
no02f80 g771962 ( .a(n_44463), .b(n_9631), .o(n_9651) );
in01f80 g763314 ( .a(n_46974), .o(n_17003) );
no02f80 g772835 ( .a(n_7903), .b(n_7869), .o(n_8269) );
in01f80 g765776 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_1_), .o(n_17193) );
in01f80 g758595 ( .a(n_22549), .o(n_22550) );
ao12f80 g766516 ( .a(n_14080), .b(n_14457), .c(n_14078), .o(n_14566) );
no02f80 g780572 ( .a(n_745), .b(n_783), .o(n_819) );
no03m80 g772368 ( .a(n_8550), .b(n_8656), .c(n_7965), .o(n_8707) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_27_ ( .ck(newNet_2267), .d(n_40552), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_) );
no02f80 g742705 ( .a(n_37397), .b(n_37098), .o(n_37410) );
na02f80 g736960 ( .a(n_43038), .b(n_42923), .o(n_43306) );
in01f80 newInst_911 ( .a(newNet_910), .o(newNet_911) );
in01f80 g760375 ( .a(n_20207), .o(n_20208) );
na02f80 g776497 ( .a(n_4356), .b(n_4063), .o(n_4538) );
no02f80 g744491 ( .a(n_35428), .b(FE_OCP_DRV_N1540_n_35427), .o(n_35535) );
in01f80 g751558 ( .a(n_28520), .o(n_28521) );
in01f80 newInst_2133 ( .a(newNet_1104), .o(newNet_2133) );
na02f80 g778391 ( .a(FE_OCP_RBN2273_n_2457), .b(n_2492), .o(n_2493) );
in01f80 FE_OCP_RBC2778_n_15595 ( .a(FE_OCP_RBN2777_n_15595), .o(FE_OCP_RBN2778_n_15595) );
no02f80 g752913 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_12_), .o(n_28297) );
na02f80 g773940 ( .a(n_7217), .b(delay_xor_ln22_unr6_stage3_stallmux_q_25_), .o(n_7278) );
in01f80 g756150 ( .a(n_24204), .o(n_25318) );
na02f80 g746028 ( .a(n_33941), .b(FE_OCP_RBN3456_n_33872), .o(n_33980) );
oa22f80 g747968 ( .a(n_31937), .b(n_31914), .c(n_31936), .d(n_31915), .o(n_31998) );
in01f80 FE_OCP_DRV_C3161_n_21419 ( .a(n_21419), .o(FE_OCP_DRV_N3161_n_21419) );
no02f80 g737077 ( .a(n_43120), .b(n_42942), .o(n_43325) );
na03f80 g740842 ( .a(n_39163), .b(n_39436), .c(n_39319), .o(n_39510) );
no02f80 g778599 ( .a(n_2705), .b(n_2803), .o(n_3351) );
in01f80 FE_OCP_RBC3823_n_44061 ( .a(n_44061), .o(FE_OCP_RBN3823_n_44061) );
oa22f80 g758200 ( .a(n_21453), .b(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .c(FE_OCP_RBN2049_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .d(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_22737) );
na02f80 g771255 ( .a(n_9371), .b(n_9302), .o(n_9546) );
no02f80 g752968 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_16_), .o(n_28259) );
no02f80 g763038 ( .a(n_17450), .b(n_17225), .o(n_17512) );
na02f80 g765008 ( .a(n_15497), .b(n_15608), .o(n_15673) );
na02f80 g771392 ( .a(n_9087), .b(FE_OCP_RBN3523_n_8242), .o(n_9142) );
no02f80 g749137 ( .a(n_30860), .b(n_30859), .o(n_30942) );
na02f80 g762901 ( .a(n_17595), .b(n_17190), .o(n_17596) );
na02f80 g776032 ( .a(n_4915), .b(FE_OCPN846_n_4046), .o(n_4957) );
in01f80 g740371 ( .a(n_39807), .o(n_39833) );
na02f80 g778977 ( .a(n_2202), .b(n_2182), .o(n_2216) );
no02f80 g747800 ( .a(n_33372), .b(n_32802), .o(n_33840) );
ao12f80 g750721 ( .a(n_29268), .b(n_29299), .c(n_29267), .o(n_29373) );
in01f80 g756314 ( .a(n_24605), .o(n_25122) );
na02f80 g777662 ( .a(n_3495), .b(n_3494), .o(n_3586) );
in01f80 g754582 ( .a(n_26926), .o(n_26927) );
in01f80 g751954 ( .a(n_28902), .o(n_28881) );
no02f80 FE_RC_2049_0 ( .a(FE_RN_689_0), .b(FE_RN_690_0), .o(FE_RN_691_0) );
in01f80 g756509 ( .a(n_23917), .o(n_23918) );
in01f80 g758238 ( .a(n_22840), .o(n_22807) );
na02f80 g762291 ( .a(n_18532), .b(n_18657), .o(n_19070) );
na02f80 g753598 ( .a(n_26723), .b(n_26655), .o(n_26750) );
in01f80 g775037 ( .a(n_5923), .o(n_5924) );
in01f80 newInst_2735 ( .a(newNet_2293), .o(newNet_2735) );
in01f80 g777304 ( .a(n_4200), .o(n_4201) );
in01f80 g778164 ( .a(n_2888), .o(n_2889) );
in01f80 FE_OCP_RBC3357_delay_xor_ln22_unr28_stage10_stallmux_q_0_ ( .a(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(FE_OCP_RBN3357_delay_xor_ln22_unr28_stage10_stallmux_q_0_) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_28_ ( .ck(newNet_1713), .d(n_22606), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_28_) );
in01f80 newInst_1709 ( .a(newNet_1708), .o(newNet_1709) );
in01f80 g748501 ( .a(n_31548), .o(n_31591) );
na02f80 FE_RC_2428_0 ( .a(FE_RN_964_0), .b(n_7270), .o(FE_RN_965_0) );
in01f80 g758624 ( .a(n_21987), .o(n_21988) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_29_ ( .ck(newNet_2630), .d(n_22875), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_29_) );
in01f80 g744237 ( .a(n_36870), .o(n_36871) );
no02f80 g752789 ( .a(n_28051), .b(n_27992), .o(n_28079) );
na02f80 FE_RC_3852_0 ( .a(FE_RN_1680_0), .b(n_19633), .o(FE_RN_1681_0) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_20_ ( .ck(newNet_2856), .d(n_11605), .o(delay_add_ln22_unr8_stage4_stallmux_q_20_) );
ao12f80 g748358 ( .a(n_32727), .b(n_32726), .c(n_32725), .o(n_33279) );
no02f80 g768965 ( .a(FE_OCP_RBN2119_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .o(n_12311) );
in01f80 newInst_873 ( .a(newNet_872), .o(newNet_873) );
na02f80 g779736 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_), .o(n_1792) );
in01f80 newInst_767 ( .a(newNet_766), .o(newNet_767) );
na02f80 g737721 ( .a(n_42195), .b(n_41505), .o(n_42239) );
na02f80 g765299 ( .a(n_15716), .b(n_15783), .o(n_16479) );
no02f80 g748318 ( .a(n_31704), .b(FE_OCPN977_n_31594), .o(n_31800) );
na02f80 g753393 ( .a(n_26882), .b(n_26754), .o(n_26970) );
ao12f80 g756829 ( .a(n_23291), .b(n_23365), .c(n_23281), .o(n_23405) );
in01f80 g767955 ( .a(n_12857), .o(n_12923) );
na02f80 g752558 ( .a(n_27598), .b(n_27297), .o(n_27600) );
na02f80 g747007 ( .a(n_32988), .b(n_32955), .o(n_33010) );
ao12f80 g768375 ( .a(n_12192), .b(n_12467), .c(n_12270), .o(n_12519) );
na02f80 g769387 ( .a(n_10388), .b(n_11507), .o(n_11571) );
na02f80 g753288 ( .a(n_27110), .b(n_26652), .o(n_27375) );
na02f80 g762696 ( .a(n_17922), .b(n_17921), .o(n_17947) );
oa22f80 FE_RC_1374_0 ( .a(n_25720), .b(n_26040), .c(n_25719), .d(n_26041), .o(n_26169) );
no02f80 g751601 ( .a(FE_OCP_RBN3404_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_27_), .o(n_28723) );
na02f80 g760450 ( .a(n_20049), .b(n_19867), .o(n_20079) );
na02f80 g741149 ( .a(n_39126), .b(n_39121), .o(n_39185) );
na02f80 g754845 ( .a(n_25389), .b(n_25388), .o(n_25487) );
in01f80 newInst_1138 ( .a(newNet_1137), .o(newNet_1138) );
in01f80 g756642 ( .a(n_23577), .o(n_23578) );
no02f80 g743042 ( .a(n_37109), .b(n_37110), .o(n_37485) );
in01f80 newInst_337 ( .a(newNet_336), .o(newNet_337) );
in01f80 g737005 ( .a(n_43387), .o(n_43420) );
no02f80 g742900 ( .a(n_37000), .b(n_37012), .o(n_37375) );
ms00f80 sin_out_reg_21_ ( .ck(newNet_55), .d(n_43899), .o(sin_out_21) );
in01f80 g762251 ( .a(n_18661), .o(n_18735) );
in01f80 newInst_2662 ( .a(newNet_2661), .o(newNet_2662) );
no02f80 g747636 ( .a(n_32328), .b(n_32020), .o(n_32359) );
no02f80 g750547 ( .a(n_30441), .b(n_29937), .o(n_30442) );
ao12f80 g742729 ( .a(n_37443), .b(n_37442), .c(n_37441), .o(n_37518) );
in01f80 newInst_474 ( .a(newNet_473), .o(newNet_474) );
na02f80 g780743 ( .a(n_591), .b(n_438), .o(n_596) );
na02f80 g761065 ( .a(n_19174), .b(n_18784), .o(n_19248) );
na02f80 g741141 ( .a(n_38988), .b(n_38588), .o(n_38989) );
in01f80 FE_RC_1567_0 ( .a(n_28334), .o(FE_RN_445_0) );
in01f80 g769847 ( .a(n_11267), .o(n_11233) );
in01f80 newInst_661 ( .a(newNet_660), .o(newNet_661) );
in01f80 g737265 ( .a(n_46938), .o(n_42953) );
no02f80 g777725 ( .a(n_3413), .b(n_3383), .o(n_3437) );
in01f80 g772610 ( .a(n_8206), .o(n_8207) );
na02f80 g750123 ( .a(FE_OCP_RBN3566_n_29857), .b(n_29055), .o(n_30007) );
no02f80 g770997 ( .a(n_9989), .b(n_9988), .o(n_10031) );
no02f80 FE_RC_2572_0 ( .a(FE_RN_1056_0), .b(n_43360), .o(FE_RN_1057_0) );
no02f80 g769208 ( .a(n_11631), .b(n_11630), .o(n_12033) );
in01f80 FE_OCP_RBC3703_n_26231 ( .a(FE_OCP_RBN2957_n_26231), .o(FE_OCP_RBN3703_n_26231) );
oa12f80 g764119 ( .a(n_16017), .b(n_16930), .c(n_16099), .o(n_16962) );
no02f80 g749928 ( .a(n_30470), .b(n_30198), .o(n_30199) );
no02f80 g778640 ( .a(n_2249), .b(n_2211), .o(n_2299) );
na02f80 g774747 ( .a(n_6265), .b(n_5636), .o(n_6292) );
in01f80 FE_OFC77_n_4117 ( .a(n_4117), .o(FE_OFN77_n_4117) );
na02f80 g763291 ( .a(n_17332), .b(n_17331), .o(n_17333) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_1_ ( .ck(newNet_1853), .d(n_16409), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_1_) );
in01f80 FE_OCPC1407_n_672 ( .a(n_672), .o(FE_OCPN1407_n_672) );
in01f80 newInst_1287 ( .a(newNet_1286), .o(newNet_1287) );
in01f80 FE_OCP_RBC3468_n_7886 ( .a(FE_OCP_RBN3462_n_7886), .o(FE_OCP_RBN3468_n_7886) );
in01f80 g778670 ( .a(n_2348), .o(n_2322) );
no02f80 g771216 ( .a(n_9720), .b(n_9407), .o(n_9757) );
na02f80 g765205 ( .a(n_15578), .b(n_15518), .o(n_15579) );
na02f80 g766502 ( .a(FE_OCPN1420_n_14003), .b(n_14004), .o(n_14101) );
no02f80 g771467 ( .a(n_9526), .b(n_9525), .o(n_9656) );
oa12f80 g781269 ( .a(n_7), .b(beta_24), .c(beta_23), .o(n_89) );
in01f80 g737845 ( .a(n_42203), .o(n_42216) );
in01f80 FE_OCP_RBC3608_n_14905 ( .a(n_14905), .o(FE_OCP_RBN3608_n_14905) );
na02f80 g759896 ( .a(n_21051), .b(n_21251), .o(n_21379) );
in01f80 newInst_3343 ( .a(newNet_3342), .o(newNet_3343) );
in01f80 g738032 ( .a(n_42150), .o(n_42197) );
in01f80 g743752 ( .a(n_36275), .o(n_36276) );
in01f80 g742059 ( .a(n_38281), .o(n_38282) );
in01f80 newInst_498 ( .a(newNet_497), .o(newNet_498) );
na02f80 g755794 ( .a(n_25060), .b(n_25059), .o(n_25061) );
na02f80 g773665 ( .a(n_7298), .b(n_7297), .o(n_7299) );
in01f80 newInst_1871 ( .a(newNet_1870), .o(newNet_1871) );
na02f80 g738416 ( .a(n_41674), .b(n_41546), .o(n_41933) );
in01f80 newInst_1577 ( .a(newNet_1191), .o(newNet_1577) );
in01f80 newInst_13 ( .a(newNet_12), .o(newNet_13) );
na02f80 g741030 ( .a(n_39007), .b(n_39006), .o(n_39008) );
na02f80 g751578 ( .a(n_28437), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_18_), .o(n_28548) );
no02f80 g752006 ( .a(n_28919), .b(n_29067), .o(n_29098) );
na02f80 g763015 ( .a(n_17667), .b(delay_add_ln22_unr11_stage5_stallmux_q_6_), .o(n_17739) );
no02f80 g745545 ( .a(n_35509), .b(n_35508), .o(n_35510) );
na02f80 g737000 ( .a(n_43097), .b(n_42955), .o(n_43339) );
no02f80 g764254 ( .a(n_16376), .b(n_16375), .o(n_16463) );
ao12f80 g745234 ( .a(n_34376), .b(n_34465), .c(n_34310), .o(n_34492) );
na02f80 g776997 ( .a(n_4208), .b(n_3941), .o(n_4145) );
no02f80 g740226 ( .a(n_40099), .b(FE_OCP_RBN3022_n_39942), .o(n_40176) );
na02f80 FE_RC_3675_0 ( .a(FE_RN_1614_0), .b(n_46969), .o(n_21044) );
ao12f80 g765588 ( .a(n_15874), .b(n_15085), .c(n_15865), .o(n_16059) );
oa12f80 g766752 ( .a(n_14084), .b(n_14085), .c(n_14083), .o(n_16246) );
no02f80 g770838 ( .a(n_10138), .b(n_10137), .o(n_10257) );
in01f80 g756669 ( .a(n_23581), .o(n_23606) );
no02f80 g773419 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_30_), .o(n_7547) );
in01f80 g758030 ( .a(n_22379), .o(n_22380) );
oa12f80 g775351 ( .a(n_5776), .b(n_5775), .c(n_5774), .o(n_5853) );
no02f80 g741252 ( .a(n_38870), .b(n_38565), .o(n_39026) );
in01f80 g738532 ( .a(n_41450), .o(n_41511) );
in01f80 FE_OCP_RBC3391_n_37557 ( .a(n_37557), .o(FE_OCP_RBN3391_n_37557) );
no02f80 g756671 ( .a(n_23507), .b(n_23506), .o(n_23508) );
in01f80 g777020 ( .a(n_3995), .o(n_3996) );
in01f80 FE_OCP_RBC2182_n_1916 ( .a(n_1916), .o(FE_OCP_RBN2182_n_1916) );
in01f80 g748899 ( .a(n_32508), .o(n_32392) );
oa12f80 g763021 ( .a(n_16986), .b(n_17483), .c(n_17515), .o(n_17516) );
oa12f80 g755283 ( .a(n_25581), .b(n_25580), .c(n_25579), .o(n_25686) );
no02f80 g743247 ( .a(n_38044), .b(n_46242), .o(n_38045) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_15_ ( .ck(newNet_1247), .d(n_5664), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_15_) );
na02f80 g753880 ( .a(n_26363), .b(n_26319), .o(n_26394) );
no02f80 g769349 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_), .o(n_11711) );
in01f80 FE_RC_3517_0 ( .a(n_23017), .o(FE_RN_1519_0) );
no02f80 g769679 ( .a(n_11247), .b(FE_OCP_RBN3038_n_47269), .o(n_11248) );
no02f80 g759104 ( .a(n_21345), .b(n_45073), .o(n_21423) );
no02f80 g739407 ( .a(n_40686), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .o(n_40728) );
no03m80 g742924 ( .a(n_37093), .b(n_37160), .c(n_37100), .o(n_37219) );
na02f80 g753564 ( .a(n_26702), .b(n_26701), .o(n_26703) );
na02f80 g764833 ( .a(n_15726), .b(n_15793), .o(n_15890) );
in01f80 g775561 ( .a(n_5739), .o(n_5740) );
na02f80 g763829 ( .a(n_17097), .b(n_17202), .o(n_17258) );
na02f80 g752345 ( .a(n_27888), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_0_), .o(n_27887) );
in01f80 g775989 ( .a(n_4925), .o(n_6030) );
na02f80 g775098 ( .a(n_6074), .b(n_5049), .o(n_6188) );
in01f80 g758156 ( .a(n_22726), .o(n_22727) );
ao12f80 g760771 ( .a(n_19627), .b(n_19626), .c(n_19625), .o(n_19715) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_19_ ( .ck(newNet_3627), .d(n_17199), .o(delay_add_ln22_unr11_stage5_stallmux_q_19_) );
na02f80 g759553 ( .a(n_20764), .b(n_20463), .o(n_20796) );
na02f80 g758886 ( .a(n_21430), .b(n_21542), .o(n_21543) );
in01f80 g778169 ( .a(n_2907), .o(n_2908) );
in01f80 FE_RC_471_0 ( .a(n_28893), .o(FE_RN_139_0) );
na02f80 g753748 ( .a(n_26448), .b(n_26472), .o(n_26553) );
in01f80 g750385 ( .a(n_29677), .o(n_29678) );
no02f80 g742599 ( .a(n_38315), .b(n_37520), .o(n_37590) );
in01f80 g778898 ( .a(n_2235), .o(n_2256) );
oa12f80 g736264 ( .a(n_322), .b(n_43900), .c(FE_OFN4_n_43918), .o(n_43914) );
no02f80 g754089 ( .a(n_26020), .b(n_23317), .o(n_26067) );
no03m80 g762060 ( .a(n_18932), .b(n_18931), .c(n_18882), .o(n_18933) );
ao12f80 g741510 ( .a(n_38724), .b(n_38742), .c(n_38755), .o(n_38774) );
na02f80 g762781 ( .a(n_17720), .b(n_17894), .o(n_17780) );
oa22f80 FE_RC_799_0 ( .a(FE_OCP_RBN3475_n_7886), .b(n_8828), .c(n_8189), .d(n_8842), .o(n_8974) );
ao12f80 g748370 ( .a(n_32442), .b(n_32674), .c(n_32588), .o(n_32750) );
no02f80 g778331 ( .a(n_2841), .b(n_2834), .o(n_2909) );
ao12f80 g774119 ( .a(n_7123), .b(n_6872), .c(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .o(n_7177) );
in01f80 g736630 ( .a(n_43625), .o(n_43646) );
na02f80 g745532 ( .a(n_34380), .b(n_34374), .o(n_34850) );
in01f80 FE_OCP_RBC3720_n_39913 ( .a(FE_OCP_RBN3719_n_39913), .o(FE_OCP_RBN3720_n_39913) );
na02f80 g775436 ( .a(n_5434), .b(n_5529), .o(n_5530) );
in01f80 newInst_96 ( .a(newNet_95), .o(newNet_96) );
no02f80 g742240 ( .a(n_44881), .b(n_37692), .o(n_38130) );
in01f80 g757505 ( .a(n_22930), .o(n_22931) );
no02f80 g760490 ( .a(n_20513), .b(n_20512), .o(n_20514) );
no02f80 g768265 ( .a(n_12623), .b(n_12610), .o(n_12611) );
in01f80 newInst_1549 ( .a(newNet_973), .o(newNet_1549) );
in01f80 FE_RC_2552_0 ( .a(n_36998), .o(FE_RN_1045_0) );
na02f80 g740237 ( .a(n_39807), .b(n_39808), .o(n_39838) );
no02f80 g760825 ( .a(n_19390), .b(n_18032), .o(n_19440) );
in01f80 g741125 ( .a(n_39299), .o(n_39300) );
in01f80 g767710 ( .a(n_13320), .o(n_13321) );
na02f80 g769090 ( .a(n_11684), .b(n_11532), .o(n_11685) );
na02f80 g738201 ( .a(n_41942), .b(n_41789), .o(n_41995) );
in01f80 FE_OCP_RBC3026_n_39942 ( .a(FE_OCP_RBN3023_n_39942), .o(FE_OCP_RBN3026_n_39942) );
na02f80 g766057 ( .a(n_14645), .b(n_14376), .o(n_14646) );
no02f80 g755381 ( .a(n_24858), .b(n_24873), .o(n_24932) );
in01f80 g781208 ( .a(n_501), .o(n_375) );
na02f80 g760614 ( .a(n_19812), .b(n_19778), .o(n_19813) );
oa12f80 g763773 ( .a(n_17015), .b(n_17263), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_7_), .o(n_17265) );
in01f80 FE_OCP_RBC1366_n_20879 ( .a(n_20879), .o(FE_OCP_RBN1366_n_20879) );
no02f80 g751976 ( .a(n_28836), .b(n_28835), .o(n_28863) );
no02f80 g760418 ( .a(n_20075), .b(n_20266), .o(n_20149) );
in01f80 g762911 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_22_), .o(n_17625) );
in01f80 FE_OCPC958_n_3951 ( .a(n_3951), .o(FE_OCPN958_n_3951) );
na02f80 g759070 ( .a(n_21494), .b(FE_OCP_DRV_N1600_n_21493), .o(n_21603) );
no02f80 g760749 ( .a(n_19603), .b(n_19362), .o(n_19635) );
no02f80 g768499 ( .a(n_45659), .b(delay_xor_ln21_unr9_stage4_stallmux_q_18_), .o(n_12372) );
na02f80 g777813 ( .a(n_3362), .b(n_3361), .o(n_3388) );
in01f80 g756995 ( .a(n_23287), .o(n_23288) );
no02f80 g743315 ( .a(n_36755), .b(n_36735), .o(n_36778) );
oa22f80 FE_RC_4131_0 ( .a(n_17085), .b(n_17247), .c(n_17086), .d(n_17245), .o(n_17348) );
in01f80 FE_RC_2379_0 ( .a(n_12168), .o(FE_RN_927_0) );
in01f80 g780663 ( .a(n_745), .o(n_779) );
no02f80 FE_RC_2401_0 ( .a(FE_RN_943_0), .b(FE_RN_946_0), .o(n_42896) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_2_ ( .ck(newNet_561), .d(n_16747), .o(delay_xor_ln22_unr12_stage5_stallmux_q_2_) );
no02f80 g754348 ( .a(n_25764), .b(n_25416), .o(n_25849) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_23_ ( .ck(newNet_1732), .d(n_22568), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_) );
no02f80 g755734 ( .a(n_25222), .b(n_25771), .o(n_25311) );
in01f80 g767204 ( .a(n_14419), .o(n_14452) );
na02f80 g770556 ( .a(FE_OCP_RBN2843_n_10326), .b(FE_OCP_RBN2621_n_44561), .o(n_10397) );
na02f80 g738197 ( .a(n_41976), .b(n_41859), .o(n_42027) );
in01f80 newInst_2010 ( .a(newNet_2009), .o(newNet_2010) );
in01f80 g768728 ( .a(n_12283), .o(n_12284) );
in01f80 newInst_1135 ( .a(newNet_1134), .o(newNet_1135) );
in01f80 newInst_371 ( .a(newNet_5), .o(newNet_371) );
no02f80 g780900 ( .a(n_374), .b(n_387), .o(n_395) );
in01f80 g752974 ( .a(n_28195), .o(n_28196) );
no02f80 g739607 ( .a(n_40624), .b(n_44610), .o(n_40626) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_22_ ( .ck(newNet_630), .d(n_46340), .o(delay_xor_ln21_unr9_stage4_stallmux_q_22_) );
in01f80 g775058 ( .a(n_6064), .o(n_6065) );
na02f80 g749290 ( .a(n_32063), .b(n_31318), .o(n_32156) );
na02f80 g749632 ( .a(n_31434), .b(n_31536), .o(n_31644) );
in01f80 newInst_1807 ( .a(newNet_98), .o(newNet_1807) );
in01f80 g736697 ( .a(n_43468), .o(n_43469) );
in01f80 g781321 ( .a(n_42), .o(n_43) );
in01f80 g758630 ( .a(n_21900), .o(n_21918) );
na02f80 g764469 ( .a(n_16160), .b(n_16189), .o(n_16423) );
in01f80 newInst_2440 ( .a(newNet_2439), .o(newNet_2440) );
no02f80 g781118 ( .a(n_223), .b(n_122), .o(n_231) );
no02f80 g775288 ( .a(FE_OCP_RBN2976_n_5555), .b(n_4759), .o(n_5600) );
ao12f80 g748769 ( .a(n_32425), .b(n_46107), .c(delay_sub_ln23_0_unr24_stage8_stallmux_q_23_), .o(n_33171) );
ao22s80 g757078 ( .a(n_23521), .b(n_23150), .c(n_23522), .d(n_23151), .o(n_23863) );
in01f80 g750666 ( .a(n_30192), .o(n_29395) );
ao22s80 FE_RC_1024_0 ( .a(n_45024), .b(n_20965), .c(n_45010), .d(n_20935), .o(n_21064) );
in01f80 newInst_193 ( .a(newNet_1), .o(newNet_193) );
oa22f80 FE_RC_1264_0 ( .a(n_6351), .b(n_6418), .c(n_6350), .d(n_6388), .o(n_6529) );
in01f80 g753591 ( .a(n_26724), .o(n_26725) );
no02f80 g750730 ( .a(n_30340), .b(n_30339), .o(n_30341) );
ao12f80 g745169 ( .a(n_34434), .b(n_34656), .c(n_34412), .o(n_34725) );
oa22f80 FE_RC_3372_0 ( .a(n_22801), .b(n_22718), .c(n_22833), .d(n_22679), .o(n_22777) );
oa22f80 g748859 ( .a(n_31778), .b(delay_sub_ln23_unr25_stage8_stallmux_q_1_), .c(n_32393), .d(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_32589) );
na02f80 g741019 ( .a(n_38965), .b(FE_OCP_RBN2638_n_38806), .o(n_39059) );
na02f80 g772844 ( .a(n_8029), .b(n_8072), .o(n_8154) );
in01f80 g744917 ( .a(n_34982), .o(n_34981) );
no02f80 g736776 ( .a(n_43352), .b(n_43351), .o(n_43398) );
in01f80 g771617 ( .a(n_10343), .o(n_10344) );
no02f80 g781299 ( .a(beta_31), .b(beta_15), .o(n_109) );
oa12f80 g752756 ( .a(n_27020), .b(n_27058), .c(n_26980), .o(n_27104) );
no02f80 g758021 ( .a(FE_OCPN991_n_22249), .b(n_22376), .o(n_22441) );
no02f80 g767776 ( .a(n_13043), .b(n_12928), .o(n_13044) );
in01f80 g767683 ( .a(n_13022), .o(n_13023) );
in01f80 newInst_2396 ( .a(newNet_2395), .o(newNet_2396) );
in01f80 g754277 ( .a(n_25934), .o(n_27217) );
in01f80 newInst_1319 ( .a(newNet_1318), .o(newNet_1319) );
ao22s80 g762066 ( .a(n_18247), .b(n_18125), .c(n_18201), .d(n_18124), .o(n_19885) );
in01f80 newInst_2880 ( .a(newNet_1963), .o(newNet_2880) );
no02f80 g767610 ( .a(n_13700), .b(n_13286), .o(n_13287) );
na02f80 g763703 ( .a(n_16719), .b(FE_OCP_RBN2741_n_15206), .o(n_16758) );
in01f80 g776231 ( .a(n_4657), .o(n_4658) );
na02f80 g780889 ( .a(n_403), .b(n_399), .o(n_438) );
in01f80 g743890 ( .a(n_35712), .o(n_35793) );
na02f80 g771874 ( .a(n_9004), .b(n_9003), .o(n_9036) );
no02f80 g759616 ( .a(n_20643), .b(n_20617), .o(n_20763) );
no02f80 g777845 ( .a(n_3259), .b(n_2913), .o(n_3269) );
no02f80 g742438 ( .a(n_37649), .b(n_37709), .o(n_37670) );
no02f80 FE_RC_3052_0 ( .a(n_35312), .b(n_35379), .o(FE_RN_1338_0) );
na02f80 g748639 ( .a(n_31488), .b(n_31490), .o(n_31489) );
no02f80 g784604 ( .a(n_5952), .b(n_5940), .o(n_46427) );
in01f80 FE_OCP_RBC2590_n_14460 ( .a(n_14460), .o(FE_OCP_RBN2590_n_14460) );
no02f80 g757966 ( .a(n_22737), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_22788) );
no02f80 g741332 ( .a(n_38805), .b(n_38816), .o(n_38857) );
oa12f80 g770484 ( .a(n_10472), .b(n_10481), .c(n_10471), .o(n_10530) );
no02f80 g751632 ( .a(n_28422), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_12_), .o(n_28439) );
no02f80 g743015 ( .a(n_46256), .b(delay_add_ln22_unr23_stage9_stallmux_q_8_), .o(n_36958) );
in01f80 newInst_2418 ( .a(newNet_2097), .o(newNet_2418) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_10_ ( .ck(newNet_2326), .d(n_40350), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_) );
in01f80 newInst_3503 ( .a(newNet_3458), .o(newNet_3503) );
na02f80 g777701 ( .a(n_3404), .b(FE_OCP_RBN3479_n_3006), .o(n_3511) );
na02f80 g763102 ( .a(n_17410), .b(n_17345), .o(n_17411) );
in01f80 FE_OCP_RBC3438_n_33750 ( .a(n_33750), .o(FE_OCP_RBN3438_n_33750) );
in01f80 newInst_2247 ( .a(newNet_2246), .o(newNet_2247) );
na02f80 g754209 ( .a(n_25974), .b(n_25973), .o(n_25975) );
no02f80 g743191 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_4_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_4_), .o(n_36923) );
na02f80 g746893 ( .a(n_33035), .b(delay_add_ln22_unr20_stage8_stallmux_q_16_), .o(n_33057) );
in01f80 g737623 ( .a(n_42398), .o(n_42399) );
ao12f80 g779443 ( .a(n_1878), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_18_), .o(n_1917) );
no02f80 g777799 ( .a(n_3252), .b(n_3223), .o(n_3338) );
in01f80 g761963 ( .a(n_18301), .o(n_18346) );
no02f80 g746887 ( .a(n_33108), .b(n_32283), .o(n_33253) );
na02f80 g746201 ( .a(n_33622), .b(n_33184), .o(n_33623) );
na02f80 g737704 ( .a(n_42285), .b(n_41956), .o(n_42332) );
oa12f80 g770432 ( .a(n_10578), .b(n_10577), .c(n_10576), .o(n_10632) );
no02f80 g767069 ( .a(n_13623), .b(n_13640), .o(n_13682) );
na02f80 g736977 ( .a(FE_OCPN913_n_43022), .b(n_43299), .o(n_43393) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_12_ ( .ck(newNet_3340), .d(n_31996), .o(delay_add_ln22_unr20_stage8_stallmux_q_12_) );
in01f80 fopt782900 ( .a(n_2308), .o(n_44344) );
na02f80 g736809 ( .a(n_43424), .b(n_43429), .o(n_43462) );
in01f80 g770396 ( .a(n_10445), .o(n_10446) );
in01f80 g749167 ( .a(n_30978), .o(n_30979) );
in01f80 newInst_1720 ( .a(newNet_1719), .o(newNet_1720) );
in01f80 g770291 ( .a(n_10667), .o(n_10694) );
na02f80 g750139 ( .a(n_29813), .b(n_29812), .o(n_29872) );
oa12f80 g778192 ( .a(n_2700), .b(n_2699), .c(n_2698), .o(n_3494) );
in01f80 FE_RC_3696_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_4_), .o(FE_RN_1625_0) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_8_ ( .ck(newNet_481), .d(n_22832), .o(delay_xor_ln22_unr15_stage6_stallmux_q_8_) );
in01f80 g739917 ( .a(n_40297), .o(n_40379) );
in01f80 g741259 ( .a(n_39226), .o(n_39227) );
in01f80 FE_OCPC3774_n_14730 ( .a(n_14730), .o(FE_OCPN3774_n_14730) );
na02f80 g751842 ( .a(n_29123), .b(n_28897), .o(n_29126) );
no02f80 g778520 ( .a(n_2484), .b(n_2483), .o(n_2541) );
in01f80 g779288 ( .a(n_1766), .o(n_1767) );
in01f80 g743859 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_7_), .o(n_35713) );
in01f80 g761783 ( .a(n_18850), .o(n_18851) );
in01f80 newInst_3240 ( .a(newNet_3239), .o(newNet_3240) );
in01f80 newInst_1227 ( .a(newNet_1226), .o(newNet_1227) );
no02f80 g748321 ( .a(n_32197), .b(n_31703), .o(n_31840) );
in01f80 FE_OCP_RBC3547_n_44575 ( .a(n_44575), .o(FE_OCP_RBN3547_n_44575) );
na02f80 g772932 ( .a(n_7875), .b(n_7874), .o(n_7984) );
in01f80 g764211 ( .a(n_16818), .o(n_16819) );
in01f80 g748960 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_46101) );
no02f80 g757907 ( .a(n_22471), .b(n_22441), .o(n_22529) );
oa12f80 g775321 ( .a(n_5864), .b(n_5863), .c(n_5862), .o(n_5922) );
na02f80 g750420 ( .a(n_29569), .b(FE_OCPN1406_n_25859), .o(n_29624) );
in01f80 FE_RC_2134_0 ( .a(n_23486), .o(FE_RN_746_0) );
in01f80 newInst_2025 ( .a(newNet_2024), .o(newNet_2025) );
na02f80 g770375 ( .a(n_10535), .b(n_10506), .o(n_10571) );
oa12f80 g742382 ( .a(n_37766), .b(n_37765), .c(n_37764), .o(n_38738) );
in01f80 g760637 ( .a(n_21246), .o(n_20327) );
oa12f80 g761742 ( .a(n_18745), .b(n_18789), .c(n_18744), .o(n_18852) );
no02f80 g776534 ( .a(n_4413), .b(n_4448), .o(n_4643) );
in01f80 FE_OCP_RBC3560_n_8809 ( .a(n_8809), .o(FE_OCP_RBN3560_n_8809) );
ao12f80 g747135 ( .a(n_32814), .b(n_32885), .c(n_32845), .o(n_32931) );
ao22s80 FE_RC_808_0 ( .a(n_7736), .b(n_8914), .c(n_7735), .d(n_8921), .o(n_9057) );
ao12f80 g746873 ( .a(n_32971), .b(n_32994), .c(n_32970), .o(n_33907) );
no02f80 g743974 ( .a(n_47267), .b(n_36035), .o(n_36069) );
in01f80 g780040 ( .a(n_1250), .o(n_1251) );
no02f80 g764735 ( .a(n_15735), .b(n_15702), .o(n_15799) );
na02f80 FE_RC_3488_0 ( .a(FE_RN_1502_0), .b(n_37380), .o(n_37377) );
in01f80 g768363 ( .a(n_12483), .o(n_12484) );
no02f80 g755065 ( .a(n_25319), .b(n_25229), .o(n_25354) );
ao12f80 g780694 ( .a(n_644), .b(n_647), .c(n_643), .o(n_867) );
in01f80 g774325 ( .a(n_6644), .o(n_6645) );
na02f80 g769885 ( .a(n_11091), .b(n_11075), .o(n_11177) );
na02f80 FE_RC_2069_0 ( .a(n_24919), .b(n_24860), .o(FE_RN_704_0) );
no02f80 g772717 ( .a(n_8148), .b(n_8132), .o(n_8229) );
oa12f80 g778927 ( .a(n_1781), .b(n_2148), .c(n_1722), .o(n_2169) );
na02f80 g742978 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_14_), .o(n_36973) );
oa12f80 g756374 ( .a(n_23503), .b(n_23691), .c(n_23481), .o(n_23827) );
na02f80 FE_RC_2543_0 ( .a(n_38902), .b(n_39260), .o(FE_RN_1040_0) );
in01f80 g776980 ( .a(n_4087), .o(n_4088) );
in01f80 g752294 ( .a(n_28028), .o(n_28029) );
in01f80 FE_RC_3760_0 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_6_), .o(FE_RN_1651_0) );
in01f80 newInst_3544 ( .a(newNet_3543), .o(newNet_3544) );
no02f80 g761138 ( .a(n_19150), .b(n_18821), .o(n_19173) );
no02f80 g752279 ( .a(FE_OCPN877_n_44734), .b(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .o(n_27968) );
na02f80 g756250 ( .a(n_24122), .b(n_23776), .o(n_24139) );
na02f80 g753401 ( .a(n_27068), .b(n_27036), .o(n_27081) );
na02f80 g781064 ( .a(cos_out_15), .b(FE_OFN2_n_43918), .o(n_350) );
na02f80 g743701 ( .a(n_36344), .b(n_35868), .o(n_36408) );
ao22s80 FE_RC_1228_0 ( .a(n_7732), .b(n_8943), .c(n_7733), .d(n_8944), .o(n_9091) );
no02f80 g770805 ( .a(n_10111), .b(n_10092), .o(n_10179) );
na02f80 g775194 ( .a(n_5957), .b(n_5688), .o(n_5978) );
ao22s80 g739611 ( .a(FE_OCP_RBN3336_n_44610), .b(n_40607), .c(n_44610), .d(delay_xor_ln21_unr28_stage10_stallmux_q_0_), .o(n_40638) );
in01f80 newInst_632 ( .a(newNet_631), .o(newNet_632) );
oa22f80 FE_RC_963_0 ( .a(n_32126), .b(n_32349), .c(n_32127), .d(n_32366), .o(n_32518) );
in01f80 FE_RC_2252_0 ( .a(n_17308), .o(FE_RN_830_0) );
oa12f80 g756287 ( .a(n_23705), .b(n_24586), .c(n_23908), .o(n_24734) );
in01f80 g761746 ( .a(n_18605), .o(n_18712) );
no02f80 g766310 ( .a(n_14333), .b(n_14270), .o(n_14370) );
in01f80 g766893 ( .a(n_14425), .o(n_14388) );
in01f80 g780414 ( .a(n_1208), .o(n_1122) );
ao12f80 g746567 ( .a(n_34815), .b(n_34810), .c(n_34497), .o(n_35042) );
na02f80 g756781 ( .a(n_23956), .b(n_24034), .o(n_24035) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_28_ ( .ck(newNet_1381), .d(n_36726), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_28_) );
ao12f80 g780780 ( .a(n_454), .b(n_430), .c(n_470), .o(n_456) );
in01f80 g737759 ( .a(n_42353), .o(n_42354) );
in01f80 fopt784010 ( .a(n_32680), .o(n_45741) );
no02f80 g763802 ( .a(n_17423), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_23_), .o(n_17465) );
in01f80 FE_OCPC1031_n_28448 ( .a(n_28448), .o(FE_OCPN1031_n_28448) );
no02f80 g737174 ( .a(n_43003), .b(n_43002), .o(n_43004) );
na02f80 g773407 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_27_), .o(n_7557) );
in01f80 g738380 ( .a(n_41515), .o(n_41516) );
na02f80 g766833 ( .a(n_13907), .b(n_14215), .o(n_14525) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_27_ ( .ck(newNet_1825), .d(n_17058), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_27_) );
in01f80 FE_OCP_RBC3721_n_39913 ( .a(FE_OCP_RBN3720_n_39913), .o(FE_OCP_RBN3721_n_39913) );
no02f80 g754139 ( .a(n_25966), .b(n_25588), .o(n_26069) );
in01f80 g741609 ( .a(n_38657), .o(n_38686) );
ao12f80 g764989 ( .a(n_15581), .b(n_15644), .c(n_15643), .o(n_15752) );
na02f80 g741045 ( .a(n_39243), .b(n_39303), .o(n_39329) );
na02f80 g781128 ( .a(n_222), .b(n_75), .o(n_224) );
ao12f80 g772871 ( .a(n_7940), .b(n_7939), .c(n_7938), .o(n_8024) );
in01f80 g775757 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_8_), .o(n_5430) );
no02f80 g737195 ( .a(FE_OCP_RBN2914_n_42947), .b(n_43012), .o(n_42978) );
in01f80 g760317 ( .a(n_20325), .o(n_20326) );
in01f80 newInst_2700 ( .a(newNet_1174), .o(newNet_2700) );
in01f80 g775909 ( .a(n_5364), .o(n_5400) );
in01f80 g755071 ( .a(n_25533), .o(n_25534) );
no02f80 g749274 ( .a(n_30676), .b(n_30373), .o(n_30739) );
in01f80 g741827 ( .a(n_39324), .o(n_38467) );
in01f80 newInst_1656 ( .a(newNet_1655), .o(newNet_1656) );
in01f80 g752435 ( .a(n_28397), .o(n_28398) );
na02f80 g744750 ( .a(n_35107), .b(n_35106), .o(n_35121) );
in01f80 g757103 ( .a(n_23178), .o(n_23179) );
in01f80 g743455 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_31_), .o(n_36650) );
ao12f80 g752475 ( .a(n_28052), .b(n_28328), .c(n_27905), .o(n_28401) );
na02f80 g755854 ( .a(n_24340), .b(n_23822), .o(n_24396) );
no02f80 g767709 ( .a(n_46414), .b(n_13127), .o(n_13211) );
in01f80 newInst_1293 ( .a(newNet_1292), .o(newNet_1293) );
in01f80 g771439 ( .a(n_9163), .o(n_9210) );
in01f80 g746237 ( .a(n_33820), .o(n_34006) );
in01f80 newInst_1648 ( .a(newNet_1647), .o(newNet_1648) );
in01f80 FE_OCP_RBC2687_n_38870 ( .a(FE_OCP_RBN2685_n_38870), .o(FE_OCP_RBN2687_n_38870) );
no02f80 g751163 ( .a(n_30303), .b(n_29908), .o(n_30381) );
no02f80 g752739 ( .a(n_28152), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_30_), .o(n_28178) );
in01f80 newInst_3427 ( .a(newNet_3426), .o(newNet_3427) );
in01f80 g741096 ( .a(n_39362), .o(n_39363) );
in01f80 newInst_1154 ( .a(newNet_1153), .o(newNet_1154) );
in01f80 g773461 ( .a(n_7513), .o(n_7514) );
no02f80 g740276 ( .a(n_40097), .b(n_39576), .o(n_40098) );
in01f80 g736699 ( .a(n_43329), .o(n_43330) );
na02f80 FE_RC_2550_0 ( .a(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .b(n_33976), .o(FE_RN_1044_0) );
in01f80 g780232 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_2_), .o(n_1107) );
na02f80 g778622 ( .a(n_2544), .b(n_2571), .o(n_2603) );
na02f80 g775952 ( .a(n_5141), .b(n_4658), .o(n_5217) );
in01f80 g749518 ( .a(n_31909), .o(n_31910) );
na02f80 g742313 ( .a(n_37819), .b(n_37818), .o(n_37820) );
in01f80 g748875 ( .a(n_32418), .o(n_32419) );
in01f80 g765070 ( .a(n_15529), .o(n_15641) );
no02f80 g777963 ( .a(n_3092), .b(n_2286), .o(n_3093) );
in01f80 g773994 ( .a(n_6990), .o(n_6991) );
na02f80 g741321 ( .a(FE_OCP_RBN2546_n_44944), .b(FE_OCP_RBN2452_n_38537), .o(n_39126) );
in01f80 fopt783491 ( .a(n_45066), .o(n_45067) );
na02f80 g774010 ( .a(n_6897), .b(n_6896), .o(n_6898) );
na02f80 g764381 ( .a(n_16364), .b(n_16436), .o(n_16388) );
no02f80 g744810 ( .a(n_35194), .b(FE_OCP_RBN2712_n_35075), .o(n_35195) );
in01f80 g737695 ( .a(n_42260), .o(n_42540) );
ao22s80 g737872 ( .a(FE_OCPN1232_n_42201), .b(n_42209), .c(n_42270), .d(n_42267), .o(n_42507) );
oa12f80 g766708 ( .a(n_13753), .b(n_13805), .c(n_13853), .o(n_14064) );
na02f80 g776214 ( .a(n_4889), .b(n_4876), .o(n_5063) );
in01f80 newInst_369 ( .a(newNet_368), .o(newNet_369) );
in01f80 FE_OCP_RBC1710_n_22150 ( .a(FE_OCP_RBN1709_n_22150), .o(FE_OCP_RBN1710_n_22150) );
na02f80 FE_RC_1337_0 ( .a(FE_RN_398_0), .b(n_5279), .o(n_47002) );
na02f80 g752704 ( .a(n_27244), .b(n_27243), .o(n_27245) );
in01f80 g775941 ( .a(n_4922), .o(n_4923) );
no02f80 g738683 ( .a(n_41525), .b(n_41297), .o(n_41722) );
no02f80 g744754 ( .a(n_35284), .b(n_35250), .o(n_35303) );
in01f80 FE_OCP_RBC2495_n_8641 ( .a(FE_OCP_RBN2494_n_8641), .o(FE_OCP_RBN2495_n_8641) );
no02f80 g763804 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_22_), .o(n_17358) );
in01f80 FE_OCPC846_n_4046 ( .a(FE_OCPN845_n_4046), .o(FE_OCPN846_n_4046) );
no02f80 g741407 ( .a(n_38800), .b(FE_OCPN3174_n_38799), .o(n_38816) );
no02f80 g736842 ( .a(n_43013), .b(n_43016), .o(n_43028) );
no02f80 g749947 ( .a(n_30470), .b(FE_OCP_RBN2632_n_30170), .o(n_30239) );
in01f80 g776990 ( .a(n_5403), .o(n_5404) );
oa22f80 FE_RC_2514_0 ( .a(n_30367), .b(n_31001), .c(n_30368), .d(n_31002), .o(n_31107) );
no02f80 g753970 ( .a(n_26318), .b(n_23590), .o(n_26354) );
na02f80 g739855 ( .a(n_40380), .b(n_40067), .o(n_40431) );
na02f80 g745969 ( .a(n_33946), .b(n_33945), .o(n_33966) );
no02f80 g744073 ( .a(n_44222), .b(n_35006), .o(n_36036) );
no02f80 g738831 ( .a(n_41656), .b(n_41562), .o(n_41328) );
no02f80 g765503 ( .a(n_15565), .b(n_15631), .o(n_15566) );
no02f80 g737519 ( .a(n_42381), .b(n_42336), .o(n_42475) );
in01f80 g750050 ( .a(n_30383), .o(n_30384) );
in01f80 g753752 ( .a(delay_sub_ln23_0_unr20_stage7_stallmux_q_13_), .o(n_27164) );
no02f80 g764467 ( .a(n_16155), .b(n_16112), .o(n_16366) );
oa22f80 g776899 ( .a(n_3814), .b(n_3029), .c(n_3746), .d(n_3862), .o(n_4028) );
in01f80 newInst_2119 ( .a(newNet_2118), .o(newNet_2119) );
no02f80 g754714 ( .a(FE_OCP_RBN2959_n_26231), .b(n_26510), .o(n_26551) );
in01f80 g779272 ( .a(n_1755), .o(n_1756) );
na02f80 g760149 ( .a(FE_OCP_RBN2740_n_20565), .b(n_20628), .o(n_20665) );
in01f80 g769306 ( .a(n_11509), .o(n_11924) );
in01f80 g751047 ( .a(n_29879), .o(n_29880) );
no02f80 g753762 ( .a(n_26458), .b(n_23509), .o(n_26579) );
no02f80 g754511 ( .a(n_26712), .b(n_26740), .o(n_26713) );
in01f80 g776660 ( .a(n_4131), .o(n_4057) );
no02f80 g743744 ( .a(n_37295), .b(n_36899), .o(n_37405) );
ao12f80 g780723 ( .a(n_613), .b(n_612), .c(n_611), .o(n_809) );
no02f80 g750946 ( .a(n_28935), .b(n_28550), .o(n_28976) );
oa12f80 g754305 ( .a(n_25536), .b(n_25819), .c(n_25556), .o(n_25900) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_0_ ( .ck(newNet_3461), .d(n_26150), .o(delay_add_ln22_unr17_stage7_stallmux_q_0_) );
ao12f80 g748737 ( .a(n_31230), .b(n_31353), .c(n_31296), .o(n_31399) );
in01f80 g754730 ( .a(n_26712), .o(n_26677) );
in01f80 newInst_2838 ( .a(newNet_2837), .o(newNet_2838) );
in01f80 g769615 ( .a(n_11384), .o(n_11385) );
no02f80 g736643 ( .a(n_43094), .b(n_43066), .o(n_43193) );
in01f80 FE_RC_3507_0 ( .a(FE_OFN787_n_25834), .o(FE_RN_1515_0) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_12_ ( .ck(newNet_3449), .d(n_27278), .o(delay_add_ln22_unr17_stage7_stallmux_q_12_) );
in01f80 g776012 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_), .o(n_5103) );
oa12f80 g770627 ( .a(n_10165), .b(n_10256), .c(n_10169), .o(n_10498) );
no02f80 g741055 ( .a(n_38986), .b(n_39103), .o(n_39415) );
ao12f80 g773780 ( .a(n_7189), .b(n_7188), .c(n_7187), .o(n_7240) );
in01f80 FE_OCP_RBC2272_n_13489 ( .a(FE_OCP_RBN2270_n_13489), .o(FE_OCP_RBN2272_n_13489) );
no02f80 g736918 ( .a(FE_OCPN910_n_43022), .b(n_42730), .o(n_43449) );
oa22f80 g761843 ( .a(n_18553), .b(n_16931), .c(n_18397), .d(n_18404), .o(n_20293) );
ao12f80 g767503 ( .a(n_12502), .b(n_12904), .c(n_12522), .o(n_13009) );
no02f80 g777168 ( .a(n_4362), .b(n_4576), .o(n_5261) );
oa12f80 g774130 ( .a(n_6655), .b(n_6654), .c(delay_add_ln22_unr5_stage3_stallmux_q_0_), .o(n_7286) );
in01f80 g742080 ( .a(n_38311), .o(n_38312) );
na02f80 g740450 ( .a(n_39769), .b(n_39768), .o(n_39806) );
ao12f80 g752452 ( .a(n_27294), .b(n_45638), .c(n_27211), .o(n_27697) );
oa12f80 g749414 ( .a(n_31572), .b(n_31911), .c(n_31321), .o(n_31977) );
in01f80 g749523 ( .a(n_30530), .o(n_30508) );
no02f80 g753633 ( .a(n_27284), .b(n_26714), .o(n_27321) );
in01f80 g758297 ( .a(n_22465), .o(n_22406) );
in01f80 FE_OFC754_n_44461 ( .a(FE_OCP_RBN2616_n_44561), .o(FE_OFN754_n_44461) );
oa12f80 g776955 ( .a(n_3986), .b(n_3985), .c(n_3984), .o(n_4089) );
no02f80 g750711 ( .a(n_29220), .b(n_29240), .o(n_29477) );
na02f80 g742595 ( .a(n_37429), .b(n_37428), .o(n_37430) );
na03f80 g765018 ( .a(n_16384), .b(n_16261), .c(n_16258), .o(n_16262) );
oa22f80 g744526 ( .a(n_36664), .b(n_36162), .c(n_36665), .d(n_36161), .o(n_36714) );
in01f80 g764357 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_11_), .o(n_18055) );
na02f80 g751533 ( .a(n_28460), .b(n_27833), .o(n_28786) );
in01f80 g766182 ( .a(n_14573), .o(n_14595) );
no02f80 g776926 ( .a(n_3996), .b(n_3912), .o(n_4222) );
in01f80 FE_OCP_RBC2177_n_1864 ( .a(n_1864), .o(FE_OCP_RBN2177_n_1864) );
oa12f80 g736286 ( .a(n_324), .b(n_43858), .c(FE_OFN3_n_43918), .o(n_43890) );
oa12f80 g749650 ( .a(n_30249), .b(n_30248), .c(n_30247), .o(n_30324) );
in01f80 g749268 ( .a(n_30800), .o(n_30801) );
in01f80 g750824 ( .a(n_29116), .o(n_29117) );
no02f80 g775783 ( .a(n_5501), .b(n_5534), .o(n_5535) );
na02f80 g759467 ( .a(n_20915), .b(n_20914), .o(n_20916) );
na02f80 g779560 ( .a(FE_OCP_RBN3249_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_1_), .o(n_1376) );
in01f80 g756515 ( .a(n_23844), .o(n_23845) );
ao12f80 g745870 ( .a(n_33923), .b(n_34017), .c(n_33963), .o(n_34069) );
no02f80 g773490 ( .a(n_7496), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_23_), .o(n_7502) );
in01f80 FE_OCP_RBC2936_n_10626 ( .a(n_10626), .o(FE_OCP_RBN2936_n_10626) );
in01f80 newInst_3378 ( .a(newNet_3377), .o(newNet_3378) );
no02f80 g738746 ( .a(n_41367), .b(n_41366), .o(n_41368) );
in01f80 FE_OCP_DRV_C1561_n_19562 ( .a(n_19562), .o(FE_OCP_DRV_N1561_n_19562) );
in01f80 FE_RC_2651_0 ( .a(FE_RN_1106_0), .o(n_12590) );
na02f80 g753823 ( .a(n_26320), .b(n_23467), .o(n_26478) );
na02f80 g736684 ( .a(n_43469), .b(n_43472), .o(n_43562) );
in01f80 g749821 ( .a(n_31564), .o(n_31565) );
oa12f80 g768616 ( .a(n_12203), .b(n_12202), .c(n_12201), .o(n_12289) );
na02f80 g756496 ( .a(n_23822), .b(n_23675), .o(n_23846) );
no02f80 g751604 ( .a(FE_OCP_RBN3404_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_28_), .o(n_28801) );
in01f80 g768477 ( .a(n_12454), .o(n_12455) );
oa12f80 g756840 ( .a(n_23336), .b(n_23385), .c(n_23335), .o(n_23476) );
in01f80 g778237 ( .a(n_2799), .o(n_3034) );
na02f80 g775535 ( .a(n_5454), .b(n_4759), .o(n_5488) );
na02f80 g737370 ( .a(n_42808), .b(n_42769), .o(n_42861) );
in01f80 g756138 ( .a(n_24981), .o(n_24998) );
na02f80 g751703 ( .a(n_28366), .b(n_28365), .o(n_28421) );
in01f80 newInst_216 ( .a(newNet_215), .o(newNet_216) );
no02f80 g772242 ( .a(n_8777), .b(n_8069), .o(n_8856) );
in01f80 fopt784024 ( .a(n_29371), .o(n_45760) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_19_ ( .ck(newNet_2764), .d(n_46973), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_19_) );
no02f80 g750667 ( .a(n_29301), .b(n_29323), .o(n_30192) );
na02f80 g766656 ( .a(n_13980), .b(n_13945), .o(n_14015) );
no02f80 g740599 ( .a(n_39575), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39595) );
no02f80 g781130 ( .a(n_222), .b(n_160), .o(n_216) );
no02f80 g742104 ( .a(n_37880), .b(n_37890), .o(n_37944) );
in01f80 g741665 ( .a(n_38609), .o(n_38610) );
in01f80 g750016 ( .a(n_30273), .o(n_30274) );
in01f80 newInst_3720 ( .a(newNet_867), .o(newNet_3720) );
in01f80 g745786 ( .a(FE_OFN627_n_34445), .o(n_34446) );
no02f80 g741021 ( .a(n_39132), .b(n_38870), .o(n_39209) );
na02f80 g738873 ( .a(n_41273), .b(n_41272), .o(n_41274) );
in01f80 g737013 ( .a(n_43451), .o(n_43452) );
in01f80 g757680 ( .a(n_22715), .o(n_22670) );
oa12f80 g770770 ( .a(n_10238), .b(n_10255), .c(n_10237), .o(n_10301) );
in01f80 g743861 ( .a(n_37898), .o(n_37189) );
in01f80 g753890 ( .a(n_26325), .o(n_26326) );
na02f80 g775741 ( .a(n_5335), .b(n_4163), .o(n_5336) );
no02f80 g752190 ( .a(n_28037), .b(n_28036), .o(n_28038) );
na02f80 g761962 ( .a(n_18357), .b(n_18393), .o(n_18396) );
in01f80 g746357 ( .a(n_33503), .o(n_33523) );
no02f80 g750923 ( .a(n_30105), .b(n_30104), .o(n_30106) );
na02f80 g746884 ( .a(FE_OCP_RBN3387_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_29_), .o(n_33325) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_14_ ( .ck(newNet_1027), .d(n_17829), .o(delay_xor_ln21_unr12_stage5_stallmux_q_14_) );
in01f80 FE_OCP_RBC3527_n_13765 ( .a(FE_OCP_RBN2459_n_13765), .o(FE_OCP_RBN3527_n_13765) );
na02f80 g770150 ( .a(n_10788), .b(n_10714), .o(n_10861) );
in01f80 newInst_3571 ( .a(newNet_3570), .o(newNet_3571) );
in01f80 newInst_197 ( .a(newNet_196), .o(newNet_197) );
na02f80 g740507 ( .a(n_39698), .b(n_38786), .o(n_39717) );
in01f80 FE_OCP_RBC2199_n_2032 ( .a(n_2032), .o(FE_OCP_RBN2199_n_2032) );
oa22f80 FE_RC_1705_0 ( .a(n_21306), .b(n_21262), .c(n_21261), .d(n_21307), .o(n_21494) );
oa12f80 g750388 ( .a(n_30617), .b(n_30634), .c(n_30616), .o(n_31184) );
in01f80 g751997 ( .a(n_29023), .o(n_29024) );
na02f80 g770513 ( .a(n_10280), .b(n_10282), .o(n_10412) );
in01f80 newInst_1290 ( .a(newNet_1289), .o(newNet_1290) );
in01f80 g762992 ( .a(n_17494), .o(n_17599) );
in01f80 g751655 ( .a(n_28467), .o(n_28460) );
na02f80 g769225 ( .a(n_11474), .b(n_11538), .o(n_11587) );
na02f80 g768079 ( .a(FE_OCPN860_n_12880), .b(n_12290), .o(n_12994) );
na02f80 g748305 ( .a(n_31793), .b(n_31862), .o(n_31895) );
oa22f80 g758739 ( .a(n_21805), .b(n_21631), .c(n_21804), .d(n_21630), .o(n_21946) );
na02f80 g780166 ( .a(n_1075), .b(n_1074), .o(n_1076) );
na02f80 g770766 ( .a(n_10334), .b(n_10302), .o(n_10303) );
no02f80 g753759 ( .a(n_26407), .b(n_26433), .o(n_26449) );
no02f80 g741983 ( .a(n_38062), .b(n_37980), .o(n_38014) );
na02f80 g772580 ( .a(n_8352), .b(n_8351), .o(n_8353) );
in01f80 newInst_375 ( .a(newNet_374), .o(newNet_375) );
no02f80 g776190 ( .a(n_4954), .b(n_4953), .o(n_4980) );
na02f80 FE_RC_70_0 ( .a(FE_RN_18_0), .b(FE_RN_19_0), .o(FE_RN_20_0) );
in01f80 g752826 ( .a(n_27402), .o(n_27430) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_4_ ( .ck(newNet_2521), .d(n_26693), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_) );
in01f80 newInst_1671 ( .a(newNet_270), .o(newNet_1671) );
in01f80 g755474 ( .a(n_24655), .o(n_24726) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_22_ ( .ck(newNet_1509), .d(n_32248), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_22_) );
in01f80 FE_RC_640_0 ( .a(n_28575), .o(FE_RN_202_0) );
na03f80 FE_RC_2615_0 ( .a(n_14511), .b(FE_RN_1087_0), .c(FE_RN_1088_0), .o(FE_RN_1089_0) );
ao12f80 g756084 ( .a(n_23713), .b(n_24145), .c(n_23768), .o(n_24166) );
ao12f80 g762812 ( .a(n_18085), .b(n_18084), .c(n_18083), .o(n_18448) );
in01f80 newInst_2097 ( .a(newNet_1360), .o(newNet_2097) );
in01f80 g738162 ( .a(n_42030), .o(n_42029) );
in01f80 g746986 ( .a(n_32934), .o(n_32935) );
in01f80 g742415 ( .a(n_37757), .o(n_37758) );
na02f80 g749717 ( .a(n_31481), .b(FE_OCP_RBN3011_n_31117), .o(n_31540) );
in01f80 newInst_3058 ( .a(newNet_3057), .o(newNet_3058) );
no02f80 FE_RC_2781_0 ( .a(n_19561), .b(n_19639), .o(FE_RN_1187_0) );
na02f80 g766835 ( .a(n_13743), .b(n_13800), .o(n_13704) );
in01f80 g769486 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11507) );
in01f80 g769722 ( .a(n_11225), .o(n_11226) );
oa12f80 g780936 ( .a(n_377), .b(n_376), .c(n_200), .o(n_378) );
in01f80 g772248 ( .a(n_8794), .o(n_8858) );
no02f80 g753833 ( .a(n_26326), .b(n_26403), .o(n_26479) );
na02f80 g740281 ( .a(n_40239), .b(n_40309), .o(n_40361) );
ao12f80 g762935 ( .a(n_17639), .b(n_17717), .c(n_17715), .o(n_17839) );
na02f80 g781011 ( .a(cos_out_0), .b(FE_OFN5_n_43918), .o(n_317) );
na02f80 g746613 ( .a(FE_OCP_RBN2598_n_34388), .b(n_33911), .o(n_34498) );
in01f80 g746054 ( .a(n_33976), .o(n_34004) );
in01f80 g762678 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_31_), .o(n_17852) );
no02f80 FE_RC_1883_0 ( .a(n_28086), .b(delay_add_ln22_unr17_stage7_stallmux_q_4_), .o(FE_RN_585_0) );
no02f80 g770839 ( .a(n_9807), .b(n_9750), .o(n_9858) );
in01f80 g778717 ( .a(n_2245), .o(n_2293) );
in01f80 newInst_2621 ( .a(newNet_2620), .o(newNet_2621) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_7_ ( .ck(newNet_2610), .d(n_21613), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_7_) );
in01f80 FE_OCP_RBC2669_n_4158 ( .a(FE_OCP_RBN2668_n_4158), .o(FE_OCP_RBN2669_n_4158) );
no02f80 g769336 ( .a(FE_OCP_RBN1993_delay_sub_ln23_0_unr8_stage4_stallmux_q_0_), .b(n_45224), .o(n_11640) );
no02f80 g780430 ( .a(n_688), .b(n_676), .o(n_739) );
no02f80 g743402 ( .a(n_36670), .b(n_36687), .o(n_36730) );
na02f80 g741191 ( .a(FE_OCP_RBN3625_n_38870), .b(n_39393), .o(n_39487) );
no02f80 g740795 ( .a(n_39314), .b(n_39313), .o(n_39355) );
in01f80 FE_OCPC915_n_7832 ( .a(FE_OCPN914_n_7832), .o(FE_OCPN915_n_7832) );
no02f80 g745189 ( .a(n_34601), .b(n_34600), .o(n_34602) );
in01f80 g754740 ( .a(n_26383), .o(n_26343) );
no02f80 g761941 ( .a(n_18268), .b(n_17555), .o(n_18398) );
na02f80 g779404 ( .a(n_1510), .b(n_1485), .o(n_1556) );
in01f80 g757956 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_12_), .o(n_23475) );
ao12f80 g761289 ( .a(n_19651), .b(n_19709), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_19769) );
in01f80 newInst_2751 ( .a(newNet_2750), .o(newNet_2751) );
no02f80 g752001 ( .a(n_28919), .b(n_28984), .o(n_29002) );
na02f80 g765644 ( .a(n_15005), .b(n_14920), .o(n_15040) );
na02f80 g781218 ( .a(n_165), .b(beta_3), .o(n_166) );
no02f80 g749119 ( .a(n_30882), .b(FE_OCP_RBN2378_n_29480), .o(n_30883) );
no02f80 g773547 ( .a(n_7442), .b(n_7441), .o(n_7443) );
in01f80 newInst_2969 ( .a(newNet_1939), .o(newNet_2969) );
na02f80 g748592 ( .a(n_32658), .b(n_32500), .o(n_32674) );
na02f80 g754103 ( .a(n_26039), .b(n_23353), .o(n_26175) );
ao12f80 g772691 ( .a(n_7349), .b(n_8106), .c(n_7382), .o(n_8191) );
in01f80 g762249 ( .a(n_18696), .o(n_18697) );
in01f80 g767018 ( .a(n_13864), .o(n_13823) );
no02f80 g779621 ( .a(n_1852), .b(delay_xor_ln22_unr3_stage2_stallmux_q_19_), .o(n_1930) );
oa22f80 g756447 ( .a(n_23602), .b(n_23537), .c(n_23666), .d(n_23538), .o(n_25044) );
no02f80 g756588 ( .a(n_23783), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_), .o(n_23851) );
no02f80 FE_RC_2924_0 ( .a(FE_RN_1272_0), .b(n_27087), .o(FE_RN_1273_0) );
in01f80 newInst_3283 ( .a(newNet_2694), .o(newNet_3283) );
na02f80 g739278 ( .a(n_40893), .b(n_40809), .o(n_40851) );
na02f80 g740242 ( .a(n_39854), .b(n_39853), .o(n_39893) );
ao12f80 g764974 ( .a(n_16312), .b(n_16176), .c(FE_OFN764_n_15670), .o(n_16313) );
no02f80 g784795 ( .a(n_6565), .b(n_6415), .o(n_47334) );
ao12f80 g739382 ( .a(n_40808), .b(n_40709), .c(n_40645), .o(n_40892) );
in01f80 newInst_3666 ( .a(newNet_3665), .o(newNet_3666) );
oa22f80 g784356 ( .a(FE_OFN775_n_46137), .b(n_5567), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5618), .o(n_46162) );
in01f80 g765194 ( .a(n_16063), .o(n_16064) );
no02f80 g772737 ( .a(n_8204), .b(n_8192), .o(n_8193) );
na02f80 g751756 ( .a(n_28306), .b(n_28305), .o(n_28344) );
na02f80 g770122 ( .a(n_10951), .b(n_10942), .o(n_10943) );
na02f80 g764961 ( .a(n_15503), .b(n_15502), .o(n_15543) );
no02f80 g742148 ( .a(FE_OCP_RBN3444_n_37945), .b(n_37568), .o(n_38111) );
no02f80 g760919 ( .a(n_19445), .b(n_17881), .o(n_19501) );
in01f80 newInst_2046 ( .a(newNet_2045), .o(newNet_2046) );
na02f80 g750691 ( .a(n_29217), .b(FE_RN_1513_0), .o(n_29241) );
in01f80 g780228 ( .a(n_1028), .o(n_1066) );
na02f80 g760823 ( .a(n_19517), .b(n_19430), .o(n_19535) );
in01f80 g768955 ( .a(delay_sub_ln21_0_unr8_stage4_stallmux_q_22_), .o(n_13024) );
in01f80 FE_OCP_RBC2924_n_5130 ( .a(FE_OCP_RBN2923_n_5130), .o(FE_OCP_RBN2924_n_5130) );
in01f80 newInst_3350 ( .a(newNet_3349), .o(newNet_3350) );
in01f80 g755805 ( .a(n_25221), .o(n_25222) );
na02f80 g758239 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_24_), .o(n_22840) );
na02f80 g739218 ( .a(n_40790), .b(n_40702), .o(n_40703) );
oa12f80 g739096 ( .a(n_41003), .b(n_41002), .c(n_41001), .o(n_41402) );
na02f80 g739223 ( .a(n_44026), .b(n_40726), .o(n_40782) );
no02f80 g741268 ( .a(FE_OCP_RBN2546_n_44944), .b(n_39025), .o(n_39094) );
in01f80 FE_OCP_RBC3050_n_11329 ( .a(n_11329), .o(FE_OCP_RBN3050_n_11329) );
no02f80 g772797 ( .a(n_8136), .b(n_8135), .o(n_8216) );
na02f80 g740836 ( .a(n_39237), .b(n_39330), .o(n_39404) );
na02f80 g737061 ( .a(n_43046), .b(n_42910), .o(n_43125) );
no02f80 g749569 ( .a(n_30405), .b(n_30010), .o(n_30436) );
ao22s80 FE_RC_541_0 ( .a(n_25859), .b(FE_OCP_RBN2340_n_29470), .c(n_29470), .d(n_29630), .o(n_29594) );
in01f80 newInst_2406 ( .a(newNet_2405), .o(newNet_2406) );
oa22f80 g784360 ( .a(FE_OFN774_n_46137), .b(n_6254), .c(FE_OCP_RBN3077_FE_OFN807_n_46195), .d(n_6297), .o(n_46166) );
na02f80 g781050 ( .a(cos_out_20), .b(n_43918), .o(n_338) );
na02f80 g766946 ( .a(n_13794), .b(n_13848), .o(n_13869) );
in01f80 FE_OCP_RBC2255_n_37844 ( .a(n_37844), .o(FE_OCP_RBN2255_n_37844) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_3_ ( .ck(newNet_1958), .d(n_9958), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_3_) );
na02f80 g736653 ( .a(n_43440), .b(n_43365), .o(n_43565) );
na02f80 g764196 ( .a(n_16368), .b(n_16491), .o(n_16529) );
na02f80 g753227 ( .a(n_27204), .b(n_26169), .o(n_27339) );
na02f80 g760662 ( .a(n_19700), .b(n_19705), .o(n_19774) );
na02f80 g773764 ( .a(n_7222), .b(n_7082), .o(n_7220) );
no02f80 g756460 ( .a(n_24195), .b(n_24194), .o(n_24196) );
no02f80 g763594 ( .a(n_17374), .b(n_17496), .o(n_17432) );
ao12f80 g743770 ( .a(n_35669), .b(n_36324), .c(n_36304), .o(n_36338) );
in01f80 FE_OCPC967_n_19342 ( .a(n_19342), .o(FE_OCPN967_n_19342) );
na02f80 g749022 ( .a(n_31018), .b(n_30822), .o(n_31079) );
in01f80 g750058 ( .a(n_30010), .o(n_30011) );
no02f80 g766426 ( .a(n_14144), .b(n_13464), .o(n_14183) );
in01f80 FE_OCP_RBC2418_n_19601 ( .a(n_19601), .o(FE_OCP_RBN2418_n_19601) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_26_ ( .ck(newNet_3404), .d(n_27772), .o(delay_add_ln22_unr17_stage7_stallmux_q_26_) );
na02f80 g775398 ( .a(n_5775), .b(n_5774), .o(n_5776) );
no02f80 g779059 ( .a(n_2043), .b(n_2040), .o(n_2041) );
in01f80 g747045 ( .a(n_32863), .o(n_32857) );
in01f80 g769867 ( .a(n_11164), .o(n_11165) );
in01f80 newInst_828 ( .a(newNet_827), .o(newNet_828) );
oa12f80 g738452 ( .a(n_41748), .b(FE_OCPN952_n_41540), .c(n_41695), .o(n_42017) );
no02f80 g744831 ( .a(n_35138), .b(n_35117), .o(n_35219) );
oa12f80 g739191 ( .a(n_40820), .b(n_40892), .c(n_40728), .o(n_40938) );
ao12f80 g748117 ( .a(n_32458), .b(n_32778), .c(n_32484), .o(n_32841) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_29_ ( .ck(newNet_2923), .d(n_6627), .o(delay_add_ln22_unr5_stage3_stallmux_q_29_) );
no02f80 g741448 ( .a(n_38796), .b(n_38779), .o(n_38830) );
in01f80 g776385 ( .a(n_4197), .o(n_4271) );
in01f80 g763747 ( .a(n_16731), .o(n_16732) );
na02f80 g783826 ( .a(n_45512), .b(n_44610), .o(n_45513) );
oa12f80 g754002 ( .a(n_26953), .b(n_26952), .c(n_26951), .o(n_27002) );
in01f80 newInst_148 ( .a(newNet_81), .o(newNet_148) );
in01f80 g745333 ( .a(n_36213), .o(n_36214) );
in01f80 newInst_953 ( .a(newNet_952), .o(newNet_953) );
na02f80 g756437 ( .a(n_24112), .b(n_24110), .o(n_24155) );
no02f80 g776588 ( .a(n_3905), .b(n_3835), .o(n_3974) );
na02f80 g739231 ( .a(n_40829), .b(n_40790), .o(n_41160) );
oa22f80 g784362 ( .a(FE_OFN86_n_46137), .b(n_5935), .c(FE_OCP_RBN3075_FE_OFN807_n_46195), .d(n_5971), .o(n_46168) );
in01f80 g742544 ( .a(n_37577), .o(n_37595) );
in01f80 FE_RC_2281_0 ( .a(FE_RN_853_0), .o(n_44827) );
ao12f80 g774021 ( .a(n_7196), .b(n_7217), .c(delay_xor_ln22_unr6_stage3_stallmux_q_22_), .o(n_7250) );
na02f80 g739349 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_12_), .o(n_41007) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_3_ ( .ck(newNet_1933), .d(n_36830), .o(delay_sub_ln21_unr24_stage9_stallmux_q_3_) );
oa22f80 g743715 ( .a(n_36273), .b(n_36287), .c(n_36274), .d(n_36288), .o(n_36371) );
in01f80 g748440 ( .a(n_31499), .o(n_31500) );
in01f80 g736439 ( .a(n_43781), .o(n_43782) );
in01f80 g757702 ( .a(n_22635), .o(n_22614) );
na02f80 g763531 ( .a(FE_OCP_RBN3079_n_16977), .b(n_16089), .o(n_17113) );
na02f80 FE_RC_3126_0 ( .a(FE_RN_1385_0), .b(n_27167), .o(n_27206) );
in01f80 g742230 ( .a(n_38247), .o(n_38248) );
in01f80 g746458 ( .a(n_34122), .o(n_33499) );
ao12f80 g779808 ( .a(n_1517), .b(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_8_), .o(n_1539) );
oa12f80 g743200 ( .a(n_36802), .b(n_36847), .c(n_36875), .o(n_36910) );
in01f80 newInst_1805 ( .a(newNet_1804), .o(newNet_1805) );
oa12f80 g743776 ( .a(n_37260), .b(n_37283), .c(n_37259), .o(n_37292) );
na02f80 g750135 ( .a(n_29839), .b(FE_OCPN1478_n_28775), .o(n_29890) );
na02f80 g753176 ( .a(n_27204), .b(n_25822), .o(n_27506) );
no02f80 g738429 ( .a(n_41742), .b(n_41788), .o(n_41812) );
in01f80 FE_OCP_RBC1695_n_19206 ( .a(n_19206), .o(FE_OCP_RBN1695_n_19206) );
na02f80 g758520 ( .a(n_21953), .b(FE_OCP_RBN1364_n_20412), .o(n_21970) );
in01f80 g754566 ( .a(n_26736), .o(n_26737) );
na02f80 g742457 ( .a(n_37665), .b(n_37647), .o(n_37762) );
oa12f80 g775426 ( .a(n_4820), .b(n_5741), .c(n_4901), .o(n_5860) );
no02f80 g772788 ( .a(n_8077), .b(n_7721), .o(n_8078) );
no02f80 g741855 ( .a(n_38363), .b(n_38362), .o(n_38364) );
no02f80 g742234 ( .a(FE_OCP_RBN2241_n_44881), .b(n_38290), .o(n_38373) );
oa22f80 g764230 ( .a(n_16798), .b(n_15959), .c(n_16770), .d(n_15960), .o(n_16846) );
in01f80 g742630 ( .a(n_37449), .o(n_37450) );
no02f80 g747634 ( .a(n_32148), .b(n_31854), .o(n_32219) );
in01f80 g744218 ( .a(n_36236), .o(n_36237) );
na02f80 g767417 ( .a(n_13521), .b(n_13520), .o(n_13522) );
na02f80 g745534 ( .a(n_34374), .b(FE_OCP_RBN1683_n_33491), .o(n_34404) );
na02f80 g739650 ( .a(n_40548), .b(n_40557), .o(n_40577) );
na02f80 g738221 ( .a(n_41944), .b(n_41943), .o(n_41945) );
na02f80 FE_RC_2384_0 ( .a(FE_RN_925_0), .b(FE_RN_931_0), .o(n_12753) );
ao12f80 g738350 ( .a(n_41595), .b(n_41474), .c(FE_OCP_RBN2312_n_41420), .o(n_41646) );
no02f80 g753260 ( .a(n_27167), .b(FE_OCP_RBN2814_n_25817), .o(n_27213) );
no02f80 g767284 ( .a(n_13608), .b(n_13569), .o(n_13610) );
in01f80 g780220 ( .a(n_45819), .o(n_997) );
na02f80 g755061 ( .a(n_25618), .b(FE_OCP_RBN2421_n_24505), .o(n_25619) );
no02f80 g755259 ( .a(n_24975), .b(n_24840), .o(n_24992) );
ao22s80 g757530 ( .a(n_23261), .b(n_22726), .c(n_23260), .d(n_22727), .o(n_23897) );
no02f80 g771934 ( .a(n_8747), .b(n_7537), .o(n_8748) );
na02f80 g744043 ( .a(n_44221), .b(n_34676), .o(n_35699) );
na02f80 g737316 ( .a(n_42851), .b(n_42757), .o(n_42885) );
in01f80 FE_RC_1190_0 ( .a(n_13693), .o(FE_RN_361_0) );
oa22f80 g751819 ( .a(n_28838), .b(n_179), .c(n_28839), .d(n_186), .o(n_28928) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_4_ ( .ck(newNet_1954), .d(n_10085), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_4_) );
in01f80 newInst_1523 ( .a(newNet_1522), .o(newNet_1523) );
oa22f80 g777901 ( .a(n_47020), .b(FE_OCP_RBN2345_FE_OCPN870_n_2737), .c(n_2741), .d(n_3231), .o(n_3259) );
in01f80 FE_OCP_RBC1341_n_19077 ( .a(n_19077), .o(FE_OCP_RBN1341_n_19077) );
oa12f80 g769391 ( .a(n_11707), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_16_), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_15_), .o(n_11976) );
in01f80 newInst_2877 ( .a(newNet_1862), .o(newNet_2877) );
in01f80 newInst_160 ( .a(newNet_159), .o(newNet_160) );
no02f80 g746835 ( .a(n_33181), .b(n_33058), .o(n_33535) );
no02f80 g759133 ( .a(n_21312), .b(n_21339), .o(n_21419) );
in01f80 newInst_2653 ( .a(newNet_2025), .o(newNet_2653) );
na02f80 g766221 ( .a(n_13141), .b(n_14283), .o(n_14379) );
in01f80 g752969 ( .a(n_28256), .o(n_28257) );
in01f80 g775056 ( .a(n_6054), .o(n_6055) );
na02f80 g750295 ( .a(n_29750), .b(n_29523), .o(n_29779) );
no02f80 g746627 ( .a(n_34666), .b(n_34474), .o(n_34911) );
in01f80 g740649 ( .a(n_39559), .o(n_39558) );
in01f80 g780457 ( .a(n_834), .o(n_883) );
in01f80 g751198 ( .a(n_29884), .o(n_29836) );
in01f80 g753769 ( .a(n_27108), .o(n_27109) );
in01f80 FE_RC_2179_0 ( .a(n_26797), .o(FE_RN_778_0) );
in01f80 newInst_3369 ( .a(newNet_162), .o(newNet_3369) );
in01f80 g736298 ( .a(n_43880), .o(n_43881) );
na02f80 g770092 ( .a(n_10983), .b(n_10982), .o(n_11015) );
no02f80 g775871 ( .a(n_5184), .b(n_5149), .o(n_5185) );
na02f80 g736940 ( .a(n_43038), .b(n_42829), .o(n_43226) );
in01f80 newInst_2448 ( .a(newNet_1861), .o(newNet_2448) );
in01f80 fopt784717 ( .a(n_5524), .o(n_47197) );
ao12f80 g767727 ( .a(n_13082), .b(n_12929), .c(delay_add_ln22_unr8_stage4_stallmux_q_31_), .o(n_13206) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_14_ ( .ck(newNet_187), .d(n_46361), .o(delay_xor_ln22_unr9_stage4_stallmux_q_14_) );
na02f80 g741575 ( .a(n_38643), .b(n_38652), .o(n_38653) );
no02f80 g764736 ( .a(n_15699), .b(n_14419), .o(n_15767) );
in01f80 g775664 ( .a(n_5661), .o(n_5662) );
in01f80 g740192 ( .a(n_39814), .o(n_39815) );
oa22f80 g739401 ( .a(FE_OCPN898_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_9_), .c(n_44775), .d(n_40460), .o(n_41111) );
in01f80 g778995 ( .a(n_2394), .o(n_2863) );
na02f80 g774771 ( .a(n_6241), .b(n_6299), .o(n_6347) );
in01f80 newInst_1418 ( .a(newNet_1417), .o(newNet_1418) );
in01f80 g752819 ( .a(n_27357), .o(n_27437) );
no02f80 g750570 ( .a(n_29446), .b(n_29424), .o(n_29518) );
oa22f80 g751294 ( .a(n_28747), .b(n_28487), .c(n_28707), .d(n_28486), .o(n_28775) );
ao22s80 FE_RC_3431_0 ( .a(FE_OCP_RBN2881_n_21272), .b(n_21464), .c(n_21272), .d(n_21420), .o(n_21640) );
no02f80 g771520 ( .a(n_8878), .b(n_8846), .o(n_8847) );
in01f80 newInst_3223 ( .a(newNet_2227), .o(newNet_3223) );
na02f80 g748845 ( .a(n_31241), .b(n_31032), .o(n_31232) );
oa12f80 g759250 ( .a(n_21114), .b(n_21263), .c(n_21174), .o(n_21415) );
na02f80 g771134 ( .a(n_9635), .b(n_9557), .o(n_9706) );
no02f80 g745935 ( .a(n_33983), .b(n_46955), .o(n_34014) );
no02f80 g745808 ( .a(n_44100), .b(n_34098), .o(n_34128) );
in01f80 FE_OCP_RBC2248_n_13017 ( .a(FE_OCP_RBN2246_n_13017), .o(FE_OCP_RBN2248_n_13017) );
oa12f80 g771632 ( .a(n_9206), .b(n_9482), .c(n_9322), .o(n_9595) );
no02f80 g746787 ( .a(n_33033), .b(n_33056), .o(n_33106) );
na02f80 g750981 ( .a(n_30100), .b(n_30099), .o(n_30101) );
no02f80 g778582 ( .a(n_2421), .b(n_1174), .o(n_2521) );
in01f80 g754484 ( .a(n_25631), .o(n_25675) );
in01f80 g768030 ( .a(n_12885), .o(n_12886) );
na02f80 g739990 ( .a(n_40148), .b(n_40072), .o(n_40195) );
na02f80 g740046 ( .a(n_40292), .b(n_40219), .o(n_40330) );
oa22f80 FE_RC_787_0 ( .a(FE_OFN803_n_46285), .b(n_12240), .c(FE_OFN771_n_46337), .d(n_12189), .o(n_46340) );
in01f80 g759735 ( .a(n_20349), .o(n_20350) );
in01f80 g772962 ( .a(n_7865), .o(n_7866) );
in01f80 newInst_2229 ( .a(newNet_2228), .o(newNet_2229) );
na02f80 g737676 ( .a(FE_OCPN887_n_42367), .b(n_42115), .o(n_42754) );
ao22s80 g736448 ( .a(n_43720), .b(n_43221), .c(n_43719), .d(n_43220), .o(n_43758) );
oa22f80 g780021 ( .a(n_1253), .b(n_988), .c(n_1254), .d(n_987), .o(n_1261) );
na02f80 FE_RC_3138_0 ( .a(FE_RN_1391_0), .b(n_16814), .o(FE_RN_1392_0) );
na02f80 g761073 ( .a(n_19641), .b(n_17900), .o(n_19119) );
in01f80 FE_RC_3829_0 ( .a(n_23229), .o(FE_RN_1669_0) );
oa12f80 g784645 ( .a(n_16787), .b(n_16755), .c(n_16728), .o(n_46975) );
in01f80 g775697 ( .a(n_5478), .o(n_5479) );
na02f80 g742845 ( .a(n_37212), .b(n_37211), .o(n_37213) );
in01f80 g741756 ( .a(n_38506), .o(n_38460) );
na02f80 FE_RC_2754_0 ( .a(n_2624), .b(n_2778), .o(FE_RN_1171_0) );
in01f80 FE_OCP_RBC3631_n_20504 ( .a(n_20504), .o(FE_OCP_RBN3631_n_20504) );
no02f80 g745854 ( .a(n_34068), .b(n_34095), .o(n_34153) );
ao12f80 g757504 ( .a(n_23322), .b(n_44066), .c(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .o(n_23029) );
in01f80 newInst_3082 ( .a(newNet_3081), .o(newNet_3082) );
in01f80 g738665 ( .a(n_41381), .o(n_41393) );
no02f80 g765009 ( .a(n_15464), .b(n_15421), .o(n_15499) );
na02f80 g744458 ( .a(n_35445), .b(n_35340), .o(n_35472) );
in01f80 g751958 ( .a(n_29071), .o(n_29040) );
ao12f80 g751778 ( .a(n_28233), .b(n_28232), .c(n_28234), .o(n_29439) );
no02f80 g765141 ( .a(n_16020), .b(n_15634), .o(n_15975) );
no02f80 g742188 ( .a(FE_OCP_RBN2241_n_44881), .b(n_37875), .o(n_38231) );
no02f80 g774861 ( .a(n_6177), .b(n_5320), .o(n_6244) );
in01f80 FE_RC_3944_0 ( .a(FE_RN_1706_0), .o(FE_OCPN1037_n_28318) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_15_ ( .ck(newNet_2674), .d(n_22359), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_) );
no02f80 g758290 ( .a(n_22187), .b(n_20978), .o(n_22213) );
na02f80 g766070 ( .a(FE_RN_1088_0), .b(n_14587), .o(n_14642) );
in01f80 g742615 ( .a(n_38298), .o(n_37490) );
oa22f80 g738099 ( .a(n_42071), .b(n_41703), .c(n_42037), .d(n_41704), .o(n_42103) );
oa12f80 g773718 ( .a(n_6667), .b(n_7264), .c(n_6741), .o(n_7281) );
na02f80 g774565 ( .a(FE_OCP_RBN1989_delay_xor_ln23_unr6_stage3_stallmux_q), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6524) );
no02f80 g743999 ( .a(n_36036), .b(n_36068), .o(n_36194) );
in01f80 g761248 ( .a(n_19912), .o(n_19766) );
in01f80 newInst_565 ( .a(newNet_163), .o(newNet_565) );
no02f80 g747516 ( .a(n_33705), .b(n_33654), .o(n_33721) );
in01f80 g767329 ( .a(n_13429), .o(n_13487) );
in01f80 g740345 ( .a(n_40271), .o(n_40272) );
in01f80 FE_OCP_RBC2615_n_35005 ( .a(n_35005), .o(FE_OCP_RBN2615_n_35005) );
no02f80 g745529 ( .a(n_34324), .b(n_34323), .o(n_34325) );
oa12f80 g737401 ( .a(n_42700), .b(n_42738), .c(n_42660), .o(n_42778) );
oa22f80 g779886 ( .a(FE_OCPN874_n_44672), .b(n_1137), .c(n_44623), .d(n_1121), .o(n_1306) );
na02f80 g773080 ( .a(n_7716), .b(n_7715), .o(n_7717) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_2_ ( .ck(newNet_498), .d(n_22581), .o(delay_xor_ln22_unr15_stage6_stallmux_q_2_) );
in01f80 drc2 ( .a(n_45808), .o(n_45809) );
oa12f80 g762599 ( .a(n_18042), .b(n_18070), .c(n_18041), .o(n_19665) );
in01f80 g745951 ( .a(n_34078), .o(n_34083) );
in01f80 g745298 ( .a(n_36052), .o(n_36053) );
na02f80 g740422 ( .a(FE_OCP_RBN3026_n_39942), .b(n_39576), .o(n_40205) );
no02f80 g753431 ( .a(n_27019), .b(n_27018), .o(n_27073) );
in01f80 g743798 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_36014) );
na02f80 g767013 ( .a(FE_OCP_RBN3529_n_13765), .b(n_13936), .o(n_14078) );
na02f80 g749658 ( .a(n_30121), .b(n_30013), .o(n_30179) );
na02f80 g772028 ( .a(n_8782), .b(n_8091), .o(n_8860) );
in01f80 g759768 ( .a(n_20677), .o(n_20960) );
no02f80 g763264 ( .a(n_16975), .b(n_17041), .o(n_17195) );
in01f80 newInst_117 ( .a(newNet_18), .o(newNet_117) );
no02f80 FE_RC_3986_0 ( .a(n_14515), .b(FE_RN_1727_0), .o(FE_RN_1728_0) );
no02f80 g755520 ( .a(n_24685), .b(n_24722), .o(n_24874) );
in01f80 g769636 ( .a(n_11275), .o(n_11279) );
no03m80 FE_RC_4046_0 ( .a(n_21351), .b(n_21319), .c(n_21540), .o(n_21638) );
in01f80 fopt784723 ( .a(n_32279), .o(n_47205) );
na02f80 g743380 ( .a(n_36612), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36692) );
ms00f80 delay_add_ln22_unr23_stage9_stallmux_q_reg_2_ ( .ck(newNet_3203), .d(n_35464), .o(delay_add_ln22_unr23_stage9_stallmux_q_2_) );
na02f80 g760493 ( .a(n_19977), .b(n_19773), .o(n_20028) );
na02f80 g770420 ( .a(n_10579), .b(FE_OCP_RBN3604_n_8981), .o(n_10608) );
in01f80 g751376 ( .a(n_28611), .o(n_28551) );
in01f80 g767587 ( .a(n_12875), .o(n_12983) );
in01f80 g770082 ( .a(n_10855), .o(n_10856) );
in01f80 newInst_2494 ( .a(newNet_2493), .o(newNet_2494) );
oa12f80 g747200 ( .a(n_33799), .b(n_33798), .c(n_33797), .o(n_34614) );
oa22f80 FE_RC_391_0 ( .a(n_1129), .b(n_44652), .c(n_1087), .d(n_44637), .o(n_1287) );
in01f80 newInst_1328 ( .a(newNet_1327), .o(newNet_1328) );
na02f80 g775998 ( .a(n_4898), .b(n_4937), .o(n_5085) );
no02f80 g744735 ( .a(n_35175), .b(n_35227), .o(n_35228) );
na02f80 g748229 ( .a(FE_OCP_RBN3731_n_31819), .b(n_30572), .o(n_32138) );
in01f80 g760643 ( .a(n_19778), .o(n_19779) );
no02f80 FE_RC_2620_0 ( .a(FE_RN_1090_0), .b(FE_RN_1091_0), .o(FE_RN_1092_0) );
na02f80 g751947 ( .a(n_28183), .b(n_28182), .o(n_28232) );
ao12f80 g755843 ( .a(n_24391), .b(n_24390), .c(n_24389), .o(n_26125) );
in01f80 newInst_2742 ( .a(newNet_335), .o(newNet_2742) );
in01f80 g738718 ( .a(n_41460), .o(n_41461) );
in01f80 FE_RC_651_0 ( .a(n_6937), .o(FE_RN_208_0) );
oa22f80 FE_RC_1590_0 ( .a(n_2776), .b(n_3274), .c(n_2664), .d(n_2829), .o(n_2930) );
no02f80 FE_RC_1556_0 ( .a(FE_RN_440_0), .b(n_8478), .o(n_8578) );
oa22f80 FE_RC_20_0 ( .a(FE_OFN84_n_46137), .b(n_6567), .c(FE_OFN806_n_46196), .d(FE_OCP_RBN3135_n_6567), .o(n_46186) );
oa22f80 FE_RC_337_0 ( .a(n_22385), .b(n_22682), .c(n_22386), .d(n_47207), .o(n_22835) );
na02f80 g780719 ( .a(n_617), .b(n_468), .o(n_626) );
na02f80 g768469 ( .a(n_12318), .b(FE_OCPN1002_n_45660), .o(n_12431) );
in01f80 newInst_2124 ( .a(newNet_2123), .o(newNet_2124) );
no02f80 g758715 ( .a(FE_OCP_RBN1705_n_21658), .b(n_21711), .o(n_21712) );
na02f80 g778370 ( .a(n_2782), .b(delay_add_ln22_unr2_stage2_stallmux_q_27_), .o(n_2874) );
in01f80 g771897 ( .a(n_9157), .o(n_9124) );
oa22f80 g780859 ( .a(n_420), .b(beta_1), .c(n_580), .d(n_353), .o(n_597) );
na02f80 g777932 ( .a(n_3144), .b(n_2913), .o(n_3145) );
in01f80 g777081 ( .a(n_3743), .o(n_3799) );
na02f80 g771126 ( .a(n_9757), .b(n_9618), .o(n_9795) );
in01f80 FE_OCP_RBC3648_n_15281 ( .a(n_15281), .o(FE_OCP_RBN3648_n_15281) );
no02f80 g764443 ( .a(n_16220), .b(n_14730), .o(n_16273) );
no02f80 g767796 ( .a(n_12929), .b(delay_add_ln22_unr8_stage4_stallmux_q_28_), .o(n_12968) );
in01f80 newInst_1359 ( .a(newNet_1358), .o(newNet_1359) );
ao12f80 g757919 ( .a(n_21960), .b(n_22132), .c(n_21961), .o(n_22204) );
in01f80 fopt784327 ( .a(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(n_46107) );
na02f80 g754982 ( .a(n_25555), .b(n_25500), .o(n_25750) );
in01f80 newInst_2517 ( .a(newNet_1050), .o(newNet_2517) );
no02f80 g737388 ( .a(n_42782), .b(n_42443), .o(n_42784) );
in01f80 FE_OCP_RBC2854_n_45462 ( .a(n_45462), .o(FE_OCP_RBN2854_n_45462) );
no02f80 g768747 ( .a(FE_OCPN867_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_14_), .o(n_12136) );
ao12f80 g766693 ( .a(n_13976), .b(n_14139), .c(n_13876), .o(n_14261) );
in01f80 newInst_2970 ( .a(newNet_2969), .o(newNet_2970) );
ao22s80 FE_RC_3911_0 ( .a(n_22038), .b(n_21988), .c(n_22039), .d(n_21987), .o(n_22068) );
na02f80 g750391 ( .a(n_29591), .b(n_29613), .o(n_29647) );
in01f80 newInst_847 ( .a(newNet_755), .o(newNet_847) );
no02f80 g736805 ( .a(n_43464), .b(n_43387), .o(n_43516) );
na02f80 g766171 ( .a(n_14836), .b(n_14835), .o(n_14837) );
na02f80 g770458 ( .a(n_10513), .b(n_44490), .o(n_10677) );
in01f80 FE_OCP_RBC1848_n_22068 ( .a(FE_OCP_RBN1846_n_22068), .o(FE_OCP_RBN1848_n_22068) );
oa12f80 g781081 ( .a(n_163), .b(n_258), .c(n_159), .o(n_262) );
no02f80 g740590 ( .a(n_45188), .b(n_39642), .o(n_39671) );
in01f80 newInst_0 ( .a(tau_clk), .o(newNet_0) );
na02f80 g771390 ( .a(n_9643), .b(FE_OCPN1402_n_9642), .o(n_9698) );
in01f80 newInst_1774 ( .a(newNet_961), .o(newNet_1774) );
in01f80 FE_RC_500_0 ( .a(n_23266), .o(FE_RN_151_0) );
in01f80 FE_RC_630_0 ( .a(n_17796), .o(FE_RN_195_0) );
na02f80 g754459 ( .a(n_26773), .b(n_26639), .o(n_26815) );
na02f80 FE_RC_3133_0 ( .a(FE_RN_1388_0), .b(FE_OCP_RBN3856_FE_RN_779_0), .o(n_22388) );
in01f80 g772813 ( .a(n_8123), .o(n_8145) );
no02f80 FE_RC_3230_0 ( .a(FE_RN_1131_0), .b(FE_RN_1432_0), .o(n_8902) );
ao22s80 FE_RC_1406_0 ( .a(n_3690), .b(n_3686), .c(FE_OCP_RBN2581_n_3734), .d(n_3687), .o(n_3945) );
in01f80 g748656 ( .a(n_31330), .o(n_31331) );
in01f80 FE_RC_855_0 ( .a(FE_OCPN912_n_43022), .o(FE_RN_255_0) );
no02f80 g764510 ( .a(n_16077), .b(n_16076), .o(n_16218) );
na02f80 g773536 ( .a(n_7412), .b(n_7444), .o(n_7452) );
in01f80 newInst_481 ( .a(newNet_480), .o(newNet_481) );
na02f80 g748666 ( .a(n_31381), .b(n_31398), .o(n_31488) );
oa12f80 g761162 ( .a(n_17783), .b(n_19006), .c(n_18987), .o(n_19153) );
no02f80 g738319 ( .a(n_41861), .b(n_41756), .o(n_41908) );
in01f80 FE_RC_4175_0 ( .a(n_33326), .o(FE_RN_1822_0) );
in01f80 newInst_2371 ( .a(newNet_2090), .o(newNet_2371) );
no02f80 g743921 ( .a(n_35649), .b(n_44223), .o(n_35706) );
no02f80 g760739 ( .a(n_20155), .b(n_20136), .o(n_20182) );
no02f80 g780618 ( .a(n_679), .b(n_693), .o(n_730) );
in01f80 newInst_180 ( .a(newNet_179), .o(newNet_180) );
oa12f80 g780709 ( .a(n_629), .b(n_628), .c(n_627), .o(n_828) );
in01f80 g778608 ( .a(n_2877), .o(n_2842) );
no02f80 g778201 ( .a(n_2871), .b(n_2870), .o(n_2808) );
in01f80 g769736 ( .a(n_11269), .o(n_11289) );
na02f80 g747473 ( .a(n_32387), .b(n_44962), .o(n_32582) );
in01f80 g748325 ( .a(n_31838), .o(n_31839) );
no02f80 g777734 ( .a(n_3425), .b(n_3406), .o(n_3431) );
in01f80 FE_RC_2935_0 ( .a(FE_RN_1280_0), .o(n_15036) );
in01f80 g758959 ( .a(n_22331), .o(n_21393) );
na02f80 g764580 ( .a(n_16506), .b(n_16505), .o(n_16507) );
na02f80 g766132 ( .a(n_14507), .b(FE_OCP_RBN3430_n_13245), .o(n_14579) );
ao12f80 g784673 ( .a(n_5161), .b(n_5123), .c(n_4723), .o(n_47003) );
no02f80 g737447 ( .a(n_42655), .b(n_42372), .o(n_42722) );
in01f80 FE_RC_179_0 ( .a(n_12296), .o(FE_RN_58_0) );
in01f80 newInst_1617 ( .a(newNet_1616), .o(newNet_1617) );
no02f80 g771470 ( .a(n_9046), .b(n_8936), .o(n_9116) );
in01f80 g753702 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_1_), .o(n_27865) );
oa22f80 FE_RC_4134_0 ( .a(FE_RN_733_0), .b(FE_RN_734_0), .c(FE_RN_735_0), .d(n_24270), .o(n_24446) );
in01f80 newInst_763 ( .a(newNet_762), .o(newNet_763) );
in01f80 g756450 ( .a(n_23771), .o(n_23772) );
ao12f80 g778219 ( .a(n_2748), .b(n_2763), .c(n_2828), .o(n_2859) );
oa12f80 g752397 ( .a(n_28256), .b(n_28401), .c(n_28297), .o(n_28435) );
in01f80 FE_OCP_RBC2047_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2047_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01f80 g759305 ( .a(n_21044), .o(n_21045) );
no02f80 g775332 ( .a(n_5586), .b(n_5654), .o(n_5655) );
in01f80 FE_OCP_RBC3084_n_31819 ( .a(n_31819), .o(FE_OCP_RBN3084_n_31819) );
na02f80 g745713 ( .a(n_34284), .b(n_34338), .o(n_34367) );
no02f80 g762085 ( .a(n_18242), .b(n_17416), .o(n_18280) );
in01f80 g763055 ( .a(n_17683), .o(n_17509) );
no02f80 g759684 ( .a(n_20508), .b(n_20480), .o(n_20597) );
oa12f80 g756531 ( .a(n_23520), .b(n_23545), .c(n_23519), .o(n_24962) );
in01f80 g758136 ( .a(n_23201), .o(n_23202) );
ao12f80 g742930 ( .a(n_37005), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_25_), .o(n_37065) );
ao22s80 g779221 ( .a(n_1761), .b(n_1838), .c(n_1760), .d(n_1811), .o(n_1880) );
in01f80 FE_OCP_RBC2410_n_13960 ( .a(n_13960), .o(FE_OCP_RBN2410_n_13960) );
in01f80 g754182 ( .a(n_25999), .o(n_25998) );
no02f80 g760613 ( .a(n_19814), .b(n_18140), .o(n_19815) );
na02f80 FE_RC_3505_0 ( .a(FE_RN_1513_0), .b(n_29030), .o(FE_RN_1514_0) );
in01f80 newInst_1156 ( .a(newNet_1155), .o(newNet_1156) );
na02f80 g770581 ( .a(n_10106), .b(n_10105), .o(n_10153) );
na02f80 FE_RC_3725_0 ( .a(FE_RN_1637_0), .b(FE_RN_1638_0), .o(FE_RN_1639_0) );
no02f80 g755534 ( .a(FE_OCP_RBN2402_n_24638), .b(FE_OFN785_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24722) );
no02f80 FE_RC_2199_0 ( .a(FE_OCPN1508_n_23414), .b(FE_RN_789_0), .o(FE_RN_790_0) );
no02f80 g767812 ( .a(n_13119), .b(n_13017), .o(n_13378) );
in01f80 newInst_1751 ( .a(newNet_1750), .o(newNet_1751) );
ao12f80 g754530 ( .a(n_25431), .b(n_25432), .c(n_25241), .o(n_25518) );
in01f80 g740238 ( .a(n_39971), .o(n_39972) );
na02f80 g757244 ( .a(n_23189), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_), .o(n_23190) );
in01f80 g753479 ( .a(n_26879), .o(n_26880) );
na02f80 g738474 ( .a(n_41660), .b(n_41320), .o(n_41808) );
na02f80 g752042 ( .a(n_28181), .b(n_28140), .o(n_28224) );
ao22s80 g759827 ( .a(n_21691), .b(n_21835), .c(n_21714), .d(n_20255), .o(n_21890) );
in01f80 g740997 ( .a(n_39084), .o(n_39085) );
in01f80 FE_OCP_RBC2901_n_44174 ( .a(n_44174), .o(FE_OCP_RBN2901_n_44174) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_0_ ( .ck(newNet_1437), .d(FE_OFN221_n_35655), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_0_) );
no02f80 g779597 ( .a(n_1800), .b(delay_xor_ln22_unr3_stage2_stallmux_q_24_), .o(n_2011) );
no02f80 g763275 ( .a(FE_OCP_RBN3213_n_44365), .b(delay_xor_ln21_unr12_stage5_stallmux_q_4_), .o(n_17197) );
na02f80 g750888 ( .a(n_29018), .b(n_29017), .o(n_29019) );
no02f80 g753256 ( .a(n_27377), .b(n_25873), .o(n_27464) );
in01f80 g745380 ( .a(n_35882), .o(n_35961) );
ao12f80 g757364 ( .a(n_23307), .b(n_44066), .c(delay_xor_ln22_unr15_stage6_stallmux_q_9_), .o(n_23017) );
no02f80 g751828 ( .a(n_28228), .b(n_28227), .o(n_28252) );
in01f80 g737588 ( .a(n_42683), .o(n_42684) );
no02f80 g740457 ( .a(n_39712), .b(n_39703), .o(n_39739) );
no02f80 g772799 ( .a(n_8123), .b(n_8121), .o(n_8245) );
na02f80 g743826 ( .a(n_37168), .b(n_46202), .o(n_37217) );
in01f80 FE_RC_4010_0 ( .a(FE_OCPN1773_n_30210), .o(FE_RN_1741_0) );
in01f80 fopt782746 ( .a(FE_OCP_RBN1911_n_20545), .o(n_44160) );
na02f80 g776021 ( .a(n_4872), .b(n_4878), .o(n_4898) );
oa22f80 FE_RC_3392_0 ( .a(n_38109), .b(n_38449), .c(n_38108), .d(n_38448), .o(n_38530) );
na02f80 g755359 ( .a(n_24914), .b(n_24961), .o(n_25020) );
in01f80 g760842 ( .a(n_19516), .o(n_19566) );
in01f80 newInst_1649 ( .a(newNet_1455), .o(newNet_1649) );
na02f80 g761489 ( .a(n_19647), .b(n_19735), .o(n_19849) );
oa12f80 g759320 ( .a(n_20917), .b(n_20956), .c(n_21041), .o(n_21074) );
no02f80 g737791 ( .a(n_42205), .b(n_42204), .o(n_42206) );
in01f80 g736615 ( .a(n_43376), .o(n_43377) );
in01f80 g773286 ( .a(n_7612), .o(n_7599) );
in01f80 FE_OCP_RBC3495_n_19390 ( .a(FE_OCP_RBN3494_n_19390), .o(FE_OCP_RBN3495_n_19390) );
no02f80 g781330 ( .a(n_7), .b(beta_21), .o(n_69) );
ao22s80 FE_RC_898_0 ( .a(n_30534), .b(n_27062), .c(FE_OCPN1410_n_27014), .d(FE_OCP_RBN2805_n_30534), .o(n_30625) );
in01f80 FE_OCP_RBC2858_n_10399 ( .a(n_10399), .o(FE_OCP_RBN2858_n_10399) );
in01f80 fopt783258 ( .a(n_44827), .o(n_44826) );
in01f80 g748158 ( .a(n_32099), .o(n_32100) );
na02f80 g777882 ( .a(n_3174), .b(n_45190), .o(n_3239) );
no02f80 g774230 ( .a(n_6578), .b(n_6552), .o(n_6665) );
na02f80 g776965 ( .a(n_3790), .b(n_3837), .o(n_3955) );
in01f80 g765104 ( .a(n_16310), .o(n_16311) );
no02f80 g741266 ( .a(FE_OCPN942_n_44925), .b(n_38473), .o(n_39318) );
in01f80 FE_OCP_RBC1349_n_19270 ( .a(FE_OCP_RBN1348_n_19270), .o(FE_OCP_RBN1349_n_19270) );
in01f80 g743930 ( .a(n_36039), .o(n_36040) );
in01f80 g762741 ( .a(n_17917), .o(n_17891) );
na02f80 g751611 ( .a(n_29252), .b(n_29251), .o(n_29253) );
in01f80 newInst_1994 ( .a(newNet_1993), .o(newNet_1994) );
ms00f80 delay_sub_ln21_unr24_stage9_stallmux_q_reg_2_ ( .ck(newNet_1935), .d(n_36776), .o(delay_sub_ln21_unr24_stage9_stallmux_q_2_) );
na02f80 g753429 ( .a(n_27019), .b(n_27018), .o(n_27068) );
no02f80 g768639 ( .a(n_12072), .b(n_12193), .o(n_12265) );
no02f80 g743094 ( .a(n_36537), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37110) );
na02f80 g758805 ( .a(n_22209), .b(n_22179), .o(n_22180) );
in01f80 g773484 ( .a(n_46992), .o(n_7518) );
na02f80 g742456 ( .a(n_37607), .b(n_37583), .o(n_37697) );
in01f80 g758396 ( .a(n_23590), .o(n_23564) );
no02f80 g761329 ( .a(n_19761), .b(n_19711), .o(n_20087) );
no02f80 FE_RC_2734_0 ( .a(FE_RN_1158_0), .b(n_22958), .o(n_46964) );
in01f80 g758772 ( .a(n_21734), .o(n_21735) );
ao12f80 g778184 ( .a(n_2774), .b(n_3006), .c(FE_OCP_RBN2290_n_2438), .o(n_2865) );
oa12f80 g759376 ( .a(n_20714), .b(n_20933), .c(n_20676), .o(n_21067) );
in01f80 FE_OCP_RBC3581_n_44944 ( .a(FE_OCP_RBN2545_n_44944), .o(FE_OCP_RBN3581_n_44944) );
oa22f80 g743636 ( .a(n_36349), .b(n_35779), .c(n_36350), .d(n_35778), .o(n_36414) );
oa22f80 FE_RC_1458_0 ( .a(n_17336), .b(n_17834), .c(n_17753), .d(n_17803), .o(n_17878) );
in01f80 newInst_95 ( .a(newNet_94), .o(newNet_95) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_19_ ( .ck(newNet_3058), .d(n_1065), .o(delay_add_ln22_unr2_stage2_stallmux_q_19_) );
in01f80 g761586 ( .a(n_20252), .o(n_22801) );
in01f80 FE_OCP_DRV_C1547_n_17643 ( .a(n_17643), .o(FE_OCP_DRV_N1547_n_17643) );
in01f80 newInst_1668 ( .a(newNet_1667), .o(newNet_1668) );
no02f80 g770730 ( .a(n_10142), .b(n_9965), .o(n_10236) );
in01f80 FE_OCP_RBC3271_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3271_n_45224) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_19_ ( .ck(newNet_2001), .d(n_11494), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_19_) );
ao22s80 g762718 ( .a(n_18210), .b(n_17356), .c(n_18157), .d(n_17357), .o(n_18529) );
na02f80 g742225 ( .a(n_44875), .b(n_38270), .o(n_37995) );
no02f80 g763368 ( .a(n_16836), .b(FE_OCP_RBN3659_n_15314), .o(n_16952) );
na02f80 g770530 ( .a(n_10362), .b(n_10397), .o(n_10513) );
no02f80 g737600 ( .a(n_42444), .b(n_42443), .o(n_42465) );
ao12f80 g772307 ( .a(n_8726), .b(n_8725), .c(n_8724), .o(n_9768) );
na02f80 g764903 ( .a(n_15473), .b(n_15502), .o(n_15622) );
in01f80 g752712 ( .a(n_27358), .o(n_27359) );
no02f80 FE_RC_1555_0 ( .a(FE_RN_438_0), .b(FE_RN_439_0), .o(FE_RN_440_0) );
no02f80 g749377 ( .a(n_30604), .b(n_30296), .o(n_30670) );
in01f80 g752319 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_30_), .o(n_27833) );
in01f80 newInst_3076 ( .a(newNet_1515), .o(newNet_3076) );
no02f80 g771452 ( .a(FE_OCP_RBN3583_n_9245), .b(n_9132), .o(n_9340) );
no02f80 g776736 ( .a(n_4257), .b(n_4179), .o(n_4436) );
na02f80 g740719 ( .a(n_39387), .b(n_39189), .o(n_39449) );
in01f80 g750091 ( .a(n_29864), .o(n_29865) );
in01f80 g779794 ( .a(n_1484), .o(n_1645) );
ao12f80 g748098 ( .a(n_32839), .b(n_32838), .c(n_32837), .o(n_32900) );
in01f80 g770181 ( .a(n_10757), .o(n_10758) );
no02f80 g750116 ( .a(FE_OCP_RBN2573_n_29922), .b(n_30191), .o(n_30278) );
in01f80 g740027 ( .a(n_39955), .o(n_39956) );
oa12f80 g746299 ( .a(n_33639), .b(n_33638), .c(n_33637), .o(n_34200) );
oa12f80 g736580 ( .a(n_301), .b(n_43655), .c(FE_OFN2_n_43918), .o(n_43693) );
oa22f80 g744528 ( .a(n_36678), .b(n_36250), .c(n_36662), .d(n_36251), .o(n_36726) );
ao12f80 g755158 ( .a(n_25021), .b(n_25020), .c(n_25049), .o(n_25100) );
na02f80 g741970 ( .a(n_38037), .b(n_38089), .o(n_38114) );
na02f80 g745325 ( .a(n_35716), .b(n_35717), .o(n_35886) );
in01f80 g765295 ( .a(n_15964), .o(n_15965) );
in01f80 g776092 ( .a(n_4789), .o(n_4790) );
na02f80 g773244 ( .a(n_7709), .b(n_7670), .o(n_7735) );
oa22f80 FE_RC_390_0 ( .a(n_1010), .b(n_44652), .c(n_993), .d(n_44637), .o(n_1301) );
no02f80 g743070 ( .a(n_37171), .b(n_36928), .o(n_37172) );
ao12f80 g755284 ( .a(n_25639), .b(n_25638), .c(n_25637), .o(n_26451) );
ao12f80 g784441 ( .a(n_37202), .b(n_37169), .c(n_46204), .o(n_46253) );
in01f80 g780074 ( .a(n_1220), .o(n_1218) );
in01f80 g776133 ( .a(n_4624), .o(n_4690) );
na03f80 g743323 ( .a(n_37773), .b(n_37854), .c(n_37789), .o(n_37920) );
in01f80 g760448 ( .a(n_20075), .o(n_20076) );
no02f80 g776839 ( .a(n_3919), .b(n_3851), .o(n_4000) );
no02f80 g769271 ( .a(n_11439), .b(n_11435), .o(n_11458) );
no02f80 g761152 ( .a(n_19131), .b(n_19170), .o(n_19171) );
na02f80 g775345 ( .a(n_5768), .b(n_5785), .o(n_5835) );
na02f80 g766415 ( .a(n_14032), .b(n_14000), .o(n_14034) );
in01f80 g743282 ( .a(n_36761), .o(n_36771) );
na02f80 g755816 ( .a(n_25316), .b(n_25318), .o(n_24316) );
in01f80 FE_RC_1317_0 ( .a(n_43143), .o(FE_RN_388_0) );
oa12f80 g776518 ( .a(n_4334), .b(n_4446), .c(n_4572), .o(n_4619) );
no02f80 g765496 ( .a(n_15664), .b(n_15747), .o(n_15781) );
in01f80 newInst_2673 ( .a(newNet_2672), .o(newNet_2673) );
in01f80 FE_OCPC1510_n_44174 ( .a(FE_OCPN1509_n_44174), .o(FE_OCPN1510_n_44174) );
in01f80 FE_OCP_RBC2507_n_13896 ( .a(FE_OCP_RBN2502_n_13896), .o(FE_OCP_RBN2507_n_13896) );
oa12f80 g749151 ( .a(n_30747), .b(n_30714), .c(n_30584), .o(n_30751) );
oa12f80 g770536 ( .a(n_10462), .b(n_10498), .c(n_10461), .o(n_10524) );
in01f80 newInst_2350 ( .a(newNet_2349), .o(newNet_2350) );
in01f80 g770394 ( .a(n_10636), .o(n_10705) );
no02f80 FE_RC_1220_0 ( .a(FE_RN_368_0), .b(n_33922), .o(n_34427) );
in01f80 g750795 ( .a(n_46960), .o(n_29327) );
ao12f80 g751068 ( .a(n_29881), .b(n_30156), .c(n_29838), .o(n_30339) );
in01f80 g761904 ( .a(n_18321), .o(n_18373) );
in01f80 FE_OCP_RBC1703_n_19560 ( .a(FE_OCP_RBN1702_n_19560), .o(FE_OCP_RBN1703_n_19560) );
no02f80 g778354 ( .a(n_2604), .b(n_2498), .o(n_2647) );
in01f80 g778008 ( .a(n_3218), .o(n_3163) );
no02f80 g760785 ( .a(n_19591), .b(FE_OCP_DRV_N1558_n_19590), .o(n_19692) );
na02f80 g776047 ( .a(n_5107), .b(n_5053), .o(n_5054) );
no02f80 g765862 ( .a(n_14879), .b(n_14855), .o(n_14979) );
na02f80 g780293 ( .a(n_1104), .b(n_1103), .o(n_1105) );
in01f80 g762664 ( .a(n_18000), .o(n_17949) );
na02f80 g742919 ( .a(n_37069), .b(n_36996), .o(n_37118) );
ao12f80 g739025 ( .a(n_41139), .b(n_41138), .c(n_41137), .o(n_41545) );
na02f80 g749354 ( .a(n_30540), .b(n_30790), .o(n_30586) );
na02f80 g758926 ( .a(n_21238), .b(n_45026), .o(n_21292) );
in01f80 g762074 ( .a(n_18354), .o(n_18425) );
no02f80 FE_RC_2648_0 ( .a(n_12176), .b(n_12069), .o(FE_RN_1105_0) );
no02f80 g743372 ( .a(n_37830), .b(n_46232), .o(n_37803) );
no02f80 g746587 ( .a(n_34666), .b(n_34735), .o(n_34809) );
na02f80 g751711 ( .a(n_28403), .b(n_28358), .o(n_28415) );
no02f80 g777826 ( .a(n_3295), .b(n_3276), .o(n_3379) );
na02f80 g772718 ( .a(n_8195), .b(FE_OCP_RBN2329_n_9003), .o(n_8196) );
no02f80 g756815 ( .a(n_23754), .b(n_23812), .o(n_23813) );
na03f80 g783833 ( .a(n_14612), .b(n_14586), .c(FE_OCP_RBN3535_n_13765), .o(n_45519) );
na02f80 g770604 ( .a(FE_OCP_RBN2797_n_10106), .b(n_9204), .o(n_10357) );
in01f80 g767028 ( .a(n_14208), .o(n_14209) );
ao12f80 g778547 ( .a(n_2617), .b(n_2620), .c(n_3029), .o(n_3434) );
na02f80 g738466 ( .a(n_41387), .b(n_41173), .o(n_41472) );
no02f80 g760305 ( .a(n_20228), .b(n_18944), .o(n_20244) );
in01f80 g775379 ( .a(n_5913), .o(n_5906) );
in01f80 g771571 ( .a(n_8974), .o(n_8975) );
no02f80 g747744 ( .a(n_33372), .b(n_33743), .o(n_33991) );
ao22s80 g780337 ( .a(n_1208), .b(n_801), .c(n_1122), .d(n_800), .o(n_897) );
na02f80 g751471 ( .a(FE_OCPN962_n_28506), .b(n_28472), .o(n_28777) );
na02f80 g768889 ( .a(n_44356), .b(n_11604), .o(n_11791) );
in01f80 g778750 ( .a(n_2420), .o(n_2421) );
in01f80 g778239 ( .a(n_2777), .o(n_2856) );
no02f80 g779572 ( .a(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_5_), .o(n_1425) );
no02f80 g783845 ( .a(n_39594), .b(n_39579), .o(n_45531) );
in01f80 g770495 ( .a(n_10330), .o(n_10331) );
in01f80 g779971 ( .a(delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .o(n_1358) );
in01f80 g753118 ( .a(n_27504), .o(n_27505) );
na02f80 g770030 ( .a(n_10833), .b(n_44498), .o(n_10894) );
ao12f80 g780298 ( .a(n_827), .b(n_995), .c(n_1002), .o(n_1056) );
in01f80 g739576 ( .a(n_40645), .o(n_40875) );
no02f80 g758811 ( .a(n_21730), .b(FE_OCP_RBN2953_n_21538), .o(n_21765) );
in01f80 FE_OCP_RBC3053_n_39913 ( .a(n_39913), .o(FE_OCP_RBN3053_n_39913) );
na02f80 g762233 ( .a(n_18135), .b(n_18133), .o(n_18134) );
in01f80 g757374 ( .a(n_24158), .o(n_24283) );
na02f80 g764690 ( .a(n_15704), .b(n_15408), .o(n_15742) );
no02f80 g771875 ( .a(n_9004), .b(n_9003), .o(n_9099) );
ao12f80 g779483 ( .a(n_1664), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln21_unr3_stage2_stallmux_q_12_), .o(n_1717) );
in01f80 g773509 ( .a(n_7676), .o(n_8453) );
na02f80 g777387 ( .a(n_3551), .b(n_3549), .o(n_3643) );
na02f80 g751882 ( .a(n_29043), .b(n_29003), .o(n_29044) );
na02f80 g752147 ( .a(n_28635), .b(n_28202), .o(n_28711) );
in01f80 g772976 ( .a(n_7799), .o(n_7835) );
in01f80 g744009 ( .a(n_36316), .o(n_36317) );
no02f80 g743101 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_), .o(n_37094) );
in01f80 FE_OCP_RBC1730_n_22492 ( .a(n_22492), .o(FE_OCP_RBN1730_n_22492) );
oa12f80 g773392 ( .a(n_7695), .b(n_7608), .c(delay_sub_ln21_0_unr5_stage3_stallmux_q_31_), .o(n_7764) );
no02f80 g741955 ( .a(n_38042), .b(n_37978), .o(n_38090) );
in01f80 g763135 ( .a(n_17882), .o(n_17883) );
oa12f80 g736499 ( .a(n_326), .b(n_43653), .c(FE_OFN3_n_43918), .o(n_43677) );
oa12f80 g750627 ( .a(n_29438), .b(n_29437), .c(n_29436), .o(n_30859) );
in01f80 newInst_1386 ( .a(newNet_1385), .o(newNet_1386) );
no02f80 g769035 ( .a(FE_OCP_RBN2119_n_45224), .b(delay_xor_ln22_unr9_stage4_stallmux_q_8_), .o(n_11840) );
na02f80 g778631 ( .a(n_2402), .b(n_2322), .o(n_2714) );
in01f80 g768789 ( .a(n_12041), .o(n_12042) );
na02f80 g776564 ( .a(n_4287), .b(n_4286), .o(n_4348) );
in01f80 g768771 ( .a(n_12098), .o(n_12099) );
no02f80 g772531 ( .a(n_8569), .b(n_8568), .o(n_8642) );
in01f80 g748341 ( .a(n_31833), .o(n_31834) );
no02f80 g779526 ( .a(n_1570), .b(n_1569), .o(n_1586) );
no02f80 g770617 ( .a(n_10428), .b(n_8687), .o(n_10429) );
na02f80 g759650 ( .a(n_21300), .b(n_21136), .o(n_21881) );
in01f80 newInst_2989 ( .a(newNet_2988), .o(newNet_2989) );
in01f80 g739333 ( .a(n_40732), .o(n_40733) );
ao12f80 g753843 ( .a(n_23414), .b(n_26218), .c(n_26078), .o(n_26366) );
in01f80 g756189 ( .a(n_24145), .o(n_24127) );
no02f80 g741280 ( .a(n_44921), .b(n_38912), .o(n_39000) );
na02f80 g757394 ( .a(n_23040), .b(n_23015), .o(n_23067) );
na02f80 g740401 ( .a(FE_OCP_RBN3027_n_39942), .b(n_39932), .o(n_39964) );
in01f80 newInst_1931 ( .a(newNet_1930), .o(newNet_1931) );
na02f80 g752586 ( .a(n_27571), .b(n_27505), .o(n_27585) );
na02f80 g753770 ( .a(n_27097), .b(n_26741), .o(n_27108) );
oa12f80 g744473 ( .a(n_35457), .b(n_35456), .c(n_35467), .o(n_35481) );
no02f80 g764760 ( .a(n_15596), .b(n_15559), .o(n_15706) );
in01f80 newInst_1239 ( .a(newNet_1238), .o(newNet_1239) );
na02f80 g756273 ( .a(n_24607), .b(n_24107), .o(n_24740) );
in01f80 newInst_2613 ( .a(newNet_116), .o(newNet_2613) );
no02f80 FE_RC_795_0 ( .a(FE_RN_242_0), .b(n_41453), .o(n_41522) );
in01f80 FE_RC_3141_0 ( .a(FE_OCP_RBN1191_n_14911), .o(FE_RN_1394_0) );
in01f80 g743703 ( .a(n_36327), .o(n_36328) );
in01f80 FE_OCP_RBC3580_n_44944 ( .a(FE_OCP_RBN2545_n_44944), .o(FE_OCP_RBN3580_n_44944) );
oa12f80 g757519 ( .a(n_22153), .b(n_22639), .c(n_22128), .o(n_22722) );
na02f80 g762692 ( .a(n_17996), .b(n_17995), .o(n_18066) );
no02f80 g745699 ( .a(n_34180), .b(n_34206), .o(n_34207) );
na02f80 g758669 ( .a(n_22397), .b(n_21780), .o(n_22489) );
oa12f80 g761934 ( .a(n_18268), .b(n_18291), .c(n_17508), .o(n_18477) );
in01f80 g763922 ( .a(n_17096), .o(n_17097) );
in01f80 g776592 ( .a(n_4482), .o(n_4483) );
no02f80 g745286 ( .a(n_36123), .b(n_35805), .o(n_36174) );
in01f80 FE_OCP_DRV_C1579_n_35482 ( .a(n_35482), .o(FE_OCP_DRV_N1579_n_35482) );
in01f80 FE_OCP_RBC2050_delay_sub_ln23_unr17_stage6_stallmux_q_1_ ( .a(FE_OCP_RBN2048_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .o(FE_OCP_RBN2050_delay_sub_ln23_unr17_stage6_stallmux_q_1_) );
in01f80 newInst_3093 ( .a(newNet_3092), .o(newNet_3093) );
ao12f80 g780790 ( .a(n_529), .b(n_528), .c(n_527), .o(n_553) );
in01f80 g776859 ( .a(n_4226), .o(n_4227) );
no02f80 g745633 ( .a(n_34289), .b(FE_OCP_DRV_N1560_n_34288), .o(n_34376) );
oa12f80 g745339 ( .a(n_35927), .b(FE_OCP_RBN2995_n_35539), .c(n_35931), .o(n_36161) );
no02f80 g754689 ( .a(FE_OCP_RBN2955_n_26231), .b(n_26451), .o(n_26486) );
no02f80 g767976 ( .a(n_13035), .b(n_12781), .o(n_13473) );
ao12f80 g746519 ( .a(n_34666), .b(n_34699), .c(n_34733), .o(n_34777) );
ao12f80 g751346 ( .a(n_29079), .b(n_29487), .c(n_29488), .o(n_29537) );
no02f80 g742127 ( .a(n_38254), .b(n_38231), .o(n_38317) );
no02f80 g744088 ( .a(n_35534), .b(n_35575), .o(n_35576) );
no02f80 g776114 ( .a(n_4558), .b(n_4557), .o(n_4559) );
na02f80 g775310 ( .a(FE_OCP_RBN2979_n_5656), .b(n_5614), .o(n_5706) );
ao22s80 FE_RC_46_0 ( .a(FE_OCPN959_n_3951), .b(n_3971), .c(n_5603), .d(n_4182), .o(n_4265) );
in01f80 g776342 ( .a(n_4880), .o(n_4881) );
no02f80 FE_RC_2869_0 ( .a(FE_RN_1239_0), .b(n_24562), .o(FE_RN_1238_0) );
in01f80 g772897 ( .a(n_8001), .o(n_8002) );
na02f80 g743832 ( .a(n_35835), .b(n_35834), .o(n_35836) );
no02f80 g761659 ( .a(n_19486), .b(n_19485), .o(n_19487) );
ao22s80 FE_RC_2147_0 ( .a(FE_RN_752_0), .b(n_15561), .c(n_15588), .d(FE_RN_756_0), .o(n_15700) );
na02f80 g780543 ( .a(n_713), .b(n_46055), .o(n_778) );
no03m80 g767235 ( .a(n_13700), .b(n_13698), .c(n_13271), .o(n_13798) );
in01f80 g754037 ( .a(n_26245), .o(n_26246) );
na02f80 g759513 ( .a(n_20649), .b(n_20555), .o(n_20691) );
na02f80 g770718 ( .a(n_10304), .b(n_10245), .o(n_10415) );
no02f80 g758941 ( .a(n_21572), .b(n_21575), .o(n_21678) );
in01f80 g769779 ( .a(n_11172), .o(n_11173) );
oa12f80 g751032 ( .a(n_29806), .b(n_29805), .c(n_29804), .o(n_29856) );
oa12f80 g761525 ( .a(n_18896), .b(n_18895), .c(n_18894), .o(n_18974) );
in01f80 g763490 ( .a(n_16838), .o(n_16876) );
no02f80 g749531 ( .a(n_31781), .b(n_31509), .o(n_31885) );
na02f80 g777258 ( .a(n_3450), .b(n_3483), .o(n_3484) );
no02f80 g736608 ( .a(n_43646), .b(n_43564), .o(n_43645) );
in01f80 FE_OCP_RBC2162_n_12312 ( .a(n_12312), .o(FE_OCP_RBN2162_n_12312) );
in01f80 g760813 ( .a(n_19476), .o(n_19477) );
in01f80 g777247 ( .a(n_3625), .o(n_3680) );
no02f80 g772592 ( .a(n_8350), .b(n_8325), .o(n_8454) );
na02f80 g748676 ( .a(n_32509), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_3_), .o(n_32562) );
no02f80 g752849 ( .a(n_27428), .b(n_27394), .o(n_27509) );
in01f80 g739426 ( .a(n_40724), .o(n_40858) );
oa22f80 FE_RC_3237_0 ( .a(n_9173), .b(n_9754), .c(n_9111), .d(n_9855), .o(n_9941) );
in01f80 newInst_109 ( .a(newNet_91), .o(newNet_109) );
in01f80 newInst_1888 ( .a(newNet_1887), .o(newNet_1888) );
oa12f80 g736377 ( .a(n_329), .b(n_43794), .c(FE_OFN2_n_43918), .o(n_43852) );
oa12f80 g751806 ( .a(n_28958), .b(n_28903), .c(n_28793), .o(n_28959) );
in01f80 FE_OCP_RBC2404_n_24638 ( .a(FE_OCP_RBN2403_n_24638), .o(FE_OCP_RBN2404_n_24638) );
ao12f80 g738233 ( .a(n_41926), .b(n_41940), .c(n_41925), .o(n_42366) );
no02f80 g768876 ( .a(n_11927), .b(n_11919), .o(n_11909) );
no02f80 g737413 ( .a(n_42719), .b(n_42620), .o(n_42753) );
in01f80 g767046 ( .a(n_14291), .o(n_14292) );
no02f80 g769949 ( .a(n_10996), .b(n_10997), .o(n_11074) );
no02f80 g753878 ( .a(n_26219), .b(n_26198), .o(n_26268) );
na02f80 g772572 ( .a(FE_OCP_RBN2371_n_8221), .b(n_7743), .o(n_8277) );
no02f80 g749878 ( .a(FE_OCP_RBN3010_n_31117), .b(n_30970), .o(n_31411) );
in01f80 g777393 ( .a(n_3576), .o(n_3577) );
ao12f80 g761670 ( .a(n_18776), .b(n_19370), .c(n_18581), .o(n_19542) );
oa22f80 g746875 ( .a(FE_OCP_RBN3390_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_13_), .c(n_33108), .d(n_32083), .o(n_33455) );
no02f80 FE_RC_175_0 ( .a(FE_RN_56_0), .b(FE_RN_55_0), .o(FE_RN_54_0) );
in01f80 g766292 ( .a(n_14441), .o(n_16215) );
oa12f80 g750452 ( .a(n_30550), .b(n_30549), .c(n_30548), .o(n_31223) );
oa22f80 FE_RC_3462_0 ( .a(n_24350), .b(n_27782), .c(n_27845), .d(n_45309), .o(n_27836) );
in01f80 g781220 ( .a(n_162), .o(n_169) );
na02f80 g742519 ( .a(n_37581), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37604) );
in01f80 g739813 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_10_), .o(n_40461) );
na02f80 g760365 ( .a(n_20212), .b(n_20211), .o(n_20213) );
in01f80 FE_OCP_RBC3698_n_35543 ( .a(FE_OCP_RBN3697_n_35543), .o(FE_OCP_RBN3698_n_35543) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_4_ ( .ck(newNet_2151), .d(n_921), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_4_) );
in01f80 g773607 ( .a(n_7414), .o(n_7415) );
no02f80 g769045 ( .a(FE_OCP_RBN3269_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_5_), .o(n_11693) );
no02f80 g784401 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_15_), .o(n_46213) );
in01f80 FE_RC_2108_0 ( .a(n_30937), .o(FE_RN_729_0) );
oa12f80 g776387 ( .a(n_4501), .b(n_4619), .c(n_4382), .o(n_4786) );
oa12f80 g772630 ( .a(n_8274), .b(n_8275), .c(n_8273), .o(n_9988) );
no02f80 g778764 ( .a(n_2354), .b(n_2030), .o(n_2382) );
na02f80 FE_RC_3980_0 ( .a(n_29630), .b(n_29417), .o(FE_RN_1725_0) );
in01f80 g754834 ( .a(n_26679), .o(n_26033) );
na02f80 g770672 ( .a(n_10057), .b(FE_OCP_RBN3597_FE_OCPN1243_n_44460), .o(n_10096) );
in01f80 g758260 ( .a(n_22695), .o(n_22646) );
na02f80 g779227 ( .a(n_1822), .b(n_1047), .o(n_1891) );
no02f80 g770912 ( .a(n_9630), .b(n_9627), .o(n_9855) );
na02f80 g745795 ( .a(n_34124), .b(n_34427), .o(n_34126) );
oa12f80 g736511 ( .a(n_43478), .b(n_43661), .c(n_43223), .o(n_43712) );
na02f80 g753495 ( .a(n_26912), .b(n_26838), .o(n_26954) );
oa22f80 g752979 ( .a(n_27044), .b(n_26915), .c(n_27045), .d(n_26916), .o(n_27090) );
no02f80 g762307 ( .a(n_18093), .b(n_18054), .o(n_18167) );
no02f80 g738034 ( .a(n_42140), .b(n_42123), .o(n_42150) );
in01f80 FE_RC_940_0 ( .a(FE_RN_278_0), .o(n_22625) );
in01f80 g752283 ( .a(n_28001), .o(n_28270) );
na02f80 g780379 ( .a(n_955), .b(n_580), .o(n_915) );
oa22f80 g743444 ( .a(n_36506), .b(n_36094), .c(FE_OCP_RBN3057_n_36506), .d(n_36093), .o(n_36594) );
na02f80 g742982 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_12_), .o(n_37079) );
in01f80 drc784095 ( .a(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_45841) );
ao12f80 g784690 ( .a(n_3093), .b(n_3092), .c(n_2286), .o(n_47020) );
na02f80 g746970 ( .a(FE_OCP_RBN2168_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .o(n_33156) );
in01f80 g750971 ( .a(n_30102), .o(n_30103) );
no02f80 g773100 ( .a(n_7759), .b(n_7711), .o(n_8096) );
na02f80 g740502 ( .a(n_39702), .b(n_39672), .o(n_39719) );
in01f80 g738846 ( .a(n_41324), .o(n_41339) );
no02f80 g756876 ( .a(n_24028), .b(n_23803), .o(n_24063) );
oa12f80 g751698 ( .a(n_28962), .b(n_28994), .c(n_28793), .o(n_29252) );
in01f80 newInst_3191 ( .a(newNet_1154), .o(newNet_3191) );
in01f80 FE_OCP_RBC2304_n_7817 ( .a(FE_OCP_RBN2303_n_7817), .o(FE_OCP_RBN2304_n_7817) );
no02f80 g772402 ( .a(n_8474), .b(FE_OCP_RBN3467_n_7886), .o(n_8529) );
na02f80 g736723 ( .a(n_43139), .b(n_43228), .o(n_43281) );
in01f80 g755104 ( .a(n_25319), .o(n_25320) );
ao12f80 g764933 ( .a(n_16312), .b(n_16264), .c(n_16384), .o(n_16385) );
na02f80 g780496 ( .a(n_977), .b(n_898), .o(n_982) );
in01f80 g738092 ( .a(n_42089), .o(n_42090) );
na02f80 FE_RC_3567_0 ( .a(FE_OCP_DRV_N1566_n_28654), .b(n_29773), .o(FE_RN_1549_0) );
ao12f80 g755405 ( .a(n_24626), .b(n_24701), .c(n_24466), .o(n_24702) );
no02f80 g773648 ( .a(n_7354), .b(n_7353), .o(n_7368) );
in01f80 newInst_2154 ( .a(newNet_2153), .o(newNet_2154) );
ao12f80 g776524 ( .a(n_4331), .b(n_4553), .c(n_4404), .o(n_4710) );
no02f80 FE_RC_365_0 ( .a(FE_RN_110_0), .b(n_374), .o(n_454) );
no02f80 g739609 ( .a(FE_OCP_RBN3338_n_44610), .b(delay_xor_ln22_unr28_stage10_stallmux_q_0_), .o(n_40601) );
no02f80 g766786 ( .a(n_14044), .b(FE_OCP_RBN1923_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_14045) );
na02f80 g750753 ( .a(n_29316), .b(n_29168), .o(n_29339) );
oa22f80 g757767 ( .a(n_22511), .b(n_22508), .c(n_22531), .d(n_22469), .o(n_22631) );
in01f80 newInst_2773 ( .a(newNet_2599), .o(newNet_2773) );
in01f80 FE_OFC781_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN781_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
no02f80 g765869 ( .a(n_14793), .b(n_14265), .o(n_14861) );
in01f80 FE_RC_2732_0 ( .a(n_22927), .o(FE_RN_1157_0) );
no02f80 g776733 ( .a(n_4075), .b(n_4003), .o(n_4235) );
in01f80 g763186 ( .a(n_17289), .o(n_17560) );
in01f80 g765665 ( .a(n_15071), .o(n_15072) );
na02f80 g775496 ( .a(n_5650), .b(n_5572), .o(n_5719) );
no02f80 g776619 ( .a(n_4220), .b(n_4165), .o(n_4259) );
ao12f80 g750158 ( .a(n_29841), .b(n_29913), .c(n_28996), .o(n_29951) );
na02f80 g761703 ( .a(n_18855), .b(FE_OCP_DRV_N1544_n_18854), .o(n_18887) );
in01f80 g759991 ( .a(n_20414), .o(n_20415) );
in01f80 FE_OCP_RBC3010_n_31117 ( .a(FE_OCP_RBN3007_n_31117), .o(FE_OCP_RBN3010_n_31117) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_22_ ( .ck(newNet_2188), .d(n_1144), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_22_) );
ao12f80 g764944 ( .a(n_15541), .b(n_15610), .c(n_15609), .o(n_15683) );
no02f80 g744938 ( .a(n_36385), .b(n_36154), .o(n_36420) );
in01f80 newInst_3389 ( .a(newNet_3388), .o(newNet_3389) );
na02f80 g743040 ( .a(n_37149), .b(n_37039), .o(n_37178) );
oa12f80 g738145 ( .a(n_41721), .b(n_42027), .c(n_41658), .o(n_42057) );
in01f80 g761555 ( .a(n_19022), .o(n_19023) );
oa12f80 g749682 ( .a(n_31347), .b(n_31457), .c(n_31456), .o(n_31512) );
oa12f80 g771884 ( .a(n_7569), .b(n_8747), .c(n_8742), .o(n_8769) );
na02f80 g747787 ( .a(n_32000), .b(n_31688), .o(n_32111) );
no02f80 g770880 ( .a(n_9853), .b(n_9868), .o(n_9869) );
in01f80 g758166 ( .a(n_22083), .o(n_22045) );
in01f80 g759240 ( .a(n_21306), .o(n_21307) );
in01f80 g775360 ( .a(n_5609), .o(n_5610) );
no02f80 g738063 ( .a(n_42088), .b(n_41882), .o(n_42118) );
in01f80 g761774 ( .a(n_19339), .o(n_19401) );
no02f80 g763439 ( .a(n_16912), .b(n_15995), .o(n_17027) );
oa22f80 g781282 ( .a(n_67), .b(n_46055), .c(n_7), .d(beta_6), .o(n_123) );
in01f80 g742929 ( .a(n_37065), .o(n_37066) );
no02f80 g738488 ( .a(FE_OCP_RBN2317_n_41420), .b(n_41347), .o(n_41588) );
ao22s80 g740565 ( .a(FE_OCP_RBN2928_n_39614), .b(n_45840), .c(n_39614), .d(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39676) );
no02f80 g753856 ( .a(n_26334), .b(n_26299), .o(n_26469) );
no02f80 g749606 ( .a(n_30375), .b(n_30019), .o(n_30407) );
oa22f80 g748048 ( .a(n_31668), .b(n_31556), .c(n_31669), .d(n_31557), .o(n_31750) );
in01f80 g755400 ( .a(n_24913), .o(n_24914) );
no02f80 g758853 ( .a(n_21703), .b(n_21463), .o(n_21730) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_19_ ( .ck(newNet_2102), .d(n_6243), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_) );
oa22f80 g748516 ( .a(n_31585), .b(n_31647), .c(n_31586), .d(n_31646), .o(n_31715) );
in01f80 g756507 ( .a(n_23680), .o(n_23681) );
no02f80 g761266 ( .a(n_20012), .b(n_19953), .o(n_20013) );
no02f80 g750125 ( .a(FE_OCP_RBN2571_n_29922), .b(FE_OCP_RBN2328_n_29378), .o(n_30258) );
no02f80 g744205 ( .a(n_36133), .b(n_35620), .o(n_36258) );
in01f80 newInst_1626 ( .a(newNet_1305), .o(newNet_1626) );
na02f80 g773818 ( .a(n_7101), .b(n_6986), .o(n_7137) );
na02f80 FE_RC_2452_0 ( .a(n_41949), .b(n_41947), .o(FE_RN_981_0) );
na02f80 g769251 ( .a(n_11475), .b(FE_OCP_RBN2891_n_10568), .o(n_11516) );
in01f80 newInst_1210 ( .a(newNet_1209), .o(newNet_1210) );
in01f80 g739242 ( .a(n_40954), .o(n_40955) );
in01f80 newInst_525 ( .a(newNet_524), .o(newNet_525) );
in01f80 newInst_1743 ( .a(newNet_1742), .o(newNet_1743) );
no02f80 g777302 ( .a(n_4219), .b(FE_OFN819_n_4298), .o(n_4576) );
in01f80 newInst_3516 ( .a(newNet_3515), .o(newNet_3516) );
in01f80 newInst_2160 ( .a(newNet_810), .o(newNet_2160) );
in01f80 g754126 ( .a(n_26974), .o(n_26949) );
in01f80 g777854 ( .a(n_3238), .o(n_3287) );
in01f80 g778641 ( .a(n_2335), .o(n_2321) );
in01f80 newInst_3492 ( .a(newNet_2085), .o(newNet_3492) );
oa12f80 g752117 ( .a(n_28621), .b(n_28620), .c(n_28619), .o(n_28984) );
ao22s80 FE_RC_842_0 ( .a(n_42166), .b(n_42157), .c(n_42156), .d(n_42173), .o(n_42179) );
in01f80 g768976 ( .a(n_12281), .o(n_12213) );
na02f80 FE_RC_1313_0 ( .a(FE_RN_386_0), .b(n_3775), .o(n_47013) );
na02f80 g765838 ( .a(n_14927), .b(n_14899), .o(n_14928) );
na02f80 g767498 ( .a(n_13265), .b(FE_OCP_DRV_N3152_n_13264), .o(n_13302) );
na02f80 g778333 ( .a(n_2664), .b(n_2438), .o(n_2665) );
in01f80 FE_OCP_RBC3266_n_45224 ( .a(FE_OCP_RBN3267_n_45224), .o(FE_OCP_RBN3266_n_45224) );
na02f80 g777056 ( .a(n_3843), .b(n_3524), .o(n_3844) );
ao12f80 g741224 ( .a(n_38997), .b(FE_OCP_RBN3579_n_44944), .c(n_38907), .o(n_39320) );
ao22s80 g780397 ( .a(n_883), .b(FE_OFN760_n_45813), .c(n_834), .d(n_1203), .o(n_916) );
na02f80 g776429 ( .a(n_4586), .b(n_4199), .o(n_4677) );
na02f80 g752227 ( .a(n_28539), .b(n_28079), .o(n_28592) );
in01f80 FE_OCP_RBC3018_n_31117 ( .a(FE_OCP_RBN3015_n_31117), .o(FE_OCP_RBN3018_n_31117) );
na02f80 g741548 ( .a(n_38714), .b(n_38713), .o(n_38742) );
ao12f80 g765253 ( .a(n_15522), .b(n_15521), .c(n_15520), .o(n_15884) );
in01f80 g748805 ( .a(n_32558), .o(n_32449) );
no02f80 g770046 ( .a(n_10732), .b(n_10733), .o(n_10767) );
na02f80 g776886 ( .a(n_3950), .b(n_3932), .o(n_4168) );
in01f80 FE_OCP_RBC2488_n_3338 ( .a(n_3338), .o(FE_OCP_RBN2488_n_3338) );
ao22s80 FE_RC_1716_0 ( .a(n_16865), .b(n_17083), .c(n_16864), .d(n_17123), .o(n_17334) );
ms00f80 cos_out_reg_1_ ( .ck(newNet_3727), .d(n_43288), .o(cos_out_1) );
oa22f80 FE_RC_1273_0 ( .a(n_14114), .b(FE_OCP_RBN2250_n_13017), .c(n_13515), .d(FE_OCP_RBN2447_n_14114), .o(n_14271) );
oa22f80 FE_RC_3252_0 ( .a(n_11279), .b(n_11296), .c(n_11275), .d(n_11274), .o(n_11377) );
in01f80 g736781 ( .a(n_43394), .o(n_43395) );
no02f80 g746229 ( .a(n_33645), .b(n_33621), .o(n_33715) );
no02f80 g766068 ( .a(n_14689), .b(n_12795), .o(n_14971) );
in01f80 g751494 ( .a(n_28624), .o(n_28625) );
no02f80 g766894 ( .a(n_13877), .b(FE_OCPN1007_n_13962), .o(n_14425) );
oa12f80 g736425 ( .a(n_346), .b(n_43748), .c(FE_OFN2_n_43918), .o(n_43796) );
no02f80 g737464 ( .a(n_42637), .b(n_42684), .o(n_42715) );
in01f80 g743168 ( .a(n_36912), .o(n_36913) );
in01f80 FE_OCPC878_n_44734 ( .a(FE_OCP_RBN3366_n_44722), .o(FE_OCPN878_n_44734) );
na02f80 g766174 ( .a(n_14836), .b(n_14295), .o(n_14868) );
in01f80 newInst_3367 ( .a(newNet_3366), .o(newNet_3367) );
in01f80 g778702 ( .a(n_2258), .o(n_2259) );
no02f80 g739146 ( .a(n_40913), .b(n_40746), .o(n_40926) );
ao22s80 g778406 ( .a(n_45486), .b(n_2069), .c(n_45487), .d(n_2068), .o(n_3217) );
na02f80 g754895 ( .a(n_25210), .b(n_24217), .o(n_25302) );
no02f80 g763576 ( .a(FE_OCP_RBN3079_n_16977), .b(n_16866), .o(n_17451) );
in01f80 newInst_672 ( .a(newNet_671), .o(newNet_672) );
in01f80 g755181 ( .a(n_25175), .o(n_25203) );
in01f80 g746078 ( .a(n_33785), .o(n_33786) );
in01f80 newInst_446 ( .a(newNet_445), .o(newNet_446) );
in01f80 newInst_3074 ( .a(newNet_3073), .o(newNet_3074) );
in01f80 g736928 ( .a(n_43087), .o(n_43108) );
in01f80 g755839 ( .a(n_24366), .o(n_24395) );
no02f80 g760869 ( .a(n_19469), .b(n_19324), .o(n_19511) );
na02f80 g769771 ( .a(n_47269), .b(n_11142), .o(n_11168) );
in01f80 g738377 ( .a(n_41789), .o(n_41790) );
na02f80 g767086 ( .a(n_13610), .b(n_13609), .o(n_13611) );
no02f80 g778433 ( .a(n_2828), .b(FE_OCPN1234_n_2414), .o(n_2565) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_13_ ( .ck(newNet_977), .d(n_22892), .o(delay_xor_ln21_unr15_stage6_stallmux_q_13_) );
no02f80 g759971 ( .a(n_20988), .b(n_20987), .o(n_20989) );
in01f80 newInst_2403 ( .a(newNet_2402), .o(newNet_2403) );
in01f80 newInst_2265 ( .a(newNet_2264), .o(newNet_2265) );
in01f80 newInst_126 ( .a(newNet_125), .o(newNet_126) );
na02f80 g745754 ( .a(n_34238), .b(FE_OCP_RBN2283_n_33846), .o(n_34259) );
no02f80 g739074 ( .a(n_41064), .b(FE_OCP_RBN2161_n_40687), .o(n_41087) );
na02f80 FE_RC_2873_0 ( .a(FE_RN_1240_0), .b(FE_OCP_RBN3561_n_29857), .o(n_29952) );
in01f80 newInst_1310 ( .a(newNet_151), .o(newNet_1310) );
no02f80 g755135 ( .a(n_25373), .b(n_25531), .o(n_25532) );
in01f80 FE_OCP_RBC3063_n_11325 ( .a(n_11325), .o(FE_OCP_RBN3063_n_11325) );
in01f80 g762454 ( .a(n_18003), .o(n_18004) );
in01f80 newInst_1346 ( .a(newNet_1345), .o(newNet_1346) );
in01f80 FE_OCP_RBC2141_FE_OCPN861_n_45450 ( .a(FE_OCPN861_n_45450), .o(FE_OCP_RBN2141_FE_OCPN861_n_45450) );
in01f80 g759621 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_21453) );
ao22s80 g757176 ( .a(n_23493), .b(n_22880), .c(n_23492), .d(n_22881), .o(n_23645) );
no02f80 g764699 ( .a(n_15853), .b(n_15404), .o(n_15854) );
no02f80 g746120 ( .a(n_33675), .b(n_34037), .o(n_33698) );
no02f80 g736839 ( .a(n_43018), .b(n_42249), .o(n_43042) );
in01f80 g749421 ( .a(n_30622), .o(n_30672) );
oa12f80 g761294 ( .a(n_19649), .b(n_19830), .c(n_19337), .o(n_19832) );
in01f80 FE_OCP_RBC3461_n_7886 ( .a(n_7886), .o(FE_OCP_RBN3461_n_7886) );
no02f80 g747981 ( .a(n_33046), .b(n_33045), .o(n_33047) );
in01f80 FE_OCPC3769_FE_OCP_RBN2375_n_8221 ( .a(FE_OCPN3768_FE_OCP_RBN2375_n_8221), .o(FE_OCPN3769_FE_OCP_RBN2375_n_8221) );
no02f80 g755684 ( .a(n_25371), .b(cordic_combinational_sub_ln23_0_unr20_z_0_), .o(n_25370) );
ao12f80 g768933 ( .a(n_12311), .b(FE_OCPN867_n_45697), .c(delay_xor_ln22_unr9_stage4_stallmux_q_10_), .o(n_11938) );
no02f80 g769823 ( .a(n_11083), .b(n_11085), .o(n_11114) );
na02f80 g745237 ( .a(n_35681), .b(n_35584), .o(n_36226) );
no02f80 g766112 ( .a(n_14540), .b(n_13515), .o(n_14606) );
in01f80 g747705 ( .a(n_33703), .o(n_33704) );
na02f80 g759427 ( .a(n_20973), .b(n_20571), .o(n_20974) );
na02f80 g776378 ( .a(n_4671), .b(FE_OCP_RBN2538_n_3645), .o(n_4672) );
no02f80 g772998 ( .a(n_7730), .b(n_7832), .o(n_7833) );
na02f80 g755618 ( .a(n_24566), .b(n_23875), .o(n_24598) );
na02f80 g766824 ( .a(n_14488), .b(n_14339), .o(n_15398) );
in01f80 FE_OCP_RBC2630_n_14912 ( .a(n_14912), .o(FE_OCP_RBN2630_n_14912) );
no02f80 g752037 ( .a(n_28117), .b(n_28029), .o(n_28144) );
no02f80 g738057 ( .a(n_42133), .b(n_42132), .o(n_42134) );
no02f80 g740687 ( .a(n_39484), .b(n_39483), .o(n_39485) );
na02f80 g780755 ( .a(n_548), .b(n_389), .o(n_576) );
oa12f80 g776516 ( .a(n_3782), .b(n_3896), .c(n_3692), .o(n_4054) );
oa12f80 g745088 ( .a(n_34686), .b(n_34714), .c(n_34685), .o(n_35742) );
no02f80 g779729 ( .a(n_1575), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_19_), .o(n_1801) );
no02f80 g778120 ( .a(n_2805), .b(n_2208), .o(n_2820) );
in01f80 g745866 ( .a(n_34266), .o(n_34267) );
in01f80 FE_OCP_RBC2149_FE_OCPN861_n_45450 ( .a(FE_OCP_RBN2146_FE_OCPN861_n_45450), .o(FE_OCP_RBN2149_FE_OCPN861_n_45450) );
in01f80 FE_RC_2385_0 ( .a(n_42285), .o(FE_RN_932_0) );
oa12f80 g738048 ( .a(n_42142), .b(n_42145), .c(n_42141), .o(n_42390) );
in01f80 FE_RC_3145_0 ( .a(n_25755), .o(FE_RN_1396_0) );
oa12f80 g774255 ( .a(n_6789), .b(n_6773), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_20_), .o(n_6851) );
in01f80 g761229 ( .a(n_19200), .o(n_19308) );
na02f80 g774017 ( .a(n_7179), .b(n_7224), .o(n_7419) );
no02f80 g771892 ( .a(n_8739), .b(n_8697), .o(n_8786) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_20_ ( .ck(newNet_2389), .d(n_36414), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_) );
na02f80 g757938 ( .a(n_22268), .b(n_22351), .o(n_22352) );
no02f80 g767351 ( .a(n_13335), .b(FE_OCP_RBN3416_n_12739), .o(n_13368) );
oa12f80 g775607 ( .a(n_5152), .b(FE_OCP_RBN2897_n_45484), .c(n_5149), .o(n_5361) );
in01f80 g746698 ( .a(n_33113), .o(n_33068) );
no02f80 g742864 ( .a(n_37343), .b(n_37163), .o(n_37253) );
in01f80 newInst_3339 ( .a(newNet_3338), .o(newNet_3339) );
in01f80 FE_OCP_RBC1223_n_22914 ( .a(n_22914), .o(FE_OCP_RBN1223_n_22914) );
in01f80 FE_OCP_RBC2572_n_29922 ( .a(FE_OCP_RBN2570_n_29922), .o(FE_OCP_RBN2572_n_29922) );
oa12f80 g751275 ( .a(FE_OCPN1032_n_28448), .b(n_28748), .c(FE_OCPN1030_n_28423), .o(n_28791) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_24_ ( .ck(newNet_2276), .d(n_40544), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_24_) );
no02f80 g739970 ( .a(n_40333), .b(n_40133), .o(n_40368) );
in01f80 FE_OCP_RBC2337_n_8269 ( .a(n_8269), .o(FE_OCP_RBN2337_n_8269) );
no02f80 g784066 ( .a(n_679), .b(n_7), .o(n_45808) );
na02f80 FE_RC_1987_0 ( .a(n_13777), .b(FE_RN_647_0), .o(FE_RN_648_0) );
in01f80 g736709 ( .a(n_43405), .o(n_43406) );
na02f80 g764746 ( .a(n_15739), .b(n_44052), .o(n_15808) );
in01f80 g775486 ( .a(n_5721), .o(n_5673) );
oa12f80 g767720 ( .a(n_12491), .b(n_12655), .c(n_12438), .o(n_12713) );
na02f80 FE_RC_1789_0 ( .a(FE_RN_523_0), .b(FE_RN_525_0), .o(FE_RN_526_0) );
no02f80 g750762 ( .a(n_29195), .b(n_29166), .o(n_29262) );
no02f80 g746180 ( .a(n_33804), .b(n_33451), .o(n_33869) );
in01f80 g741885 ( .a(n_38434), .o(n_38404) );
oa22f80 FE_RC_961_0 ( .a(n_32566), .b(n_32516), .c(n_28336), .d(n_32465), .o(n_32567) );
no02f80 g752336 ( .a(n_44723), .b(delay_xor_ln21_unr18_stage7_stallmux_q_6_), .o(n_27999) );
oa12f80 g746474 ( .a(n_34940), .b(n_34891), .c(n_34666), .o(n_35187) );
in01f80 FE_OCPC1453_n_18559 ( .a(n_18559), .o(FE_OCPN1453_n_18559) );
na02f80 g779034 ( .a(n_2063), .b(n_1891), .o(n_2058) );
in01f80 FE_RC_1599_0 ( .a(n_27204), .o(FE_RN_447_0) );
na02f80 g760692 ( .a(n_19658), .b(n_19704), .o(n_19722) );
in01f80 newInst_1255 ( .a(newNet_1254), .o(newNet_1255) );
in01f80 newInst_2813 ( .a(newNet_2812), .o(newNet_2813) );
na02f80 g756006 ( .a(FE_OCP_RBN2525_n_24902), .b(n_24257), .o(n_25003) );
no02f80 g778075 ( .a(n_2972), .b(n_2867), .o(n_3035) );
in01f80 newInst_1407 ( .a(newNet_1406), .o(newNet_1407) );
in01f80 newInst_1115 ( .a(newNet_1114), .o(newNet_1115) );
na02f80 g745846 ( .a(n_35373), .b(n_35372), .o(n_35374) );
na02f80 FE_RC_468_0 ( .a(FE_RN_137_0), .b(n_28386), .o(n_28453) );
oa12f80 g740808 ( .a(n_39061), .b(n_39264), .c(n_38885), .o(n_39311) );
in01f80 g759319 ( .a(n_21074), .o(n_21183) );
ao12f80 g757060 ( .a(n_23086), .b(n_23546), .c(n_23051), .o(n_23648) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_2_ ( .ck(newNet_2726), .d(n_15168), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_2_) );
no02f80 g755856 ( .a(n_24340), .b(n_24016), .o(n_24363) );
in01f80 g750865 ( .a(n_29154), .o(n_29210) );
in01f80 newInst_2212 ( .a(newNet_2211), .o(newNet_2212) );
na02f80 g759520 ( .a(n_20930), .b(n_20903), .o(n_20959) );
na02f80 g751422 ( .a(n_28475), .b(n_28467), .o(n_28511) );
in01f80 FE_RC_2448_0 ( .a(n_13312), .o(FE_RN_978_0) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_14_ ( .ck(newNet_842), .d(n_1300), .o(delay_xor_ln21_unr3_stage2_stallmux_q_14_) );
no02f80 g776311 ( .a(n_4703), .b(n_4374), .o(n_4814) );
in01f80 g754544 ( .a(n_26738), .o(n_26739) );
in01f80 g755752 ( .a(n_24489), .o(n_24490) );
in01f80 g757791 ( .a(n_22450), .o(n_22543) );
in01f80 g766381 ( .a(n_14238), .o(n_14239) );
in01f80 FE_OCP_RBC2934_n_31010 ( .a(n_31010), .o(FE_OCP_RBN2934_n_31010) );
in01f80 g751438 ( .a(n_28530), .o(n_28531) );
in01f80 g765277 ( .a(n_15785), .o(n_15881) );
na02f80 g772359 ( .a(n_8521), .b(n_8477), .o(n_8545) );
na02f80 g751536 ( .a(n_28460), .b(n_27860), .o(n_28719) );
no02f80 g756616 ( .a(n_24078), .b(n_24149), .o(n_24195) );
oa12f80 g769957 ( .a(n_10825), .b(n_10857), .c(FE_OCP_RBN3653_n_10100), .o(n_10946) );
na02f80 g754070 ( .a(n_26166), .b(n_26147), .o(n_26318) );
na02f80 g747319 ( .a(n_32529), .b(n_44962), .o(n_32791) );
na02f80 g754906 ( .a(n_25481), .b(n_24518), .o(n_25564) );
no02f80 g738751 ( .a(n_41384), .b(n_41383), .o(n_41397) );
no02f80 g756025 ( .a(n_25188), .b(n_25027), .o(n_25134) );
ms00f80 delay_sub_ln21_0_unr17_stage7_stallmux_q_reg_15_ ( .ck(newNet_2581), .d(n_27443), .o(delay_sub_ln21_0_unr17_stage7_stallmux_q_15_) );
ao12f80 g763093 ( .a(n_17546), .b(n_17545), .c(n_17544), .o(n_18953) );
in01f80 g755352 ( .a(n_24860), .o(n_24923) );
na02f80 g768694 ( .a(n_12108), .b(n_11852), .o(n_12154) );
no02f80 g758673 ( .a(n_21743), .b(n_21553), .o(n_21793) );
ao22s80 FE_RC_3783_0 ( .a(n_17268), .b(n_17446), .c(n_17269), .d(n_17452), .o(n_17587) );
na02f80 g761698 ( .a(n_18853), .b(n_18432), .o(n_18916) );
in01f80 newInst_2301 ( .a(newNet_2300), .o(newNet_2301) );
na02f80 g768817 ( .a(n_44859), .b(n_11729), .o(n_11921) );
in01f80 newInst_2034 ( .a(newNet_2033), .o(newNet_2034) );
in01f80 newInst_3404 ( .a(newNet_3403), .o(newNet_3404) );
na02f80 g779786 ( .a(n_1780), .b(n_1131), .o(n_1442) );
in01f80 g766343 ( .a(n_14328), .o(n_14327) );
no02f80 g764586 ( .a(n_15998), .b(n_15985), .o(n_16077) );
in01f80 newInst_757 ( .a(newNet_756), .o(newNet_757) );
no02f80 g748390 ( .a(n_31476), .b(n_30507), .o(n_31555) );
no02f80 g758902 ( .a(n_46966), .b(n_21728), .o(n_21761) );
no02f80 g760489 ( .a(n_19923), .b(n_18677), .o(n_20029) );
in01f80 FE_OCP_RBC2598_n_34388 ( .a(n_34388), .o(FE_OCP_RBN2598_n_34388) );
na02f80 g751547 ( .a(n_28419), .b(delay_add_ln22_unr17_stage7_stallmux_q_14_), .o(n_28474) );
in01f80 g774295 ( .a(n_6642), .o(n_6571) );
in01f80 g763650 ( .a(n_46975), .o(n_16895) );
na02f80 g745400 ( .a(n_34226), .b(n_34209), .o(n_34210) );
in01f80 newInst_2595 ( .a(newNet_2594), .o(newNet_2595) );
na02f80 g768436 ( .a(n_12374), .b(n_12397), .o(n_12560) );
na02f80 g742837 ( .a(n_37270), .b(n_37096), .o(n_37255) );
na02f80 g775453 ( .a(n_5433), .b(n_5336), .o(n_5526) );
in01f80 newInst_3648 ( .a(newNet_3451), .o(newNet_3648) );
in01f80 FE_OCP_RBC2351_n_38534 ( .a(n_38534), .o(FE_OCP_RBN2351_n_38534) );
no02f80 g774372 ( .a(n_6593), .b(n_6562), .o(n_6672) );
na03f80 g745021 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_4_), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_3_), .o(n_36434) );
no02f80 g778415 ( .a(n_2722), .b(n_2137), .o(n_2786) );
na02f80 g753242 ( .a(n_27167), .b(n_25907), .o(n_27216) );
no02f80 g755811 ( .a(FE_OCP_RBN2334_n_24359), .b(n_24288), .o(n_24427) );
in01f80 newInst_1480 ( .a(newNet_1479), .o(newNet_1480) );
na02f80 g760572 ( .a(n_19806), .b(n_18230), .o(n_19843) );
no02f80 g761540 ( .a(n_18755), .b(n_18682), .o(n_18828) );
ao22s80 g776747 ( .a(FE_OCP_RBN2624_n_3848), .b(n_3029), .c(n_3848), .d(n_3082), .o(n_4011) );
in01f80 g757168 ( .a(n_23671), .o(n_23700) );
ao12f80 g752459 ( .a(n_28352), .b(n_28378), .c(n_28351), .o(n_28835) );
no02f80 g764619 ( .a(n_15951), .b(n_14524), .o(n_15952) );
in01f80 g757773 ( .a(delay_xor_ln22_unr15_stage6_stallmux_q_0_), .o(n_22517) );
na02f80 g774282 ( .a(n_6705), .b(n_6628), .o(n_6706) );
ao12f80 g767398 ( .a(n_13402), .b(n_13401), .c(n_13400), .o(n_13478) );
in01f80 g752520 ( .a(n_27743), .o(n_27793) );
in01f80 newInst_1079 ( .a(newNet_1078), .o(newNet_1079) );
oa22f80 g769012 ( .a(n_12219), .b(FE_OCP_RBN1925_cordic_combinational_sub_ln23_0_unr12_z_0__), .c(n_12218), .d(FE_OCP_RBN1926_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(n_12671) );
na02f80 g754409 ( .a(FE_OCP_RBN2763_n_25732), .b(n_25760), .o(n_25761) );
in01f80 g765364 ( .a(n_16253), .o(n_16254) );
in01f80 FE_OCP_RBC2116_n_45224 ( .a(FE_OCP_RBN3266_n_45224), .o(FE_OCP_RBN2116_n_45224) );
na02f80 FE_RC_3604_0 ( .a(FE_RN_1574_0), .b(n_20542), .o(FE_RN_1575_0) );
na02f80 g753249 ( .a(n_27287), .b(n_27416), .o(n_27527) );
no02f80 g775091 ( .a(n_5987), .b(n_5709), .o(n_6009) );
na02f80 g763525 ( .a(n_15912), .b(FE_OCP_RBN1208_n_16814), .o(n_17032) );
no02f80 FE_RC_4074_0 ( .a(n_36011), .b(FE_RN_1775_0), .o(n_36474) );
na02f80 g767555 ( .a(n_13012), .b(n_13005), .o(n_13094) );
no02f80 g744156 ( .a(n_35553), .b(n_35520), .o(n_35670) );
no02f80 g742190 ( .a(n_44869), .b(n_38209), .o(n_37874) );
in01f80 g778811 ( .a(n_3106), .o(n_3862) );
oa12f80 g784698 ( .a(FE_OFN751_n_45003), .b(n_20250), .c(n_20229), .o(n_47174) );
in01f80 FE_OCP_RBC2874_n_10477 ( .a(n_10477), .o(FE_OCP_RBN2874_n_10477) );
oa22f80 g779335 ( .a(FE_OCP_RBN2157_n_1614), .b(n_1438), .c(n_1614), .d(n_1439), .o(n_1701) );
in01f80 g736887 ( .a(n_43593), .o(n_43594) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_23_ ( .ck(newNet_2279), .d(n_40525), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_23_) );
no02f80 g768288 ( .a(n_12641), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_), .o(n_12656) );
no02f80 g755516 ( .a(n_24651), .b(n_24622), .o(n_24750) );
in01f80 FE_OCP_RBC2326_n_29378 ( .a(n_29378), .o(FE_OCP_RBN2326_n_29378) );
in01f80 FE_OCP_RBC2151_n_22822 ( .a(n_22822), .o(FE_OCP_RBN2151_n_22822) );
oa22f80 FE_RC_3436_0 ( .a(n_32287), .b(n_32519), .c(n_28336), .d(n_32469), .o(n_32569) );
in01f80 g745349 ( .a(n_36157), .o(n_36158) );
no02f80 g755881 ( .a(n_25086), .b(n_25085), .o(n_25087) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_16_ ( .ck(newNet_3637), .d(n_16810), .o(delay_add_ln22_unr11_stage5_stallmux_q_16_) );
in01f80 newInst_3238 ( .a(newNet_3237), .o(newNet_3238) );
in01f80 g748492 ( .a(n_31783), .o(n_31819) );
in01f80 FE_RC_519_0 ( .a(n_24182), .o(FE_RN_162_0) );
na02f80 g763158 ( .a(n_17048), .b(n_16909), .o(n_17092) );
in01f80 FE_OCPC3787_n_22156 ( .a(FE_OCPN3786_n_22156), .o(FE_OCPN3787_n_22156) );
in01f80 newInst_659 ( .a(newNet_12), .o(newNet_659) );
no02f80 g780779 ( .a(n_534), .b(n_533), .o(n_535) );
no02f80 g773605 ( .a(n_7381), .b(n_7374), .o(n_7375) );
oa22f80 g750039 ( .a(n_29896), .b(n_29501), .c(n_29869), .d(n_29530), .o(n_30347) );
na02f80 g765573 ( .a(n_15142), .b(n_14821), .o(n_15403) );
na02f80 g779010 ( .a(n_2106), .b(n_2095), .o(n_2096) );
oa12f80 g747133 ( .a(n_32733), .b(n_32774), .c(n_32695), .o(n_32799) );
na02f80 g773756 ( .a(n_7218), .b(n_7041), .o(n_7219) );
in01f80 g756471 ( .a(n_23661), .o(n_23662) );
na02f80 g777607 ( .a(n_3530), .b(n_3552), .o(n_3674) );
in01f80 FE_RC_2435_0 ( .a(n_32712), .o(FE_RN_970_0) );
oa12f80 g741927 ( .a(n_37972), .b(n_38092), .c(n_37887), .o(n_38124) );
in01f80 g738459 ( .a(n_41851), .o(n_41852) );
in01f80 g779145 ( .a(n_1956), .o(n_1957) );
ms00f80 sin_out_reg_16_ ( .ck(newNet_73), .d(n_43873), .o(sin_out_16) );
ao22s80 g757408 ( .a(FE_OCP_RBN3823_n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .c(n_22939), .d(n_44061), .o(n_22992) );
in01f80 g737176 ( .a(n_43001), .o(n_43007) );
in01f80 g765513 ( .a(n_15787), .o(n_15716) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_29_ ( .ck(newNet_1083), .d(n_11433), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_29_) );
in01f80 g764164 ( .a(n_16555), .o(n_16556) );
na02f80 g769970 ( .a(n_10995), .b(n_10956), .o(n_11045) );
oa12f80 g780809 ( .a(n_598), .b(n_597), .c(beta_0), .o(n_600) );
na02f80 g739592 ( .a(n_40641), .b(n_40654), .o(n_40642) );
na02f80 g763074 ( .a(n_17201), .b(n_17043), .o(n_17293) );
in01f80 g765383 ( .a(n_15578), .o(n_15516) );
oa12f80 g765179 ( .a(n_16343), .b(n_16342), .c(n_16341), .o(n_16408) );
in01f80 newInst_1513 ( .a(newNet_1512), .o(newNet_1513) );
oa12f80 g751282 ( .a(n_29743), .b(n_29742), .c(n_29741), .o(n_30030) );
no02f80 g774034 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_28_), .b(delay_add_ln22_unr5_stage3_stallmux_q_29_), .o(n_6707) );
na02f80 g775973 ( .a(n_5108), .b(n_5033), .o(n_5171) );
na02f80 g757780 ( .a(n_22482), .b(n_22347), .o(n_22536) );
in01f80 g770162 ( .a(n_46988), .o(n_10980) );
in01f80 FE_RC_2553_0 ( .a(FE_RN_206_0), .o(FE_RN_1046_0) );
in01f80 g778315 ( .a(n_2904), .o(n_2905) );
oa12f80 g742574 ( .a(n_37508), .b(n_37507), .c(n_37506), .o(n_38270) );
in01f80 g763615 ( .a(n_16864), .o(n_16865) );
in01f80 g743698 ( .a(n_36376), .o(n_36411) );
na02f80 g738086 ( .a(n_42107), .b(n_42542), .o(n_42106) );
no02f80 g767957 ( .a(n_12855), .b(n_12854), .o(n_12856) );
na02f80 g760389 ( .a(n_20099), .b(n_19884), .o(n_20148) );
na03f80 g784655 ( .a(n_12761), .b(n_12461), .c(n_12495), .o(n_46985) );
no02f80 g746219 ( .a(n_35087), .b(n_35086), .o(n_35088) );
na02f80 g738509 ( .a(FE_OCP_RBN2314_n_41420), .b(n_41219), .o(n_41632) );
oa12f80 g748680 ( .a(n_32446), .b(n_32539), .c(n_32508), .o(n_32610) );
no02f80 g784389 ( .a(n_6305), .b(n_5341), .o(n_46195) );
na02f80 g744530 ( .a(n_35369), .b(n_35353), .o(n_35428) );
in01f80 g736446 ( .a(n_43822), .o(n_43790) );
no02f80 g753687 ( .a(n_26522), .b(n_25013), .o(n_26584) );
na03f80 FE_RC_3220_0 ( .a(n_11195), .b(n_11110), .c(n_11076), .o(n_11196) );
oa22f80 FE_RC_777_0 ( .a(FE_OCPN1011_n_7802), .b(n_8548), .c(FE_OCP_RBN3467_n_7886), .d(n_8549), .o(n_8696) );
na02f80 g758370 ( .a(n_22187), .b(n_20868), .o(n_22351) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_5_ ( .ck(newNet_2347), .d(n_35507), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_5_) );
na02f80 g754862 ( .a(n_25977), .b(n_25950), .o(n_25951) );
ao12f80 g781267 ( .a(n_7), .b(beta_24), .c(beta_23), .o(n_120) );
no02f80 g781233 ( .a(n_109), .b(n_68), .o(n_143) );
oa12f80 g745174 ( .a(n_34187), .b(n_34494), .c(n_34128), .o(n_34658) );
in01f80 g744000 ( .a(n_36268), .o(n_36269) );
ao12f80 g756225 ( .a(n_24708), .b(n_24707), .c(n_24706), .o(n_25136) );
in01f80 g776146 ( .a(n_4986), .o(n_5059) );
ao12f80 g765060 ( .a(n_15514), .b(n_16347), .c(n_15788), .o(n_15789) );
na02f80 FE_RC_2173_0 ( .a(n_26292), .b(n_26218), .o(FE_RN_774_0) );
in01f80 newInst_3478 ( .a(newNet_1413), .o(newNet_3478) );
oa12f80 g780738 ( .a(n_446), .b(n_596), .c(n_433), .o(n_608) );
no02f80 g740232 ( .a(n_39772), .b(n_39754), .o(n_39798) );
no02f80 g760127 ( .a(n_20428), .b(FE_OCPN1782_FE_OCP_RBN1701_n_19353), .o(n_20532) );
no02f80 g784763 ( .a(n_33594), .b(n_34037), .o(n_47249) );
oa12f80 g739849 ( .a(n_40090), .b(n_40265), .c(n_39954), .o(n_40300) );
no02f80 g773153 ( .a(n_7886), .b(n_7877), .o(n_7964) );
in01f80 g746915 ( .a(n_33151), .o(n_33200) );
na02f80 FE_RC_269_0 ( .a(FE_RN_80_0), .b(n_44275), .o(n_22170) );
in01f80 FE_OCP_RBC2405_n_24638 ( .a(FE_OCP_RBN2403_n_24638), .o(FE_OCP_RBN2405_n_24638) );
no02f80 g750400 ( .a(n_29645), .b(n_29644), .o(n_29660) );
in01f80 newInst_2960 ( .a(newNet_2941), .o(newNet_2960) );
in01f80 g747250 ( .a(n_32813), .o(n_32814) );
na02f80 g741089 ( .a(n_38883), .b(n_38868), .o(n_39002) );
in01f80 g738545 ( .a(n_41453), .o(n_41424) );
na02f80 g749770 ( .a(n_31572), .b(n_31280), .o(n_31631) );
in01f80 g756267 ( .a(n_24094), .o(n_24095) );
no02f80 g765983 ( .a(n_14672), .b(n_13404), .o(n_14697) );
ao22s80 FE_RC_2980_0 ( .a(n_29262), .b(FE_RN_1301_0), .c(n_29296), .d(n_29451), .o(n_29577) );
oa12f80 g769845 ( .a(n_10208), .b(n_11180), .c(n_10119), .o(n_11213) );
oa12f80 g775307 ( .a(n_5423), .b(n_44862), .c(n_5446), .o(n_5561) );
no02f80 g766028 ( .a(n_14662), .b(n_14661), .o(n_14741) );
in01f80 g765304 ( .a(n_15962), .o(n_15963) );
in01f80 newInst_609 ( .a(newNet_608), .o(newNet_609) );
oa12f80 g744330 ( .a(n_35440), .b(n_35503), .c(n_35465), .o(n_35556) );
in01f80 g780918 ( .a(n_560), .o(n_561) );
na04m80 FE_RC_3937_0 ( .a(n_22944), .b(n_22824), .c(FE_OCP_RBN2151_n_22822), .d(n_22866), .o(n_23044) );
na02f80 g767984 ( .a(n_13114), .b(n_13109), .o(n_13679) );
no02f80 g749307 ( .a(n_30727), .b(FE_OCPN1410_n_27014), .o(n_30760) );
no02f80 g752794 ( .a(n_28077), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_27_), .o(n_28129) );
in01f80 g761781 ( .a(n_18518), .o(n_18562) );
in01f80 g778929 ( .a(n_2170), .o(n_2171) );
in01f80 g776643 ( .a(n_4296), .o(n_4427) );
ao12f80 g769955 ( .a(n_10836), .b(n_11019), .c(FE_OCP_RBN3002_n_10805), .o(n_11096) );
oa12f80 g749700 ( .a(n_31229), .b(n_31228), .c(n_31227), .o(n_31293) );
na02f80 g756848 ( .a(n_23328), .b(n_23179), .o(n_23350) );
in01f80 FE_RC_3522_0 ( .a(n_34406), .o(FE_RN_1522_0) );
no02f80 g776179 ( .a(n_4895), .b(n_4424), .o(n_5024) );
na02f80 g778246 ( .a(n_2725), .b(n_3127), .o(n_2726) );
oa12f80 g748168 ( .a(n_32403), .b(n_32780), .c(n_32483), .o(n_32807) );
in01f80 newInst_1054 ( .a(newNet_1053), .o(newNet_1054) );
na02f80 g749763 ( .a(n_31115), .b(n_31089), .o(n_31227) );
oa12f80 g756944 ( .a(n_23864), .b(n_24188), .c(n_23802), .o(n_24628) );
in01f80 newInst_1171 ( .a(newNet_1170), .o(newNet_1171) );
in01f80 newInst_3345 ( .a(newNet_3344), .o(newNet_3345) );
in01f80 FE_OFC793_n_45813 ( .a(FE_OFN40_n_45813), .o(FE_OFN793_n_45813) );
na02f80 g777789 ( .a(n_3255), .b(n_3104), .o(n_3322) );
oa12f80 g747581 ( .a(n_33480), .b(n_33479), .c(n_33392), .o(n_34074) );
in01f80 g769326 ( .a(n_11974), .o(n_11893) );
ao12f80 g767302 ( .a(n_13672), .b(n_13678), .c(n_13671), .o(n_14256) );
na02f80 g748826 ( .a(n_31236), .b(n_31200), .o(n_31237) );
in01f80 g766437 ( .a(n_14123), .o(n_14124) );
in01f80 g748559 ( .a(n_31476), .o(n_31518) );
in01f80 g772802 ( .a(n_8133), .o(n_8134) );
na02f80 g758576 ( .a(n_21936), .b(n_21922), .o(n_21997) );
in01f80 g741590 ( .a(n_38662), .o(n_38663) );
in01f80 FE_RC_1362_0 ( .a(n_5426), .o(FE_RN_406_0) );
in01f80 fopt783174 ( .a(n_6487), .o(n_44711) );
in01f80 g757352 ( .a(n_23101), .o(n_23126) );
no02f80 g780596 ( .a(n_694), .b(n_719), .o(n_732) );
na02f80 g770954 ( .a(n_10041), .b(n_8429), .o(n_10162) );
oa12f80 g747115 ( .a(n_33445), .b(n_33953), .c(n_33572), .o(n_34022) );
no02f80 g742376 ( .a(n_37806), .b(n_37817), .o(n_37807) );
na02f80 g747739 ( .a(n_33417), .b(n_33415), .o(n_33416) );
no02f80 g737885 ( .a(n_42270), .b(n_42570), .o(n_42608) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_22_ ( .ck(newNet_333), .d(n_1309), .o(delay_xor_ln22_unr3_stage2_stallmux_q_22_) );
na02f80 g755335 ( .a(n_24787), .b(n_24705), .o(n_24900) );
no02f80 g773557 ( .a(n_7405), .b(n_7257), .o(n_7422) );
oa12f80 g750987 ( .a(n_30035), .b(n_29996), .c(n_29944), .o(n_30098) );
na02f80 g770177 ( .a(n_10795), .b(n_10773), .o(n_10820) );
in01f80 newInst_2239 ( .a(newNet_827), .o(newNet_2239) );
na02f80 g761317 ( .a(n_19981), .b(n_19901), .o(n_19982) );
in01f80 g756036 ( .a(n_24954), .o(n_24955) );
na02f80 g772496 ( .a(n_8400), .b(n_8292), .o(n_8415) );
in01f80 g745272 ( .a(n_36176), .o(n_36177) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_6_ ( .ck(newNet_2144), .d(n_934), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_6_) );
na03f80 FE_RC_3297_0 ( .a(n_34460), .b(n_34398), .c(n_34401), .o(n_34461) );
no02f80 g780478 ( .a(n_831), .b(n_754), .o(n_755) );
na02f80 g759586 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_21485) );
oa12f80 g739204 ( .a(n_40741), .b(n_40740), .c(n_40739), .o(n_40863) );
ao22s80 g771712 ( .a(n_8995), .b(FE_OCP_RBN3547_n_44575), .c(n_9032), .d(FE_OCP_RBN3552_n_44575), .o(n_9275) );
no02f80 g742766 ( .a(n_37389), .b(n_37205), .o(n_37390) );
no02f80 g739453 ( .a(n_44769), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_), .o(n_40904) );
ao12f80 g750967 ( .a(n_30097), .b(n_30166), .c(n_30165), .o(n_30185) );
in01f80 g774183 ( .a(n_6635), .o(n_6636) );
in01f80 g760102 ( .a(n_20215), .o(n_20216) );
ao22s80 g784438 ( .a(n_36902), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .c(n_36942), .d(n_46204), .o(n_46250) );
oa12f80 g743809 ( .a(n_35643), .b(n_36335), .c(n_35706), .o(n_36046) );
no02f80 g747335 ( .a(n_32810), .b(n_32684), .o(n_32685) );
na03f80 FE_RC_1060_0 ( .a(n_41730), .b(n_41749), .c(n_41748), .o(n_41750) );
in01f80 g779087 ( .a(n_2766), .o(n_2031) );
in01f80 g763617 ( .a(n_17471), .o(n_17541) );
na02f80 g767966 ( .a(FE_OCPN860_n_12880), .b(n_13163), .o(n_13251) );
na02f80 g774369 ( .a(n_6857), .b(n_6887), .o(n_7392) );
na02f80 g746481 ( .a(n_34814), .b(n_34810), .o(n_34942) );
in01f80 FE_OCP_RBC3267_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3267_n_45224) );
in01f80 g739309 ( .a(n_40902), .o(n_40903) );
oa22f80 FE_RC_25_0 ( .a(n_6078), .b(n_6130), .c(n_6059), .d(n_6115), .o(n_6214) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_10_ ( .ck(newNet_678), .d(n_46367), .o(delay_xor_ln21_unr9_stage4_stallmux_q_10_) );
oa22f80 g744622 ( .a(n_36571), .b(n_36164), .c(n_36572), .d(n_36165), .o(n_36641) );
na02f80 g779158 ( .a(n_1885), .b(n_1884), .o(n_1886) );
no02f80 g778265 ( .a(n_2920), .b(n_3857), .o(n_2982) );
oa12f80 g770634 ( .a(n_10242), .b(n_10355), .c(n_10190), .o(n_10377) );
na02f80 g749141 ( .a(n_31046), .b(n_31045), .o(n_31016) );
in01f80 g772689 ( .a(n_8211), .o(n_8212) );
in01f80 newInst_3311 ( .a(newNet_3310), .o(newNet_3311) );
oa22f80 g763966 ( .a(n_16851), .b(n_16300), .c(n_16850), .d(n_16301), .o(n_16967) );
in01f80 g778808 ( .a(n_3106), .o(n_4093) );
no02f80 g741491 ( .a(n_38743), .b(n_38715), .o(n_38758) );
in01f80 g764927 ( .a(n_15723), .o(n_15724) );
na02f80 g772018 ( .a(FE_OCP_RBN3647_n_44490), .b(n_9647), .o(n_9692) );
in01f80 g779747 ( .a(n_1527), .o(n_1518) );
oa12f80 g749490 ( .a(n_30203), .b(n_30498), .c(n_30202), .o(n_30558) );
no02f80 g740743 ( .a(n_39413), .b(n_39445), .o(n_39889) );
no02f80 g764288 ( .a(FE_OCP_RBN2906_n_16230), .b(n_14618), .o(n_16335) );
in01f80 FE_OCP_RBC2329_n_9003 ( .a(n_9003), .o(FE_OCP_RBN2329_n_9003) );
in01f80 g780121 ( .a(n_1188), .o(n_1186) );
in01f80 newInst_614 ( .a(newNet_613), .o(newNet_614) );
na02f80 g746469 ( .a(n_34498), .b(n_34553), .o(n_35017) );
na02f80 g781030 ( .a(sin_out_28), .b(FE_OFN4_n_43918), .o(n_322) );
na02f80 FE_RC_1568_0 ( .a(FE_RN_444_0), .b(FE_RN_445_0), .o(FE_RN_446_0) );
na02f80 g776452 ( .a(n_4588), .b(n_4587), .o(n_4649) );
in01f80 g758377 ( .a(n_21999), .o(n_22014) );
oa12f80 g779240 ( .a(n_1843), .b(n_1853), .c(n_1842), .o(n_1905) );
no02f80 g768831 ( .a(n_11941), .b(delay_add_ln22_unr8_stage4_stallmux_q_2_), .o(n_12069) );
na02f80 g757852 ( .a(n_22445), .b(n_22446), .o(n_22447) );
in01f80 g737665 ( .a(n_42659), .o(n_42660) );
na02f80 g772568 ( .a(n_8557), .b(n_8556), .o(n_8558) );
in01f80 g750817 ( .a(n_29144), .o(n_29145) );
in01f80 g754755 ( .a(n_25403), .o(n_25461) );
in01f80 g771558 ( .a(n_9441), .o(n_9442) );
no02f80 g736979 ( .a(FE_OCPN1246_n_43120), .b(n_42972), .o(n_43505) );
na02f80 g770750 ( .a(FE_OCP_RBN3654_n_10100), .b(n_10183), .o(n_10185) );
no02f80 g749063 ( .a(n_30890), .b(n_30887), .o(n_30891) );
na02f80 FE_RC_491_0 ( .a(FE_RN_144_0), .b(FE_RN_145_0), .o(FE_RN_146_0) );
na02f80 g736988 ( .a(n_43242), .b(n_42774), .o(n_43453) );
oa12f80 g772376 ( .a(FE_OCP_RBN2416_n_8293), .b(n_8392), .c(n_8460), .o(n_8553) );
in01f80 g750647 ( .a(n_29466), .o(n_29467) );
na02f80 g740095 ( .a(n_40187), .b(n_39924), .o(n_40289) );
in01f80 newInst_2750 ( .a(newNet_2749), .o(newNet_2750) );
in01f80 g770823 ( .a(n_9862), .o(n_10017) );
in01f80 newInst_1061 ( .a(newNet_454), .o(newNet_1061) );
no02f80 g745588 ( .a(FE_OCPN1732_n_34369), .b(FE_OCPN3749_n_34296), .o(n_34764) );
in01f80 g766607 ( .a(n_14115), .o(n_14049) );
oa12f80 g751855 ( .a(n_28919), .b(n_29068), .c(n_29067), .o(n_29028) );
in01f80 newInst_707 ( .a(newNet_706), .o(newNet_707) );
oa12f80 g771464 ( .a(n_7678), .b(n_8878), .c(n_8846), .o(n_8914) );
in01f80 newInst_2553 ( .a(newNet_2552), .o(newNet_2553) );
ao12f80 g738561 ( .a(n_41423), .b(n_41422), .c(n_41421), .o(n_41504) );
no02f80 g754268 ( .a(n_26688), .b(n_26716), .o(n_26717) );
ao12f80 g784122 ( .a(n_45874), .b(n_45846), .c(n_45866), .o(n_45875) );
in01f80 g768374 ( .a(n_12519), .o(n_12482) );
in01f80 g739796 ( .a(n_40425), .o(n_40426) );
in01f80 FE_OCP_DRV_C1537_n_13646 ( .a(n_13646), .o(FE_OCP_DRV_N1537_n_13646) );
oa12f80 g775071 ( .a(n_47270), .b(n_6036), .c(n_5891), .o(n_6112) );
ao12f80 g741844 ( .a(n_38255), .b(n_38363), .c(n_38316), .o(n_38394) );
na02f80 g763384 ( .a(FE_OCP_RBN3725_n_16975), .b(n_15983), .o(n_17221) );
no02f80 FE_RC_3091_0 ( .a(FE_RN_1364_0), .b(n_21424), .o(FE_RN_1365_0) );
in01f80 g736633 ( .a(n_43623), .o(n_43624) );
no02f80 g779818 ( .a(FE_OCP_RBN3248_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln23_unr3_stage2_stallmux_q), .o(n_1780) );
no02f80 g775895 ( .a(n_4991), .b(n_4952), .o(n_5163) );
ao12f80 g751500 ( .a(n_28608), .b(n_28458), .c(delay_sub_ln21_0_unr17_stage7_stallmux_q_19_), .o(n_28676) );
na02f80 g742110 ( .a(n_37995), .b(n_37620), .o(n_38050) );
na02f80 g741082 ( .a(n_39006), .b(n_39100), .o(n_39187) );
in01f80 g781005 ( .a(n_276), .o(n_277) );
no02f80 g747616 ( .a(n_32280), .b(n_31991), .o(n_32302) );
in01f80 newInst_1076 ( .a(newNet_1075), .o(newNet_1076) );
in01f80 g770595 ( .a(n_10292), .o(n_10293) );
na02f80 g745238 ( .a(n_34592), .b(n_34627), .o(n_34655) );
in01f80 FE_OCP_RBC3108_n_40586 ( .a(n_40586), .o(FE_OCP_RBN3108_n_40586) );
ao22s80 g736598 ( .a(n_43241), .b(n_43578), .c(n_43240), .d(n_43577), .o(n_43648) );
na02f80 g756299 ( .a(n_24609), .b(n_23862), .o(n_24610) );
no02f80 g741570 ( .a(n_45192), .b(n_38662), .o(n_38688) );
in01f80 g752719 ( .a(n_27239), .o(n_27240) );
in01f80 g738153 ( .a(n_42076), .o(n_42077) );
na02f80 g776416 ( .a(n_4608), .b(n_4561), .o(n_4562) );
no02f80 g744273 ( .a(n_44174), .b(n_35567), .o(n_35617) );
in01f80 FE_OCPC1256_n_13831 ( .a(FE_OCP_RBN2361_n_13818), .o(FE_OCPN1256_n_13831) );
in01f80 FE_OCP_RBC2704_n_9411 ( .a(n_9411), .o(FE_OCP_RBN2704_n_9411) );
ao22s80 FE_RC_393_0 ( .a(n_12647), .b(n_13299), .c(n_12648), .d(n_13298), .o(n_13388) );
in01f80 newInst_1562 ( .a(newNet_1561), .o(newNet_1562) );
na02f80 g741949 ( .a(n_38140), .b(n_38247), .o(n_38284) );
ao12f80 g777411 ( .a(n_2631), .b(n_3400), .c(n_2658), .o(n_3492) );
no02f80 FE_RC_2461_0 ( .a(n_13900), .b(n_13937), .o(FE_RN_987_0) );
no02f80 g741144 ( .a(n_38993), .b(n_38890), .o(n_38891) );
na02f80 g775770 ( .a(n_5003), .b(FE_OCPN846_n_4046), .o(n_5045) );
oa12f80 g759699 ( .a(n_21256), .b(n_21255), .c(cordic_combinational_sub_ln23_0_unr16_z_0_), .o(n_21338) );
no02f80 g749252 ( .a(n_30841), .b(n_30843), .o(n_30904) );
na02f80 g773423 ( .a(n_7559), .b(FE_OCP_RBN2226_n_7531), .o(n_7586) );
na02f80 g765200 ( .a(n_15272), .b(n_15273), .o(n_15274) );
in01f80 FE_OCP_RBC2354_n_13858 ( .a(FE_OCP_RBN1171_n_13858), .o(FE_OCP_RBN2354_n_13858) );
no02f80 g746348 ( .a(n_35633), .b(n_36111), .o(n_35108) );
na02f80 g738494 ( .a(FE_OCP_RBN2316_n_41420), .b(n_41628), .o(n_41701) );
in01f80 newInst_3166 ( .a(newNet_1621), .o(newNet_3166) );
in01f80 newInst_1737 ( .a(newNet_1736), .o(newNet_1737) );
no02f80 g767355 ( .a(n_13492), .b(n_13491), .o(n_13493) );
in01f80 g749295 ( .a(n_30867), .o(n_30868) );
no02f80 g766820 ( .a(n_14300), .b(n_14350), .o(n_14351) );
na02f80 g765079 ( .a(n_15237), .b(FE_OCP_RBN2751_n_15239), .o(n_15313) );
na02f80 g759915 ( .a(n_21051), .b(n_21249), .o(n_21297) );
ms00f80 sin_out_reg_28_ ( .ck(newNet_37), .d(n_43914), .o(sin_out_28) );
in01f80 newInst_3025 ( .a(newNet_3024), .o(newNet_3025) );
na02f80 g746376 ( .a(n_33387), .b(n_33018), .o(n_33434) );
no02f80 g741583 ( .a(n_38645), .b(n_38650), .o(n_38683) );
in01f80 g761887 ( .a(n_18509), .o(n_18510) );
ao12f80 g779134 ( .a(n_1929), .b(n_1928), .c(n_1927), .o(n_2357) );
na02f80 g755739 ( .a(n_24315), .b(n_24041), .o(n_24405) );
no02f80 g776639 ( .a(n_4300), .b(n_3951), .o(n_4374) );
na02f80 g749800 ( .a(n_31222), .b(n_31221), .o(n_31580) );
na02f80 g762228 ( .a(n_18114), .b(n_18079), .o(n_18179) );
in01f80 g772894 ( .a(n_7949), .o(n_7969) );
in01f80 FE_OCP_RBC2398_n_38586 ( .a(n_38586), .o(FE_OCP_RBN2398_n_38586) );
na02f80 g767646 ( .a(n_12771), .b(n_12753), .o(n_12803) );
in01f80 g751507 ( .a(n_28699), .o(n_28700) );
in01f80 FE_OCP_RBC3652_n_10100 ( .a(n_10100), .o(FE_OCP_RBN3652_n_10100) );
in01f80 g757010 ( .a(n_23373), .o(n_23325) );
no02f80 g760742 ( .a(n_20180), .b(n_20198), .o(n_20199) );
oa12f80 g751263 ( .a(n_28778), .b(n_28790), .c(n_28777), .o(n_28829) );
in01f80 g759707 ( .a(n_20638), .o(n_20680) );
no02f80 g755768 ( .a(n_24427), .b(n_24397), .o(n_24484) );
in01f80 g754553 ( .a(n_26901), .o(n_26902) );
oa12f80 g775162 ( .a(n_5727), .b(n_5959), .c(n_5657), .o(n_6025) );
na02f80 g770994 ( .a(n_9667), .b(FE_OFN755_n_44461), .o(n_9820) );
no02f80 g747638 ( .a(n_32170), .b(n_31763), .o(n_32218) );
in01f80 g774042 ( .a(n_6842), .o(n_6843) );
oa12f80 g747771 ( .a(n_33817), .b(n_33571), .c(n_33512), .o(n_33930) );
in01f80 g753293 ( .a(n_27044), .o(n_27045) );
in01f80 g759556 ( .a(n_20957), .o(n_20958) );
in01f80 FE_OCPC977_n_31594 ( .a(FE_OCPN976_n_31594), .o(FE_OCPN977_n_31594) );
na02f80 g741524 ( .a(n_38677), .b(n_38778), .o(n_38704) );
no02f80 FE_RC_3090_0 ( .a(n_45072), .b(n_21384), .o(FE_RN_1364_0) );
na02f80 g749624 ( .a(n_31461), .b(n_31169), .o(n_31582) );
ao12f80 g757222 ( .a(n_23127), .b(n_44219), .c(n_23188), .o(n_23301) );
no02f80 g769339 ( .a(FE_OCP_RBN2002_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_1_), .o(n_11607) );
no02f80 g760965 ( .a(n_19374), .b(n_19498), .o(n_19449) );
in01f80 g751979 ( .a(n_29170), .o(n_29171) );
in01f80 g758521 ( .a(n_22183), .o(n_22184) );
in01f80 newInst_255 ( .a(newNet_38), .o(newNet_255) );
in01f80 FE_RC_3625_0 ( .a(n_45069), .o(FE_RN_1588_0) );
no02f80 g774112 ( .a(n_6734), .b(n_6708), .o(n_6723) );
na02f80 g776972 ( .a(n_4035), .b(n_3958), .o(n_4003) );
in01f80 g740727 ( .a(n_39473), .o(n_39474) );
in01f80 g761478 ( .a(n_19826), .o(n_19827) );
in01f80 g738838 ( .a(n_41340), .o(n_41605) );
in01f80 g754786 ( .a(FE_OCP_RBN2966_n_26231), .o(n_26541) );
in01f80 g768361 ( .a(n_12490), .o(n_12465) );
in01f80 g741033 ( .a(n_39276), .o(n_39277) );
na02f80 g780838 ( .a(n_426), .b(n_405), .o(n_578) );
in01f80 g758236 ( .a(n_23052), .o(n_22950) );
no02f80 g762380 ( .a(FE_OCP_RBN3410_n_45120), .b(n_18420), .o(n_18694) );
ao12f80 g773569 ( .a(n_7457), .b(n_7456), .c(n_7455), .o(n_7683) );
in01f80 g749832 ( .a(n_31254), .o(n_31220) );
in01f80 g762705 ( .a(n_17915), .o(n_17916) );
oa12f80 g737543 ( .a(n_42386), .b(n_42375), .c(n_42367), .o(n_42494) );
na02f80 g773913 ( .a(n_7003), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_7_), .o(n_7081) );
in01f80 newInst_3739 ( .a(newNet_3738), .o(newNet_3739) );
in01f80 g776082 ( .a(n_4878), .o(n_4879) );
in01f80 g774197 ( .a(n_7040), .o(n_7041) );
in01f80 g756415 ( .a(n_24162), .o(n_23825) );
in01f80 FE_OCP_RBC3559_n_8809 ( .a(n_8809), .o(FE_OCP_RBN3559_n_8809) );
na02f80 g777376 ( .a(n_3674), .b(FE_OCPN1042_n_3673), .o(n_3782) );
na02f80 g740069 ( .a(n_40036), .b(n_40071), .o(n_40113) );
oa12f80 g780750 ( .a(n_579), .b(n_584), .c(n_578), .o(n_712) );
ao12f80 g745551 ( .a(n_34357), .b(FE_OCPN1732_n_34369), .c(n_34294), .o(n_34783) );
oa12f80 g768102 ( .a(n_12736), .b(FE_OCP_RBN2219_n_12698), .c(n_12734), .o(n_12816) );
na02f80 g764836 ( .a(n_15888), .b(n_15886), .o(n_15887) );
no02f80 FE_RC_3479_0 ( .a(FE_RN_1495_0), .b(n_40406), .o(n_40422) );
in01f80 FE_OCPC1465_n_13014 ( .a(n_13014), .o(FE_OCPN1465_n_13014) );
oa22f80 g750029 ( .a(FE_OCPN1786_n_30134), .b(n_29059), .c(FE_OCP_RBN3563_n_29857), .d(n_29913), .o(n_30485) );
in01f80 g737949 ( .a(n_42372), .o(n_42293) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_24_ ( .ck(newNet_2935), .d(FE_OCP_RBN3114_n_6379), .o(delay_add_ln22_unr5_stage3_stallmux_q_24_) );
in01f80 g744613 ( .a(n_35375), .o(n_35376) );
na02f80 g750126 ( .a(FE_OCPN1786_n_30134), .b(n_30310), .o(n_30372) );
in01f80 g776476 ( .a(n_4422), .o(n_4423) );
no02f80 g759594 ( .a(n_20756), .b(n_20760), .o(n_20795) );
na02f80 g763648 ( .a(n_16671), .b(n_16714), .o(n_16814) );
in01f80 g773226 ( .a(n_7957), .o(n_7941) );
in01f80 FE_RC_3124_0 ( .a(n_27416), .o(FE_RN_1384_0) );
in01f80 newInst_1844 ( .a(newNet_1843), .o(newNet_1844) );
in01f80 FE_OCPUNCOC1808_n_31435 ( .a(FE_OCPUNCON1807_n_31435), .o(FE_OCPUNCON1808_n_31435) );
na02f80 g739005 ( .a(n_41098), .b(n_40869), .o(n_41161) );
in01f80 g771089 ( .a(n_9718), .o(n_9719) );
in01f80 FE_OCP_RBC3296_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3296_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
in01f80 FE_RC_901_0 ( .a(n_30535), .o(FE_RN_265_0) );
in01f80 g780344 ( .a(n_918), .o(n_958) );
no02f80 g743928 ( .a(n_35786), .b(n_44223), .o(n_35867) );
in01f80 g750917 ( .a(n_28979), .o(n_29018) );
oa12f80 g753801 ( .a(n_26371), .b(n_26370), .c(n_26369), .o(n_26439) );
in01f80 g772217 ( .a(n_8765), .o(n_10105) );
in01f80 g740487 ( .a(n_39787), .o(n_39942) );
in01f80 newInst_3252 ( .a(newNet_3251), .o(newNet_3252) );
ao12f80 g767715 ( .a(n_13371), .b(n_13317), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n_13419) );
in01f80 g773283 ( .a(n_7617), .o(n_7650) );
in01f80 g772972 ( .a(n_7731), .o(n_7749) );
ao22s80 g773891 ( .a(n_6916), .b(n_6852), .c(n_6941), .d(n_6853), .o(n_7022) );
in01f80 g778950 ( .a(n_2305), .o(n_2279) );
in01f80 g763048 ( .a(FE_OCP_DRV_N1548_n_17643), .o(n_17644) );
in01f80 fopt783127 ( .a(n_8875), .o(n_44592) );
ao12f80 g772822 ( .a(n_7301), .b(n_7949), .c(n_7326), .o(n_8042) );
oa22f80 FE_RC_4135_0 ( .a(n_14976), .b(n_15059), .c(n_14975), .d(n_15060), .o(n_15206) );
in01f80 g777318 ( .a(n_5001), .o(n_4972) );
in01f80 g740152 ( .a(n_39918), .o(n_39983) );
no02f80 g771279 ( .a(n_9341), .b(n_9588), .o(n_9720) );
na02f80 g750284 ( .a(n_29779), .b(n_29786), .o(n_29861) );
oa12f80 g747759 ( .a(n_31747), .b(n_32000), .c(n_31554), .o(n_32143) );
na02f80 g773976 ( .a(n_6875), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_5_), .o(n_6993) );
oa12f80 g746759 ( .a(FE_OCP_RBN3385_n_33108), .b(n_33180), .c(delay_add_ln22_unr20_stage8_stallmux_q_21_), .o(n_33189) );
no02f80 g780577 ( .a(n_745), .b(n_744), .o(n_1191) );
in01f80 FE_OCP_RBC2348_n_13702 ( .a(n_13702), .o(FE_OCP_RBN2348_n_13702) );
no02f80 g755945 ( .a(n_24185), .b(n_24210), .o(n_24319) );
in01f80 g779039 ( .a(n_2149), .o(n_2150) );
in01f80 newInst_1100 ( .a(newNet_1099), .o(newNet_1100) );
na02f80 g769928 ( .a(n_11005), .b(n_9798), .o(n_11035) );
no02f80 g756372 ( .a(n_24380), .b(n_24379), .o(n_24381) );
in01f80 g740625 ( .a(n_39638), .o(n_39639) );
in01f80 newInst_1362 ( .a(newNet_1361), .o(newNet_1362) );
in01f80 FE_OCP_RBC3077_FE_OFN807_n_46195 ( .a(FE_OFN807_n_46195), .o(FE_OCP_RBN3077_FE_OFN807_n_46195) );
in01f80 g753394 ( .a(n_27042), .o(n_27043) );
oa22f80 g739675 ( .a(n_40563), .b(n_40306), .c(n_45196), .d(n_45306), .o(n_40593) );
in01f80 g738436 ( .a(n_41906), .o(n_41907) );
in01f80 FE_OCPC3780_n_16440 ( .a(n_16440), .o(FE_OCPN3780_n_16440) );
na02f80 g747341 ( .a(n_32577), .b(n_32437), .o(n_32575) );
in01f80 newInst_2242 ( .a(newNet_2241), .o(newNet_2242) );
in01f80 FE_OCP_RBC1843_n_20910 ( .a(FE_OCP_RBN1842_n_20910), .o(FE_OCP_RBN1843_n_20910) );
oa12f80 g781224 ( .a(beta_22), .b(n_152), .c(beta_31), .o(n_157) );
na02f80 g773575 ( .a(n_7383), .b(n_7373), .o(n_7440) );
oa22f80 g743720 ( .a(n_36372), .b(n_36318), .c(n_36309), .d(n_36319), .o(n_36407) );
in01f80 g747104 ( .a(n_32831), .o(n_32832) );
na02f80 g767306 ( .a(n_13500), .b(n_13452), .o(n_13541) );
oa22f80 g781167 ( .a(n_178), .b(n_131), .c(n_182), .d(n_132), .o(n_470) );
no02f80 g743117 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_12_), .o(n_37147) );
no02f80 FE_RC_1191_0 ( .a(FE_RN_360_0), .b(FE_RN_361_0), .o(FE_RN_362_0) );
no02f80 g754332 ( .a(n_25869), .b(n_25750), .o(n_25894) );
no02f80 g761661 ( .a(n_18940), .b(n_18888), .o(n_18999) );
oa22f80 g743536 ( .a(n_36529), .b(n_36299), .c(n_36530), .d(n_36300), .o(n_36629) );
in01f80 g750334 ( .a(n_29728), .o(n_29729) );
in01f80 newInst_1374 ( .a(newNet_65), .o(newNet_1374) );
in01f80 FE_RC_162_0 ( .a(n_11997), .o(FE_RN_48_0) );
oa22f80 g739914 ( .a(n_40049), .b(n_39919), .c(n_40087), .d(n_39920), .o(n_40198) );
in01f80 FE_OCPC3761_n_2466 ( .a(FE_OCPN3760_n_2466), .o(FE_OCPN3761_n_2466) );
in01f80 g770717 ( .a(n_10415), .o(n_10416) );
no02f80 g773067 ( .a(n_7855), .b(n_7922), .o(n_7951) );
ao12f80 g757667 ( .a(n_22370), .b(n_22463), .c(n_44364), .o(n_22744) );
in01f80 g744506 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_26_), .o(n_36747) );
na02f80 g741338 ( .a(FE_OCP_RBN2546_n_44944), .b(n_38554), .o(n_39130) );
in01f80 fopt783291 ( .a(n_44871), .o(n_44872) );
no02f80 g760097 ( .a(n_20518), .b(n_20124), .o(n_20577) );
in01f80 g754871 ( .a(n_25622), .o(n_25623) );
oa12f80 g779167 ( .a(n_1910), .b(n_2494), .c(n_1909), .o(n_3944) );
no02f80 g771866 ( .a(n_9309), .b(n_9282), .o(n_9880) );
no02f80 g750382 ( .a(n_29695), .b(n_29595), .o(n_29696) );
in01f80 g757613 ( .a(n_24119), .o(n_22767) );
na02f80 g753566 ( .a(n_26775), .b(n_26819), .o(n_26835) );
in01f80 newInst_3138 ( .a(newNet_1792), .o(newNet_3138) );
in01f80 newInst_3679 ( .a(newNet_2128), .o(newNet_3679) );
na02f80 g741198 ( .a(FE_OCP_RBN2639_n_38806), .b(FE_OCP_RBN2351_n_38534), .o(n_38985) );
na02f80 g747004 ( .a(n_32834), .b(n_32736), .o(n_32876) );
in01f80 newInst_1707 ( .a(newNet_1706), .o(newNet_1707) );
no02f80 FE_RC_3080_0 ( .a(FE_OCPN3775_n_14730), .b(n_16333), .o(FE_RN_1358_0) );
ao12f80 g752291 ( .a(n_27864), .b(n_44723), .c(delay_xor_ln22_unr18_stage7_stallmux_q_4_), .o(n_27895) );
in01f80 g770512 ( .a(n_10412), .o(n_10413) );
na02f80 g737197 ( .a(n_42959), .b(n_43012), .o(n_42977) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_15_ ( .ck(newNet_3642), .d(n_46977), .o(delay_add_ln22_unr11_stage5_stallmux_q_15_) );
na02f80 g755871 ( .a(n_25194), .b(n_25081), .o(n_25641) );
no02f80 g777187 ( .a(n_4170), .b(n_4107), .o(n_4561) );
no02f80 g736951 ( .a(FE_OCPN1246_n_43120), .b(n_42926), .o(n_43511) );
no02f80 g779385 ( .a(n_1440), .b(n_1533), .o(n_1541) );
na02f80 g740902 ( .a(n_39262), .b(n_39144), .o(n_39342) );
ao22s80 FE_RC_728_0 ( .a(n_7438), .b(n_8044), .c(n_7437), .d(n_8043), .o(n_8163) );
in01f80 g779555 ( .a(n_1664), .o(n_1665) );
in01f80 FE_OCP_RBC2627_n_14590 ( .a(n_14590), .o(FE_OCP_RBN2627_n_14590) );
no02f80 g747954 ( .a(n_33122), .b(n_33121), .o(n_33123) );
in01f80 g779696 ( .a(delay_xor_ln22_unr3_stage2_stallmux_q_2_), .o(n_1367) );
in01f80 g764499 ( .a(n_16615), .o(n_16630) );
in01f80 g744999 ( .a(n_35824), .o(n_34861) );
no02f80 FE_RC_2948_0 ( .a(FE_RN_1287_0), .b(n_22237), .o(n_22446) );
no02f80 g751152 ( .a(n_30097), .b(n_29817), .o(n_30332) );
na02f80 g765184 ( .a(n_15082), .b(n_15118), .o(n_15235) );
na02f80 g747331 ( .a(n_32688), .b(n_44962), .o(n_32689) );
in01f80 newInst_2964 ( .a(newNet_2249), .o(newNet_2964) );
in01f80 g774246 ( .a(n_6660), .o(n_6661) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_4_ ( .ck(newNet_216), .d(n_46162), .o(delay_xor_ln22_unr6_stage3_stallmux_q_4_) );
in01f80 g748041 ( .a(n_33004), .o(n_32981) );
na02f80 g771538 ( .a(n_9075), .b(FE_OCP_RBN3550_n_44575), .o(n_9101) );
no02f80 g772946 ( .a(n_7799), .b(n_7689), .o(n_7843) );
in01f80 newInst_2545 ( .a(newNet_2544), .o(newNet_2545) );
in01f80 g758635 ( .a(n_22487), .o(n_22488) );
na02f80 g768650 ( .a(n_12101), .b(n_10493), .o(n_12270) );
in01f80 newInst_1722 ( .a(newNet_1556), .o(newNet_1722) );
no02f80 g742141 ( .a(FE_OCPN1239_n_37945), .b(n_37590), .o(n_38167) );
in01f80 g770278 ( .a(n_10618), .o(n_10619) );
no02f80 g781075 ( .a(n_267), .b(n_266), .o(n_268) );
oa12f80 g755369 ( .a(n_22393), .b(n_24875), .c(n_24874), .o(n_24876) );
na02f80 g748371 ( .a(FE_OCPN1052_n_31674), .b(n_31795), .o(n_31897) );
oa12f80 g771568 ( .a(n_9781), .b(n_9332), .c(n_9331), .o(n_9428) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_30_ ( .ck(newNet_1966), .d(n_12197), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_30_) );
in01f80 g777423 ( .a(n_3564), .o(n_3596) );
na02f80 g744279 ( .a(n_44174), .b(n_34924), .o(n_35687) );
in01f80 g747371 ( .a(n_32577), .o(n_32599) );
in01f80 g769563 ( .a(n_11464), .o(n_11465) );
no02f80 g784108 ( .a(n_6866), .b(n_45858), .o(n_45861) );
na02f80 g778613 ( .a(n_2491), .b(n_2140), .o(n_2549) );
no02f80 g762041 ( .a(n_18195), .b(n_18076), .o(n_18204) );
in01f80 g774985 ( .a(n_6233), .o(n_6212) );
na02f80 g781067 ( .a(sin_out_16), .b(FE_OFN3_n_43918), .o(n_332) );
in01f80 g745465 ( .a(n_34653), .o(n_34654) );
na02f80 g741894 ( .a(n_38338), .b(n_37956), .o(n_38190) );
oa12f80 g763136 ( .a(n_17820), .b(n_17819), .c(n_17818), .o(n_17882) );
in01f80 g756237 ( .a(n_24099), .o(n_24100) );
na02f80 g742091 ( .a(FE_OCP_RBN3451_n_37945), .b(n_37551), .o(n_38137) );
in01f80 g766875 ( .a(n_14343), .o(n_14344) );
no02f80 g764686 ( .a(n_46980), .b(n_16111), .o(n_15944) );
ms00f80 delay_xor_ln21_unr3_stage2_stallmux_q_reg_11_ ( .ck(newNet_848), .d(n_1298), .o(delay_xor_ln21_unr3_stage2_stallmux_q_11_) );
na02f80 g778711 ( .a(n_2365), .b(n_2363), .o(n_2389) );
na02f80 g738366 ( .a(n_41709), .b(n_41643), .o(n_41773) );
na02f80 g747988 ( .a(n_33048), .b(n_32563), .o(n_33072) );
na02f80 g750612 ( .a(FE_OCP_RBN2332_n_29380), .b(n_29327), .o(n_29403) );
ao12f80 g769236 ( .a(n_11970), .b(n_45659), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_22_), .o(n_12493) );
in01f80 g753274 ( .a(n_27211), .o(n_27254) );
in01f80 g762016 ( .a(n_18633), .o(n_18705) );
na02f80 g736850 ( .a(n_43460), .b(n_43226), .o(n_43547) );
in01f80 newInst_2458 ( .a(newNet_907), .o(newNet_2458) );
no02f80 FE_RC_2678_0 ( .a(FE_RN_1120_0), .b(n_4166), .o(FE_RN_1121_0) );
no02f80 g761812 ( .a(n_18347), .b(n_18245), .o(n_18411) );
in01f80 FE_RC_4158_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_17_), .o(FE_RN_1810_0) );
na02f80 g769089 ( .a(n_11568), .b(n_11358), .o(n_11599) );
in01f80 g737787 ( .a(n_42208), .o(n_42218) );
na02f80 g761918 ( .a(n_18284), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_21_), .o(n_18401) );
no02f80 g768326 ( .a(n_12490), .b(n_12488), .o(n_12489) );
no02f80 g770173 ( .a(n_10759), .b(n_10601), .o(n_10789) );
oa12f80 g784623 ( .a(FE_OCPN1460_n_37232), .b(n_37377), .c(n_37019), .o(n_46952) );
in01f80 g753716 ( .a(n_27203), .o(n_27198) );
no02f80 g736923 ( .a(FE_OCP_RBN3699_n_43015), .b(n_43021), .o(n_43035) );
in01f80 FE_OCP_RBC3016_n_31117 ( .a(FE_OCP_RBN3014_n_31117), .o(FE_OCP_RBN3016_n_31117) );
in01f80 newInst_2339 ( .a(newNet_1587), .o(newNet_2339) );
na03f80 FE_RC_731_0 ( .a(n_41577), .b(n_41488), .c(n_41479), .o(n_41578) );
in01f80 newInst_1245 ( .a(newNet_1244), .o(newNet_1245) );
ao12f80 g756524 ( .a(n_23969), .b(n_23843), .c(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n_24009) );
no02f80 g772355 ( .a(n_8627), .b(FE_OCP_RBN2480_n_8595), .o(n_8659) );
ao12f80 g743064 ( .a(n_37093), .b(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_27_), .o(n_37140) );
in01f80 newInst_2904 ( .a(newNet_1728), .o(newNet_2904) );
no02f80 g764171 ( .a(n_16582), .b(FE_OCP_RBN1188_n_14823), .o(n_16600) );
na02f80 g750082 ( .a(n_30952), .b(n_30951), .o(n_30953) );
no03m80 g746468 ( .a(n_33380), .b(n_33453), .c(n_33160), .o(n_33381) );
in01f80 FE_OCP_RBC3283_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3283_n_44365) );
in01f80 newInst_2916 ( .a(newNet_2915), .o(newNet_2916) );
na02f80 g746306 ( .a(n_33638), .b(n_33637), .o(n_33639) );
no02f80 g744642 ( .a(n_35326), .b(n_35283), .o(n_35343) );
no02f80 g779324 ( .a(n_1716), .b(n_1450), .o(n_1732) );
oa12f80 g766469 ( .a(n_14495), .b(n_14494), .c(n_14493), .o(n_15786) );
no02f80 g743882 ( .a(n_35826), .b(n_35869), .o(n_35918) );
na02f80 g762268 ( .a(n_18840), .b(n_18611), .o(n_19491) );
na02f80 g746470 ( .a(n_34554), .b(n_34645), .o(n_34617) );
ao12f80 g742723 ( .a(n_37341), .b(n_37340), .c(n_37339), .o(n_38209) );
na02f80 g764630 ( .a(n_16142), .b(n_16140), .o(n_16141) );
na02f80 g764743 ( .a(n_16265), .b(n_16211), .o(n_16450) );
in01f80 g738910 ( .a(n_41298), .o(n_41332) );
in01f80 newInst_3623 ( .a(newNet_3622), .o(newNet_3623) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_7_ ( .ck(newNet_1565), .d(n_26973), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_) );
no02f80 g738275 ( .a(n_41844), .b(n_41620), .o(n_41891) );
na02f80 g775769 ( .a(n_5251), .b(n_5199), .o(n_5310) );
oa12f80 g772714 ( .a(n_8196), .b(n_8195), .c(FE_OCP_RBN2329_n_9003), .o(n_8271) );
ao12f80 g780850 ( .a(n_369), .b(n_420), .c(n_362), .o(n_518) );
ao12f80 g772465 ( .a(n_8306), .b(n_8385), .c(FE_OCP_RBN2301_n_7817), .o(n_8413) );
na02f80 g766230 ( .a(n_14334), .b(n_14191), .o(n_14377) );
oa22f80 g740747 ( .a(n_39448), .b(n_39457), .c(n_39355), .d(n_39458), .o(n_39932) );
in01f80 newInst_2870 ( .a(newNet_927), .o(newNet_2870) );
na02f80 g746599 ( .a(n_34666), .b(n_34739), .o(n_34800) );
na02f80 g771094 ( .a(n_9843), .b(n_9999), .o(n_10132) );
oa22f80 g780150 ( .a(n_1091), .b(FE_OFN760_n_45813), .c(n_1090), .d(n_1203), .o(n_1169) );
in01f80 newInst_683 ( .a(newNet_257), .o(newNet_683) );
na02f80 FE_RC_3561_0 ( .a(n_12914), .b(FE_RN_1546_0), .o(n_13529) );
na02f80 g759420 ( .a(n_21000), .b(n_20999), .o(n_21001) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_19_ ( .ck(newNet_2659), .d(n_22640), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_) );
na02f80 FE_RC_2160_0 ( .a(n_14420), .b(n_15433), .o(FE_RN_765_0) );
in01f80 g744013 ( .a(n_36359), .o(n_36360) );
no02f80 g762888 ( .a(n_17595), .b(n_17444), .o(n_17694) );
no02f80 g740753 ( .a(n_39312), .b(n_39367), .o(n_39445) );
in01f80 fopt783658 ( .a(n_45304), .o(n_45301) );
no02f80 g756806 ( .a(n_23452), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_11_), .o(n_23471) );
in01f80 g779440 ( .a(n_1960), .o(n_1961) );
in01f80 g766303 ( .a(n_45521), .o(n_14384) );
in01f80 newInst_3204 ( .a(newNet_848), .o(newNet_3204) );
in01f80 g736775 ( .a(n_43398), .o(n_43399) );
oa22f80 g775740 ( .a(n_4964), .b(n_4938), .c(n_4965), .d(n_4939), .o(n_5130) );
no02f80 g758214 ( .a(FE_OCP_RBN2044_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_12_), .o(n_23295) );
no02f80 g750813 ( .a(n_30335), .b(n_30256), .o(n_30306) );
no02f80 g770943 ( .a(n_9895), .b(FE_OCPN903_n_44581), .o(n_9899) );
no02f80 g738852 ( .a(n_41319), .b(n_41337), .o(n_41349) );
na02f80 FE_RC_3581_0 ( .a(n_14478), .b(FE_RN_1559_0), .o(FE_RN_1560_0) );
na02f80 g740618 ( .a(n_39542), .b(delay_sub_ln23_0_unr26_stage9_stallmux_q_2_), .o(n_39560) );
in01f80 g739411 ( .a(n_40981), .o(n_40982) );
oa22f80 g753412 ( .a(n_27586), .b(n_26829), .c(n_27587), .d(n_26830), .o(n_27625) );
in01f80 g767360 ( .a(n_13451), .o(n_13452) );
in01f80 FE_OCP_RBC2623_n_3631 ( .a(n_3631), .o(FE_OCP_RBN2623_n_3631) );
no02f80 FE_RC_2693_0 ( .a(FE_RN_1127_0), .b(n_3933), .o(FE_RN_1128_0) );
na02f80 g736945 ( .a(n_43038), .b(n_43181), .o(n_43514) );
in01f80 FE_RC_3311_0 ( .a(n_13913), .o(FE_RN_1457_0) );
in01f80 newInst_3553 ( .a(newNet_3552), .o(newNet_3553) );
no02f80 g746074 ( .a(n_33898), .b(n_33402), .o(n_33922) );
in01f80 FE_OCP_RBC3499_n_8187 ( .a(n_8187), .o(FE_OCP_RBN3499_n_8187) );
in01f80 g748726 ( .a(n_31358), .o(n_31359) );
na02f80 g762382 ( .a(n_45118), .b(n_18526), .o(n_18665) );
ms00f80 sin_out_reg_18_ ( .ck(newNet_67), .d(n_43889), .o(sin_out_18) );
no02f80 g751061 ( .a(n_30380), .b(n_30037), .o(n_30635) );
in01f80 g764215 ( .a(n_16602), .o(n_16579) );
no02f80 g770053 ( .a(n_10907), .b(n_9629), .o(n_11047) );
na02f80 g779178 ( .a(n_1898), .b(delay_add_ln22_unr2_stage2_stallmux_q_10_), .o(n_1935) );
na02f80 g775401 ( .a(n_5712), .b(n_5572), .o(n_5743) );
in01f80 FE_OCP_RBC2461_n_14273 ( .a(n_14273), .o(FE_OCP_RBN2461_n_14273) );
in01f80 g770957 ( .a(n_10129), .o(n_10130) );
in01f80 g754587 ( .a(n_26892), .o(n_26893) );
no02f80 g770740 ( .a(n_10059), .b(n_9933), .o(n_10060) );
oa12f80 FE_RC_3053_0 ( .a(FE_RN_1337_0), .b(FE_RN_1338_0), .c(n_35345), .o(n_35377) );
no02f80 g743584 ( .a(n_37586), .b(n_46200), .o(n_37584) );
na02f80 g759321 ( .a(n_21148), .b(n_21176), .o(n_21344) );
in01f80 g775525 ( .a(n_46999), .o(n_5723) );
in01f80 FE_RC_1218_0 ( .a(n_33898), .o(FE_RN_367_0) );
in01f80 newInst_1641 ( .a(newNet_1640), .o(newNet_1641) );
na02f80 g776038 ( .a(n_5114), .b(n_4497), .o(n_5164) );
no02f80 g765874 ( .a(n_14819), .b(n_14711), .o(n_14883) );
ao12f80 g743416 ( .a(n_37748), .b(n_36775), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37813) );
na02f80 g750398 ( .a(n_29645), .b(n_29644), .o(n_29698) );
in01f80 g772616 ( .a(n_8419), .o(n_8420) );
in01f80 FE_OCPC1448_n_27463 ( .a(FE_OCPN1447_n_27463), .o(FE_OCPN1448_n_27463) );
no02f80 g740669 ( .a(n_39570), .b(n_39589), .o(n_39617) );
no02f80 g739369 ( .a(n_40901), .b(n_40900), .o(n_41243) );
no02f80 g765525 ( .a(n_15874), .b(n_15865), .o(n_15967) );
in01f80 newInst_1508 ( .a(newNet_1507), .o(newNet_1508) );
in01f80 FE_OCP_RBC1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1985_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01f80 g759782 ( .a(n_21695), .o(n_21696) );
in01f80 g758620 ( .a(n_22526), .o(n_22525) );
oa12f80 g741078 ( .a(n_39013), .b(FE_OCP_RBN2689_n_38870), .c(n_38964), .o(n_39455) );
no02f80 g748900 ( .a(n_32393), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .o(n_32508) );
in01f80 FE_OCP_RBC3603_n_8981 ( .a(n_8981), .o(FE_OCP_RBN3603_n_8981) );
na02f80 g751451 ( .a(n_28741), .b(n_28786), .o(n_28802) );
oa12f80 g770971 ( .a(n_10003), .b(n_10045), .c(n_10002), .o(n_10085) );
in01f80 newInst_1572 ( .a(newNet_1571), .o(newNet_1572) );
na02f80 FE_RC_4071_0 ( .a(FE_RN_1772_0), .b(n_36376), .o(n_36410) );
ao12f80 g739021 ( .a(n_41101), .b(n_41100), .c(n_41099), .o(n_41462) );
in01f80 newInst_3032 ( .a(newNet_3031), .o(newNet_3032) );
no02f80 g747424 ( .a(FE_OCP_RBN3331_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_5_), .o(n_32820) );
in01f80 g742774 ( .a(n_37290), .o(n_37608) );
no02f80 g763320 ( .a(n_17220), .b(n_17137), .o(n_17386) );
ao12f80 g778970 ( .a(n_2133), .b(n_2132), .c(n_2131), .o(n_2577) );
oa12f80 g743074 ( .a(n_36987), .b(n_36986), .c(n_36985), .o(n_37800) );
in01f80 FE_OCP_RBC2745_n_47011 ( .a(n_47011), .o(FE_OCP_RBN2745_n_47011) );
in01f80 g761333 ( .a(n_19906), .o(n_19875) );
na02f80 g781034 ( .a(sin_out_3), .b(FE_OFN5_n_43918), .o(n_304) );
in01f80 newInst_16 ( .a(newNet_15), .o(newNet_16) );
no02f80 g753793 ( .a(n_26375), .b(n_26411), .o(n_26531) );
in01f80 newInst_3382 ( .a(newNet_3381), .o(newNet_3382) );
no02f80 g775392 ( .a(n_5417), .b(n_5422), .o(n_5446) );
in01f80 newInst_3127 ( .a(newNet_1873), .o(newNet_3127) );
na02f80 g781300 ( .a(n_7), .b(n_47), .o(n_46) );
na02f80 g774038 ( .a(n_6780), .b(delay_add_ln22_unr5_stage3_stallmux_q_3_), .o(n_6903) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_6_ ( .ck(newNet_1944), .d(n_10389), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_6_) );
no02f80 g770451 ( .a(FE_OCP_RBN2858_n_10399), .b(FE_OCP_RBN3594_n_44561), .o(n_10452) );
oa12f80 g742160 ( .a(n_38253), .b(FE_OCP_RBN2241_n_44881), .c(n_38251), .o(n_38379) );
oa22f80 FE_RC_2403_0 ( .a(n_6598), .b(FE_OCP_RBN3374_n_6745), .c(FE_OCP_RBN2128_n_6745), .d(n_6599), .o(n_6780) );
na02f80 g776478 ( .a(n_4313), .b(n_3297), .o(n_4464) );
in01f80 newInst_1330 ( .a(newNet_1329), .o(newNet_1330) );
ao22s80 FE_RC_1369_0 ( .a(n_43849), .b(n_43602), .c(n_43601), .d(n_43848), .o(n_43879) );
na02f80 g757851 ( .a(n_22389), .b(FE_OCP_RBN3857_FE_RN_779_0), .o(n_22423) );
no02f80 g770034 ( .a(n_10778), .b(FE_OCP_RBN3643_n_44490), .o(n_10860) );
in01f80 newInst_3600 ( .a(newNet_3370), .o(newNet_3600) );
in01f80 FE_OCP_RBC3456_n_33872 ( .a(n_33872), .o(FE_OCP_RBN3456_n_33872) );
in01f80 FE_RC_4041_0 ( .a(FE_RN_1756_0), .o(n_16461) );
in01f80 g746909 ( .a(n_33160), .o(n_33053) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_21_ ( .ck(newNet_2189), .d(n_1152), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_21_) );
in01f80 g778601 ( .a(n_2720), .o(n_2721) );
no02f80 g755172 ( .a(n_24946), .b(n_23628), .o(n_25050) );
no02f80 g745700 ( .a(n_34181), .b(n_34224), .o(n_34225) );
in01f80 FE_OCP_RBC3395_n_28651 ( .a(n_28651), .o(FE_OCP_RBN3395_n_28651) );
in01f80 FE_RC_1914_0 ( .a(n_19170), .o(FE_RN_602_0) );
na02f80 g737595 ( .a(n_42754), .b(n_42801), .o(n_42817) );
na02f80 g750442 ( .a(n_29532), .b(n_29529), .o(n_29634) );
in01f80 g751168 ( .a(n_29977), .o(n_30099) );
in01f80 g739993 ( .a(n_40022), .o(n_40023) );
no02f80 g745767 ( .a(n_34164), .b(n_34036), .o(n_34180) );
oa12f80 g768729 ( .a(n_12178), .b(n_12177), .c(n_12176), .o(n_12283) );
in01f80 newInst_649 ( .a(newNet_648), .o(newNet_649) );
in01f80 newInst_2240 ( .a(newNet_2239), .o(newNet_2240) );
na02f80 FE_RC_3079_0 ( .a(FE_RN_1355_0), .b(FE_RN_1357_0), .o(FE_RN_565_0) );
in01f80 FE_OCP_RBC2239_n_44881 ( .a(FE_OCP_RBN3427_n_44881), .o(FE_OCP_RBN2239_n_44881) );
oa12f80 g752488 ( .a(n_27302), .b(n_27691), .c(n_27401), .o(n_27715) );
in01f80 newInst_2685 ( .a(newNet_2684), .o(newNet_2685) );
no02f80 g777284 ( .a(n_3938), .b(n_4018), .o(n_4170) );
na02f80 g740863 ( .a(n_39310), .b(n_39331), .o(n_39378) );
in01f80 g758221 ( .a(n_22839), .o(n_22809) );
na02f80 g766192 ( .a(n_14380), .b(n_14250), .o(n_14478) );
na02f80 g766935 ( .a(n_14385), .b(n_14294), .o(n_15063) );
no02f80 g767041 ( .a(FE_OCP_RBN2457_n_13765), .b(n_13787), .o(n_13821) );
in01f80 newInst_1435 ( .a(newNet_1434), .o(newNet_1435) );
no02f80 g764449 ( .a(FE_OCP_RBN2919_n_16084), .b(n_14730), .o(n_16162) );
in01f80 fopt783924 ( .a(n_45631), .o(n_45630) );
in01f80 FE_OCP_RBC1915_n_20965 ( .a(FE_OCP_RBN1913_n_20965), .o(FE_OCP_RBN1915_n_20965) );
no02f80 g745708 ( .a(n_34223), .b(FE_OCPN3172_n_34222), .o(n_34272) );
na02f80 g769126 ( .a(n_11481), .b(n_11392), .o(n_11553) );
in01f80 FE_RC_213_0 ( .a(n_12477), .o(FE_RN_69_0) );
in01f80 g769295 ( .a(n_11578), .o(n_11613) );
in01f80 newInst_1661 ( .a(newNet_644), .o(newNet_1661) );
in01f80 FE_OCPC1261_n_20242 ( .a(FE_OCP_RBN1334_n_20249), .o(FE_OCPN1261_n_20242) );
in01f80 g739051 ( .a(n_41173), .o(n_41174) );
in01f80 FE_OCP_RBC3576_n_4528 ( .a(n_4528), .o(FE_OCP_RBN3576_n_4528) );
oa22f80 FE_RC_992_0 ( .a(n_24059), .b(n_27799), .c(n_27796), .d(n_27766), .o(n_27855) );
oa22f80 g780533 ( .a(n_890), .b(FE_OCPN1408_n_672), .c(n_923), .d(n_556), .o(n_1103) );
oa22f80 g763538 ( .a(n_16810), .b(FE_OFN767_n_15670), .c(n_16781), .d(n_16339), .o(n_16873) );
in01f80 g770475 ( .a(n_10404), .o(n_10440) );
no02f80 g744855 ( .a(n_35133), .b(n_35093), .o(n_35167) );
na02f80 g753302 ( .a(n_27207), .b(n_26250), .o(n_27302) );
no02f80 g772201 ( .a(n_8759), .b(n_8200), .o(n_8875) );
in01f80 newInst_2145 ( .a(newNet_1844), .o(newNet_2145) );
in01f80 g743244 ( .a(n_36832), .o(n_36833) );
na02f80 g741042 ( .a(n_39061), .b(n_38922), .o(n_39057) );
in01f80 newInst_3488 ( .a(newNet_248), .o(newNet_3488) );
ao12f80 g746102 ( .a(n_33919), .b(n_33918), .c(n_33917), .o(n_34007) );
in01f80 fopt783212 ( .a(n_12196), .o(n_44766) );
no02f80 g742772 ( .a(n_37387), .b(n_37386), .o(n_37388) );
oa12f80 g739196 ( .a(n_45149), .b(n_40700), .c(delay_add_ln22_unr27_stage10_stallmux_q_23_), .o(n_40794) );
no02f80 g768647 ( .a(FE_OCPN858_n_45697), .b(delay_xor_ln22_unr9_stage4_stallmux_q_15_), .o(n_12319) );
in01f80 g737379 ( .a(n_42812), .o(n_42823) );
na02f80 g760916 ( .a(n_19414), .b(n_18099), .o(n_19427) );
in01f80 g767243 ( .a(n_13597), .o(n_13598) );
no02f80 g748156 ( .a(n_31869), .b(n_32055), .o(n_32101) );
ao12f80 g757072 ( .a(n_23236), .b(n_23235), .c(n_23234), .o(n_23282) );
na02f80 g771808 ( .a(n_8839), .b(n_8849), .o(n_8964) );
no02f80 g765477 ( .a(n_15042), .b(n_15097), .o(n_15149) );
na02f80 g745828 ( .a(n_44102), .b(n_33706), .o(n_34196) );
in01f80 g741612 ( .a(n_38654), .o(n_38628) );
in01f80 g740094 ( .a(n_40289), .o(n_40290) );
in01f80 g736743 ( .a(n_43225), .o(n_43278) );
oa12f80 g750265 ( .a(n_30839), .b(n_30838), .c(n_30837), .o(n_30920) );
in01f80 newInst_623 ( .a(newNet_424), .o(newNet_623) );
no02f80 g767819 ( .a(n_13064), .b(n_12926), .o(n_13736) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_3_ ( .ck(newNet_2715), .d(n_15406), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_3_) );
no02f80 g769683 ( .a(n_11146), .b(n_44511), .o(n_11171) );
no02f80 g776300 ( .a(n_4475), .b(n_4403), .o(n_4535) );
in01f80 g748163 ( .a(n_32134), .o(n_32135) );
ao12f80 g756221 ( .a(n_24677), .b(n_24676), .c(n_24675), .o(n_25251) );
na02f80 g756853 ( .a(n_23404), .b(n_23403), .o(n_23455) );
na02f80 g759330 ( .a(n_21071), .b(n_21120), .o(n_21242) );
in01f80 newInst_267 ( .a(newNet_266), .o(newNet_267) );
no02f80 g744720 ( .a(n_35204), .b(n_35167), .o(n_35205) );
no02f80 g748274 ( .a(FE_OCP_RBN3084_n_31819), .b(n_30738), .o(n_31992) );
ao12f80 g756161 ( .a(n_24846), .b(n_24864), .c(n_24845), .o(n_25258) );
in01f80 newInst_1282 ( .a(newNet_1166), .o(newNet_1282) );
in01f80 g766861 ( .a(n_13661), .o(n_13659) );
in01f80 FE_OCP_RBC2824_n_10068 ( .a(n_10068), .o(FE_OCP_RBN2824_n_10068) );
na02f80 g777640 ( .a(n_3538), .b(n_3499), .o(n_3627) );
ao12f80 g752619 ( .a(n_27269), .b(n_27554), .c(n_27233), .o(n_27604) );
oa12f80 g754883 ( .a(n_25158), .b(n_25187), .c(n_25157), .o(n_26873) );
oa12f80 g763622 ( .a(n_17498), .b(n_17573), .c(delay_sub_ln23_0_unr12_stage5_stallmux_q_29_), .o(n_17665) );
na02f80 g778167 ( .a(n_2843), .b(n_2579), .o(n_2872) );
no02f80 g756786 ( .a(n_23405), .b(n_23264), .o(n_23456) );
na02f80 g757051 ( .a(n_23700), .b(n_23699), .o(n_23808) );
no02f80 g772596 ( .a(n_9304), .b(n_8285), .o(n_8350) );
in01f80 g765802 ( .a(n_15324), .o(n_15325) );
oa12f80 g753540 ( .a(n_26616), .b(n_26701), .c(n_26557), .o(n_26767) );
no02f80 g738456 ( .a(n_41380), .b(n_41388), .o(n_41517) );
ao12f80 g751849 ( .a(n_29129), .b(n_28919), .c(n_29026), .o(n_29746) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_21_ ( .ck(newNet_236), .d(n_46189), .o(delay_xor_ln22_unr6_stage3_stallmux_q_21_) );
oa22f80 g759820 ( .a(n_21714), .b(n_21626), .c(n_21691), .d(n_21719), .o(n_21853) );
na02f80 g778325 ( .a(n_2528), .b(n_2518), .o(n_2519) );
na02f80 g763377 ( .a(FE_OCP_RBN3724_n_16975), .b(FE_OCP_RBN3670_n_46982), .o(n_17185) );
na02f80 g741122 ( .a(n_39200), .b(n_39246), .o(n_39272) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_29_ ( .ck(newNet_2265), .d(n_40577), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_29_) );
na02f80 g744090 ( .a(n_44040), .b(n_35901), .o(n_36192) );
na02f80 g759235 ( .a(n_21891), .b(n_21890), .o(n_21892) );
oa12f80 g784148 ( .a(n_38525), .b(n_38174), .c(n_45890), .o(n_45898) );
na02f80 g762193 ( .a(n_18113), .b(n_17973), .o(n_18170) );
ao12f80 g771793 ( .a(n_8933), .b(n_8932), .c(n_8931), .o(n_9028) );
na02f80 g746553 ( .a(n_34839), .b(n_34756), .o(n_34840) );
no02f80 g750857 ( .a(n_29157), .b(n_29155), .o(n_29158) );
oa12f80 g766007 ( .a(n_15031), .b(n_15030), .c(n_15029), .o(n_15833) );
no02f80 g740886 ( .a(n_39397), .b(n_39429), .o(n_39869) );
oa22f80 g741258 ( .a(FE_OCP_RBN3582_n_44944), .b(n_39040), .c(FE_OCPN942_n_44925), .d(n_38538), .o(n_39451) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_12_ ( .ck(newNet_1543), .d(n_32004), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_12_) );
na02f80 g757984 ( .a(n_22271), .b(n_22131), .o(n_22272) );
na02f80 g767900 ( .a(n_13199), .b(n_13251), .o(n_13769) );
no02f80 g760298 ( .a(n_20264), .b(FE_OCP_RBN1713_FE_RN_664_0), .o(n_20281) );
in01f80 FE_OCPC1763_n_13646 ( .a(n_13646), .o(FE_OCPN1763_n_13646) );
in01f80 fopt782906 ( .a(n_8231), .o(n_44352) );
in01f80 g749500 ( .a(n_30465), .o(n_30464) );
in01f80 g780201 ( .a(delay_sub_ln21_0_unr2_stage2_stallmux_q_19_), .o(n_1141) );
in01f80 g780076 ( .a(n_1215), .o(n_1220) );
no02f80 g757912 ( .a(n_22978), .b(n_22925), .o(n_23437) );
in01f80 g737078 ( .a(n_43383), .o(n_43384) );
na02f80 g758855 ( .a(n_21546), .b(n_21545), .o(n_21547) );
na02f80 g766957 ( .a(n_14296), .b(n_14295), .o(n_14835) );
ao12f80 g769255 ( .a(n_12080), .b(n_45659), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n_12740) );
in01f80 FE_OCP_RBC1906_n_29080 ( .a(FE_OCP_RBN1905_n_29080), .o(FE_OCP_RBN1906_n_29080) );
no02f80 g770920 ( .a(n_9671), .b(n_9675), .o(n_9809) );
no02f80 g743673 ( .a(n_37436), .b(n_37434), .o(n_37477) );
in01f80 FE_OCPC1747_n_23354 ( .a(n_23354), .o(FE_OCPN1747_n_23354) );
in01f80 FE_OCPC3776_n_43019 ( .a(n_43019), .o(FE_OCPN3776_n_43019) );
in01f80 FE_RC_1043_0 ( .a(n_32706), .o(FE_RN_303_0) );
no02f80 g744139 ( .a(n_35739), .b(n_35736), .o(n_35778) );
na02f80 g740206 ( .a(n_39812), .b(n_39534), .o(n_39944) );
na02f80 g755548 ( .a(n_24508), .b(n_24472), .o(n_24761) );
in01f80 g740438 ( .a(n_39792), .o(n_39804) );
no02f80 g750271 ( .a(n_30893), .b(n_30892), .o(n_30894) );
in01f80 newInst_1273 ( .a(newNet_193), .o(newNet_1273) );
oa22f80 FE_RC_1622_0 ( .a(n_17584), .b(n_17811), .c(n_16339), .d(n_17781), .o(n_17855) );
in01f80 g776793 ( .a(n_4329), .o(n_4330) );
in01f80 g743606 ( .a(n_36543), .o(n_36544) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_30_ ( .ck(newNet_1079), .d(FE_OCP_RBN3711_n_46337), .o(n_45224) );
ao12f80 g750911 ( .a(n_29016), .b(n_29015), .c(n_29014), .o(n_29113) );
na02f80 g779205 ( .a(n_1953), .b(n_1952), .o(n_2095) );
no02f80 g752962 ( .a(n_27948), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_25_), .o(n_28107) );
no02f80 g763827 ( .a(n_17462), .b(n_17099), .o(n_17711) );
na02f80 g748265 ( .a(FE_OCP_RBN3735_n_31819), .b(n_30626), .o(n_32051) );
in01f80 newInst_970 ( .a(newNet_969), .o(newNet_970) );
ao22s80 FE_RC_3887_0 ( .a(n_16716), .b(n_16665), .c(n_16735), .d(n_16666), .o(n_16791) );
oa12f80 g742833 ( .a(n_37198), .b(n_37200), .c(n_37197), .o(n_37836) );
na02f80 g738425 ( .a(n_41672), .b(n_41499), .o(n_41673) );
in01f80 g750145 ( .a(n_29954), .o(n_30019) );
in01f80 g761133 ( .a(n_19116), .o(n_19117) );
na02f80 g761694 ( .a(n_19405), .b(n_19406), .o(n_19492) );
oa12f80 g775648 ( .a(n_4966), .b(n_45318), .c(n_4956), .o(n_5206) );
na02f80 g775256 ( .a(n_5857), .b(n_5778), .o(n_5858) );
in01f80 g773988 ( .a(n_7026), .o(n_7027) );
na02f80 g778282 ( .a(n_47026), .b(n_2702), .o(n_2775) );
in01f80 g743613 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n_36470) );
na02f80 g776069 ( .a(n_4947), .b(n_4920), .o(n_5101) );
na02f80 g775036 ( .a(n_5893), .b(n_4875), .o(n_5965) );
na02f80 g751743 ( .a(n_29050), .b(n_29049), .o(n_29051) );
in01f80 g763317 ( .a(n_16884), .o(n_16917) );
na02f80 g758652 ( .a(n_21961), .b(n_22012), .o(n_22032) );
oa22f80 g778749 ( .a(n_2191), .b(n_1499), .c(n_2225), .d(n_1500), .o(n_2807) );
na03f80 FE_RC_3748_0 ( .a(n_40654), .b(n_40653), .c(n_40647), .o(n_40664) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_5_ ( .ck(newNet_905), .d(n_27748), .o(delay_xor_ln21_unr18_stage7_stallmux_q_5_) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_8_ ( .ck(newNet_2433), .d(n_31715), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_8_) );
no02f80 g779030 ( .a(n_2127), .b(delay_add_ln22_unr2_stage2_stallmux_q_16_), .o(n_2141) );
in01f80 g777310 ( .a(n_4106), .o(n_4107) );
ao12f80 g778350 ( .a(n_2366), .b(n_2308), .c(n_2508), .o(n_2575) );
in01f80 g757639 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_20_), .o(n_23658) );
no02f80 g767529 ( .a(n_12976), .b(n_12947), .o(n_13062) );
in01f80 g757321 ( .a(n_23069), .o(n_23070) );
no02f80 g746207 ( .a(n_33664), .b(n_34037), .o(n_33663) );
in01f80 g761500 ( .a(n_18873), .o(n_18874) );
in01f80 g741544 ( .a(n_38707), .o(n_38691) );
ao22s80 FE_RC_550_0 ( .a(FE_OCP_RBN2347_n_29448), .b(n_29690), .c(n_30310), .d(n_29689), .o(n_29753) );
no02f80 g779125 ( .a(n_2445), .b(n_1687), .o(n_1980) );
in01f80 g737305 ( .a(n_46940), .o(n_42936) );
na02f80 g755289 ( .a(n_25580), .b(n_25579), .o(n_25581) );
oa22f80 FE_RC_24_0 ( .a(FE_OFN774_n_46137), .b(n_6436), .c(FE_OFN806_n_46196), .d(n_6476), .o(n_46180) );
na02f80 g766529 ( .a(n_14025), .b(n_13999), .o(n_14114) );
ao12f80 g780051 ( .a(n_816), .b(n_1231), .c(n_1052), .o(n_1242) );
ao12f80 g777409 ( .a(n_2601), .b(n_3386), .c(n_2666), .o(n_3450) );
no02f80 g772789 ( .a(n_8342), .b(FE_OCP_RBN3453_FE_OCPN1240_n_7721), .o(n_8157) );
in01f80 g771498 ( .a(n_9087), .o(n_9088) );
in01f80 g771068 ( .a(n_9743), .o(n_9744) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_9_ ( .ck(newNet_1273), .d(n_1135), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_9_) );
no02f80 FE_RC_637_0 ( .a(FE_RN_198_0), .b(FE_RN_199_0), .o(FE_RN_200_0) );
no02f80 FE_RC_1697_0 ( .a(FE_RN_468_0), .b(FE_RN_469_0), .o(FE_RN_470_0) );
in01f80 newInst_2376 ( .a(newNet_2375), .o(newNet_2376) );
in01f80 g738725 ( .a(n_41499), .o(n_41458) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_11_ ( .ck(newNet_1144), .d(n_10420), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_11_) );
ao22s80 g737233 ( .a(n_42912), .b(n_42800), .c(n_42913), .d(n_42799), .o(n_42968) );
na02f80 g764848 ( .a(n_15439), .b(n_15477), .o(n_15595) );
no02f80 g767551 ( .a(n_12983), .b(n_12975), .o(n_12976) );
na02f80 g743488 ( .a(n_36562), .b(n_36550), .o(n_36626) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_7_ ( .ck(newNet_898), .d(n_27858), .o(delay_xor_ln21_unr18_stage7_stallmux_q_7_) );
no02f80 g749826 ( .a(n_29834), .b(n_29848), .o(n_29905) );
na02f80 g771987 ( .a(n_44464), .b(n_9478), .o(n_9601) );
no02f80 g741550 ( .a(n_38714), .b(n_38713), .o(n_38724) );
ao12f80 g767655 ( .a(n_13069), .b(n_13213), .c(n_11785), .o(n_13214) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_11_ ( .ck(newNet_468), .d(n_27846), .o(delay_xor_ln22_unr18_stage7_stallmux_q_11_) );
na02f80 g777192 ( .a(n_3991), .b(n_4090), .o(n_4419) );
no02f80 g768422 ( .a(n_12428), .b(delay_add_ln22_unr8_stage4_stallmux_q_11_), .o(n_12438) );
na02f80 g776101 ( .a(n_5063), .b(n_5062), .o(n_5116) );
ao12f80 g750175 ( .a(n_29739), .b(n_29736), .c(n_29611), .o(n_29740) );
in01f80 g753281 ( .a(n_27461), .o(n_27411) );
no02f80 g759661 ( .a(n_20383), .b(n_20421), .o(n_20510) );
na02f80 g755703 ( .a(n_24429), .b(n_24520), .o(n_24522) );
na02f80 g766697 ( .a(n_13728), .b(n_13724), .o(n_13780) );
in01f80 newInst_1411 ( .a(newNet_1410), .o(newNet_1411) );
na02f80 g737002 ( .a(FE_OCP_RBN3067_n_43230), .b(n_46936), .o(n_43355) );
in01f80 g752910 ( .a(n_27791), .o(n_27792) );
in01f80 g774229 ( .a(n_6665), .o(n_6666) );
ao12f80 g762898 ( .a(n_17070), .b(n_17494), .c(n_16991), .o(n_17626) );
no02f80 g750369 ( .a(n_30663), .b(n_30635), .o(n_30636) );
na02f80 g754535 ( .a(n_26238), .b(n_26237), .o(n_26239) );
ao12f80 g757172 ( .a(n_23182), .b(n_44995), .c(n_23117), .o(n_23592) );
na02f80 g773765 ( .a(n_7258), .b(n_7036), .o(n_7259) );
no02f80 g746096 ( .a(n_44842), .b(n_33854), .o(n_33957) );
in01f80 g780192 ( .a(n_1143), .o(n_1165) );
oa12f80 g736454 ( .a(n_330), .b(n_43723), .c(FE_OFN2_n_43918), .o(n_43766) );
oa12f80 g762461 ( .a(n_17896), .b(n_18000), .c(n_17849), .o(n_18080) );
in01f80 g762012 ( .a(n_18338), .o(n_18339) );
in01f80 g754591 ( .a(n_26888), .o(n_26889) );
oa12f80 g776678 ( .a(n_3701), .b(n_3786), .c(n_3648), .o(n_3896) );
in01f80 g743021 ( .a(n_36955), .o(n_36956) );
no02f80 g771435 ( .a(n_8974), .b(FE_OCP_RBN3475_n_7886), .o(n_9112) );
na02f80 g756319 ( .a(n_24000), .b(n_23684), .o(n_24042) );
oa22f80 g756153 ( .a(n_24181), .b(n_24100), .c(n_24161), .d(n_24099), .o(n_24270) );
in01f80 newInst_3756 ( .a(newNet_3755), .o(newNet_3756) );
na02f80 g773406 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_), .o(n_7709) );
ao12f80 g750722 ( .a(n_30341), .b(n_30340), .c(n_30339), .o(n_31145) );
na02f80 g776710 ( .a(n_4015), .b(n_3814), .o(n_4068) );
in01f80 g756743 ( .a(n_23482), .o(n_23463) );
na02f80 g763357 ( .a(n_17632), .b(n_17532), .o(n_17633) );
in01f80 g773384 ( .a(n_7609), .o(n_7610) );
in01f80 g737254 ( .a(n_42975), .o(n_42940) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_18_ ( .ck(newNet_2768), .d(n_17128), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_18_) );
no02f80 g754100 ( .a(n_26044), .b(FE_OFN737_n_22641), .o(n_26119) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_0_ ( .ck(newNet_202), .d(n_46380), .o(n_45209) );
na02f80 g757292 ( .a(n_23438), .b(n_22923), .o(n_23469) );
in01f80 newInst_1262 ( .a(newNet_1261), .o(newNet_1262) );
no02f80 g779211 ( .a(n_1924), .b(n_1695), .o(n_1959) );
in01f80 g765341 ( .a(n_15153), .o(n_15154) );
no02f80 g752174 ( .a(n_28592), .b(n_28176), .o(n_28593) );
no02f80 g779614 ( .a(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_15_), .o(n_1797) );
no02f80 g767941 ( .a(n_12711), .b(n_12710), .o(n_12712) );
in01f80 fopt783465 ( .a(n_45073), .o(n_45072) );
no02f80 g748898 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_7_), .o(n_32442) );
in01f80 newInst_1778 ( .a(newNet_1009), .o(newNet_1778) );
in01f80 newInst_471 ( .a(newNet_402), .o(newNet_471) );
in01f80 newInst_346 ( .a(newNet_101), .o(newNet_346) );
na02f80 g773854 ( .a(n_7069), .b(n_7102), .o(n_7108) );
in01f80 fopt783803 ( .a(n_45487), .o(n_45486) );
in01f80 newInst_529 ( .a(newNet_528), .o(newNet_529) );
oa12f80 g739043 ( .a(n_41091), .b(n_41090), .c(n_41089), .o(n_41494) );
oa12f80 g755316 ( .a(n_25473), .b(n_25472), .c(n_25471), .o(n_25685) );
na02f80 g765842 ( .a(n_14865), .b(n_13656), .o(n_14908) );
in01f80 newInst_1711 ( .a(newNet_1710), .o(newNet_1711) );
na02f80 g776040 ( .a(n_4976), .b(n_5026), .o(n_5082) );
na02f80 g770089 ( .a(n_10892), .b(n_10747), .o(n_10929) );
na02f80 g740512 ( .a(n_39748), .b(n_39747), .o(n_39775) );
no02f80 g771898 ( .a(n_9019), .b(n_8959), .o(n_9157) );
na02f80 g784764 ( .a(n_12823), .b(n_12834), .o(n_47250) );
oa12f80 g736501 ( .a(n_313), .b(n_43708), .c(FE_OFN2_n_43918), .o(n_43738) );
na02f80 g750746 ( .a(n_29165), .b(n_28851), .o(n_29279) );
oa12f80 g773513 ( .a(n_7475), .b(n_7474), .c(n_7473), .o(n_7885) );
no02f80 g768012 ( .a(n_12629), .b(n_12498), .o(n_12630) );
na02f80 g770065 ( .a(n_10897), .b(n_10898), .o(n_10958) );
in01f80 newInst_3510 ( .a(newNet_3509), .o(newNet_3510) );
na02f80 g773006 ( .a(n_7796), .b(n_7795), .o(n_7797) );
in01f80 g755423 ( .a(n_26230), .o(n_25605) );
oa12f80 g752022 ( .a(n_28715), .b(n_28714), .c(n_28713), .o(n_29068) );
na02f80 g750423 ( .a(n_29621), .b(n_29520), .o(n_29656) );
na02f80 g752764 ( .a(n_28110), .b(n_28154), .o(n_28155) );
in01f80 g745415 ( .a(n_35679), .o(n_35654) );
in01f80 newInst_2721 ( .a(newNet_963), .o(newNet_2721) );
na02f80 g737620 ( .a(n_42240), .b(n_42237), .o(n_42238) );
na02f80 g740914 ( .a(n_39283), .b(n_39267), .o(n_39309) );
ms00f80 delay_sub_ln21_0_unr11_stage5_stallmux_q_reg_24_ ( .ck(newNet_2741), .d(n_17648), .o(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_) );
na02f80 g771939 ( .a(n_8896), .b(n_8799), .o(n_8960) );
no02f80 FE_RC_4091_0 ( .a(n_21087), .b(n_21080), .o(FE_RN_1789_0) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_17_ ( .ck(newNet_2109), .d(n_6146), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_17_) );
in01f80 g778289 ( .a(n_2725), .o(n_2697) );
in01f80 g745524 ( .a(n_34378), .o(n_34379) );
no02f80 g742997 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_20_), .o(n_37012) );
na02f80 g765093 ( .a(n_15459), .b(n_15458), .o(n_15580) );
ao12f80 g780697 ( .a(n_642), .b(n_646), .c(n_641), .o(n_905) );
na02f80 g768972 ( .a(n_11852), .b(n_11751), .o(n_12193) );
no02f80 g757904 ( .a(n_22235), .b(n_22233), .o(n_22276) );
in01f80 g769250 ( .a(n_11516), .o(n_11517) );
in01f80 FE_OCP_RBC2654_n_9198 ( .a(n_9198), .o(FE_OCP_RBN2654_n_9198) );
no02f80 g748758 ( .a(n_31111), .b(n_27536), .o(n_31201) );
no02f80 g752189 ( .a(FE_OCP_RBN2126_n_44734), .b(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .o(n_28065) );
no02f80 g773388 ( .a(n_7671), .b(n_7638), .o(n_7732) );
na02f80 g767841 ( .a(n_12955), .b(n_12954), .o(n_12997) );
na02f80 g743642 ( .a(n_36441), .b(n_36203), .o(n_36514) );
no02f80 g765352 ( .a(n_15215), .b(n_15250), .o(n_15297) );
na02f80 g767375 ( .a(n_13449), .b(n_13448), .o(n_13450) );
na02f80 g781253 ( .a(n_127), .b(n_91), .o(n_147) );
oa12f80 g776503 ( .a(n_2927), .b(n_4131), .c(n_4073), .o(n_4132) );
na02f80 g748202 ( .a(n_32015), .b(n_32044), .o(n_32122) );
na02f80 g764827 ( .a(n_16178), .b(n_16136), .o(n_16359) );
in01f80 newInst_2746 ( .a(newNet_2745), .o(newNet_2746) );
na02f80 g737900 ( .a(n_42202), .b(n_41867), .o(n_42215) );
na02f80 g741778 ( .a(n_38455), .b(n_38454), .o(n_38456) );
in01f80 g746494 ( .a(n_33291), .o(n_33255) );
oa22f80 g739706 ( .a(n_40475), .b(n_40146), .c(n_40476), .d(n_40145), .o(n_40506) );
oa12f80 g745145 ( .a(n_34659), .b(n_34658), .c(n_34657), .o(n_35667) );
in01f80 g764176 ( .a(n_16532), .o(n_16553) );
na02f80 g776650 ( .a(n_4069), .b(FE_OCP_RBN2626_n_3848), .o(n_4163) );
oa22f80 g784534 ( .a(n_12131), .b(FE_OFN803_n_46285), .c(n_12060), .d(FE_OFN771_n_46337), .o(n_46355) );
na02f80 g768009 ( .a(n_12612), .b(delay_add_ln22_unr8_stage4_stallmux_q_19_), .o(n_12683) );
in01f80 g756024 ( .a(n_25134), .o(n_25194) );
oa12f80 g763181 ( .a(n_17439), .b(n_17438), .c(n_17437), .o(n_18479) );
na02f80 g750655 ( .a(n_31145), .b(n_30393), .o(n_30432) );
in01f80 g771628 ( .a(n_8817), .o(n_8878) );
no02f80 g744235 ( .a(n_46225), .b(n_36859), .o(n_37727) );
na02f80 g777905 ( .a(n_3168), .b(n_3216), .o(n_3220) );
no02f80 g745439 ( .a(n_35541), .b(n_35524), .o(n_36118) );
oa12f80 g751019 ( .a(n_29909), .b(n_29977), .c(n_30086), .o(n_30036) );
ao12f80 g750320 ( .a(n_30691), .b(n_30690), .c(n_30689), .o(n_31288) );
no02f80 FE_RC_1760_0 ( .a(FE_RN_501_0), .b(n_12051), .o(FE_RN_502_0) );
in01f80 newInst_2138 ( .a(newNet_1637), .o(newNet_2138) );
no02f80 g777157 ( .a(n_4685), .b(n_4613), .o(n_5294) );
in01f80 newInst_2943 ( .a(newNet_2942), .o(newNet_2943) );
in01f80 g763699 ( .a(n_17706), .o(n_17707) );
oa22f80 g779021 ( .a(n_45717), .b(n_1498), .c(n_45716), .d(n_1497), .o(n_2432) );
in01f80 g750102 ( .a(n_30051), .o(n_30076) );
in01f80 g774762 ( .a(n_6373), .o(n_6356) );
no02f80 g764129 ( .a(n_16498), .b(n_16535), .o(n_16536) );
no02f80 g764825 ( .a(n_15652), .b(n_14419), .o(n_15653) );
in01f80 FE_OCP_RBC2203_n_18242 ( .a(n_18242), .o(FE_OCP_RBN2203_n_18242) );
na02f80 g766060 ( .a(n_14948), .b(n_14427), .o(n_14949) );
na02f80 g774885 ( .a(n_6182), .b(n_6033), .o(n_6208) );
na02f80 g773612 ( .a(n_7376), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .o(n_7432) );
na02f80 g739904 ( .a(n_40341), .b(n_40084), .o(n_40342) );
in01f80 g775422 ( .a(n_5899), .o(n_5900) );
na02f80 g736546 ( .a(n_43629), .b(n_43091), .o(n_43639) );
in01f80 g761713 ( .a(n_18682), .o(n_18716) );
na02f80 FE_RC_2388_0 ( .a(FE_RN_933_0), .b(FE_RN_934_0), .o(FE_RN_935_0) );
in01f80 g748996 ( .a(FE_OCP_RBN2933_n_31010), .o(n_31034) );
oa12f80 g737284 ( .a(n_42624), .b(n_42842), .c(n_42556), .o(n_42914) );
na02f80 g760876 ( .a(n_19437), .b(n_19436), .o(n_19465) );
no02f80 g779542 ( .a(FE_OCP_RBN3363_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_8_), .o(n_1519) );
na02f80 g775674 ( .a(n_5510), .b(n_5481), .o(n_5482) );
na02f80 g743553 ( .a(n_36474), .b(FE_OCPN1788_n_36034), .o(n_36492) );
in01f80 g771672 ( .a(n_10284), .o(n_10250) );
no02f80 g736872 ( .a(n_43507), .b(n_43538), .o(n_43607) );
in01f80 g748524 ( .a(n_31698), .o(n_31699) );
na02f80 g766225 ( .a(n_14677), .b(n_14676), .o(n_14998) );
in01f80 FE_OCPC1245_n_43120 ( .a(n_43120), .o(FE_OCPN1245_n_43120) );
in01f80 g768209 ( .a(FE_OCP_RBN3420_n_12739), .o(n_13017) );
na02f80 g766549 ( .a(n_13930), .b(FE_OCP_RBN2246_n_13017), .o(n_14000) );
no02f80 g748577 ( .a(n_31383), .b(n_31201), .o(n_31386) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_6_ ( .ck(newNet_1467), .d(n_31671), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_6_) );
no02f80 g756080 ( .a(n_24248), .b(n_23946), .o(n_24264) );
ao12f80 g774236 ( .a(n_7100), .b(n_6806), .c(delay_xor_ln22_unr6_stage3_stallmux_q_17_), .o(n_7190) );
in01f80 FE_OCP_RBC3003_n_10805 ( .a(n_10805), .o(FE_OCP_RBN3003_n_10805) );
in01f80 g773018 ( .a(n_7766), .o(n_7813) );
in01f80 newInst_2650 ( .a(newNet_2649), .o(newNet_2650) );
na02f80 g773587 ( .a(n_7420), .b(n_7224), .o(n_7442) );
ao12f80 g739067 ( .a(n_40851), .b(n_41081), .c(n_40810), .o(n_41135) );
na03f80 g767833 ( .a(n_12860), .b(n_12863), .c(n_12718), .o(n_12861) );
no02f80 g760512 ( .a(n_19891), .b(n_18397), .o(n_19978) );
in01f80 g765027 ( .a(n_15242), .o(n_15286) );
na02f80 g772579 ( .a(n_8359), .b(n_8358), .o(n_8360) );
ao12f80 g753470 ( .a(n_26766), .b(FE_OCP_RBN2983_n_26767), .c(n_26617), .o(n_26786) );
no02f80 g758786 ( .a(n_21509), .b(n_21429), .o(n_21557) );
na02f80 g763066 ( .a(n_17635), .b(n_17634), .o(n_17636) );
in01f80 g740848 ( .a(n_39470), .o(n_39894) );
no02f80 g763290 ( .a(n_16952), .b(n_16808), .o(n_16953) );
na03f80 g755343 ( .a(n_25169), .b(n_25409), .c(n_24999), .o(n_25580) );
in01f80 FE_RC_515_0 ( .a(FE_RN_161_0), .o(n_23199) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_13_ ( .ck(newNet_3557), .d(n_22107), .o(delay_add_ln22_unr14_stage6_stallmux_q_13_) );
no02f80 g753734 ( .a(n_26579), .b(n_26521), .o(n_26614) );
na02f80 g768342 ( .a(n_12554), .b(n_12583), .o(n_12592) );
ao22s80 FE_RC_906_0 ( .a(n_30316), .b(n_30610), .c(n_30317), .d(n_30609), .o(n_30711) );
no02f80 g756563 ( .a(n_23843), .b(delay_add_ln22_unr14_stage6_stallmux_q_29_), .o(n_23969) );
no02f80 g746232 ( .a(n_33707), .b(n_33264), .o(n_33753) );
no02f80 g769014 ( .a(n_11641), .b(FE_OCP_RBN3093_n_11475), .o(n_11723) );
na02f80 g740977 ( .a(n_39139), .b(n_39007), .o(n_39140) );
no02f80 g753806 ( .a(n_26376), .b(FE_OCPN1048_n_24819), .o(n_26377) );
in01f80 newInst_3316 ( .a(newNet_3315), .o(newNet_3316) );
na02f80 g767004 ( .a(n_13765), .b(n_13764), .o(n_13848) );
in01f80 g740171 ( .a(n_40037), .o(n_40119) );
in01f80 FE_OCP_RBC2153_n_32772 ( .a(n_32772), .o(FE_OCP_RBN2153_n_32772) );
in01f80 FE_OCP_RBC2478_n_8599 ( .a(n_8599), .o(FE_OCP_RBN2478_n_8599) );
no02f80 g754925 ( .a(n_25481), .b(FE_OCP_RBN2405_n_24638), .o(n_25673) );
in01f80 g775214 ( .a(n_5813), .o(n_5790) );
na02f80 g745155 ( .a(n_34658), .b(n_34657), .o(n_34659) );
na02f80 g767357 ( .a(n_13390), .b(n_13385), .o(n_13408) );
no02f80 g768348 ( .a(n_12514), .b(n_12066), .o(n_12535) );
oa12f80 g759965 ( .a(FE_OCP_RBN3677_n_21051), .b(n_21294), .c(n_20327), .o(n_21334) );
no02f80 g762146 ( .a(n_18739), .b(n_18576), .o(n_18774) );
oa22f80 g743662 ( .a(n_36408), .b(n_35828), .c(n_36409), .d(n_35829), .o(n_36455) );
ao22s80 FE_RC_4113_0 ( .a(n_23717), .b(n_24094), .c(n_23716), .d(n_24095), .o(n_24175) );
na04m80 g742385 ( .a(n_37754), .b(n_37756), .c(n_37755), .d(FE_OCP_RBN2186_n_37686), .o(n_37772) );
in01f80 FE_OFC3_n_43918 ( .a(FE_OFN0_n_43918), .o(FE_OFN3_n_43918) );
no02f80 g737465 ( .a(n_42650), .b(n_42683), .o(n_42702) );
na02f80 g759219 ( .a(n_20980), .b(n_20944), .o(n_20981) );
no02f80 g744979 ( .a(n_34971), .b(n_34624), .o(n_34976) );
no02f80 g747386 ( .a(n_32436), .b(n_32435), .o(n_32547) );
na02f80 g771678 ( .a(n_9232), .b(n_9330), .o(n_9389) );
ao22s80 FE_RC_4118_0 ( .a(n_27719), .b(n_44759), .c(delay_xor_ln22_unr18_stage7_stallmux_q_0_), .d(FE_OCP_RBN3308_n_44722), .o(n_27773) );
in01f80 newInst_3112 ( .a(newNet_2241), .o(newNet_3112) );
in01f80 FE_OCP_RBC2694_n_15083 ( .a(n_15083), .o(FE_OCP_RBN2694_n_15083) );
no02f80 g776025 ( .a(n_5055), .b(n_4616), .o(n_5140) );
no02f80 g736866 ( .a(n_43356), .b(n_43505), .o(n_43611) );
ao12f80 g759739 ( .a(FE_OCP_RBN3679_n_21051), .b(n_21379), .c(n_21591), .o(n_21409) );
in01f80 FE_OCPC1497_n_26360 ( .a(n_26360), .o(FE_OCPN1497_n_26360) );
na02f80 g745652 ( .a(n_34221), .b(n_34219), .o(n_34287) );
in01f80 newInst_2817 ( .a(newNet_2816), .o(newNet_2817) );
na02f80 g736729 ( .a(n_43149), .b(n_43183), .o(n_43150) );
no02f80 g772980 ( .a(n_7766), .b(n_7680), .o(n_7834) );
oa22f80 FE_RC_1269_0 ( .a(n_38778), .b(n_38545), .c(FE_OCP_RBN2368_n_38545), .d(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38594) );
in01f80 g739959 ( .a(n_40089), .o(n_40046) );
in01f80 g748403 ( .a(n_31553), .o(n_32168) );
no02f80 g755121 ( .a(n_25374), .b(n_24310), .o(n_25375) );
ao12f80 g773803 ( .a(n_7171), .b(n_7180), .c(n_7170), .o(n_7715) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_30_ ( .ck(newNet_2625), .d(n_22874), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_30_) );
na02f80 g743311 ( .a(n_36691), .b(n_36750), .o(n_36724) );
oa12f80 g743052 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_17_), .c(delay_add_ln22_unr23_stage9_stallmux_q_16_), .o(n_37135) );
in01f80 g778786 ( .a(n_2414), .o(n_2438) );
in01f80 g761682 ( .a(n_18938), .o(n_18939) );
no02f80 g745131 ( .a(n_36127), .b(n_36126), .o(n_36179) );
in01f80 g770062 ( .a(n_11061), .o(n_11036) );
ao12f80 g761124 ( .a(n_19237), .b(n_19200), .c(n_19166), .o(n_19300) );
no02f80 g765831 ( .a(n_14823), .b(FE_OCP_RBN2505_n_13896), .o(n_14864) );
na02f80 g738769 ( .a(n_41353), .b(n_41329), .o(n_41355) );
in01f80 g752428 ( .a(n_27868), .o(n_27751) );
in01f80 g771028 ( .a(n_10042), .o(n_10043) );
no02f80 g757864 ( .a(n_22205), .b(n_22003), .o(n_22279) );
in01f80 g740102 ( .a(n_40285), .o(n_40286) );
na02f80 g748135 ( .a(n_32779), .b(n_32586), .o(n_32838) );
in01f80 g740378 ( .a(n_39852), .o(n_40152) );
na02f80 FE_RC_2493_0 ( .a(n_1358), .b(FE_RN_1009_0), .o(FE_RN_1010_0) );
in01f80 g757250 ( .a(n_23208), .o(n_23209) );
na02f80 g774335 ( .a(n_6542), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6543) );
in01f80 g743988 ( .a(n_36367), .o(n_36368) );
na02f80 g764514 ( .a(n_15953), .b(n_16005), .o(n_16169) );
na02f80 FE_RC_821_0 ( .a(FE_RN_246_0), .b(FE_RN_247_0), .o(FE_RN_248_0) );
na02f80 g764193 ( .a(n_16580), .b(n_16515), .o(n_16594) );
no02f80 g778493 ( .a(n_2406), .b(FE_OFN812_n_2405), .o(n_2407) );
no02f80 g739408 ( .a(FE_OCPN898_n_44776), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_8_), .o(n_41052) );
na02f80 g739355 ( .a(n_45153), .b(n_40702), .o(n_40814) );
na02f80 g768690 ( .a(n_12099), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_5_), .o(n_12252) );
in01f80 g780925 ( .a(n_498), .o(n_499) );
na02f80 g746118 ( .a(n_33827), .b(n_33870), .o(n_33900) );
ms00f80 delay_sub_ln23_0_unr5_stage3_stallmux_q_reg_11_ ( .ck(newNet_1260), .d(n_5371), .o(delay_sub_ln23_0_unr5_stage3_stallmux_q_11_) );
in01f80 newInst_1961 ( .a(newNet_1960), .o(newNet_1961) );
ao12f80 g781271 ( .a(n_81), .b(n_46055), .c(beta_14), .o(n_113) );
in01f80 g758519 ( .a(n_21970), .o(n_22002) );
no02f80 g779381 ( .a(n_1547), .b(n_1436), .o(n_1548) );
na02f80 g740750 ( .a(n_39356), .b(n_39035), .o(n_39357) );
in01f80 g748225 ( .a(n_31805), .o(n_31848) );
in01f80 g740588 ( .a(n_39704), .o(n_39705) );
in01f80 g776156 ( .a(n_4927), .o(n_4928) );
ao22s80 FE_RC_1349_0 ( .a(n_15295), .b(n_15655), .c(n_15294), .d(n_15698), .o(n_15861) );
na02f80 g736970 ( .a(FE_OCPN913_n_43022), .b(n_43208), .o(n_43248) );
na02f80 g736832 ( .a(n_43260), .b(n_43125), .o(n_43309) );
in01f80 newInst_3257 ( .a(newNet_3256), .o(newNet_3257) );
no02f80 g772876 ( .a(n_7895), .b(n_7957), .o(n_7958) );
in01f80 newInst_3568 ( .a(newNet_3567), .o(newNet_3568) );
in01f80 newInst_2381 ( .a(newNet_271), .o(newNet_2381) );
na02f80 g769603 ( .a(n_11325), .b(n_11345), .o(n_11353) );
no02f80 g777061 ( .a(n_4973), .b(n_4972), .o(n_4974) );
in01f80 g753012 ( .a(delay_sub_ln23_unr21_stage7_stallmux_q_1_), .o(n_27762) );
no02f80 g778272 ( .a(n_2647), .b(n_3084), .o(n_2650) );
in01f80 g744908 ( .a(n_35029), .o(n_35053) );
no02f80 g776254 ( .a(n_4931), .b(n_4774), .o(n_4935) );
na02f80 g771708 ( .a(n_9180), .b(n_9119), .o(n_9306) );
oa12f80 g736380 ( .a(n_309), .b(n_43784), .c(n_43918), .o(n_43844) );
no02f80 g780086 ( .a(n_1198), .b(n_1191), .o(n_1192) );
oa12f80 g768808 ( .a(n_11684), .b(n_11870), .c(n_11915), .o(n_11954) );
in01f80 g770804 ( .a(n_10179), .o(n_10180) );
no02f80 g768495 ( .a(n_12357), .b(n_12356), .o(n_12358) );
no04s80 g747171 ( .a(n_32706), .b(n_32572), .c(n_32643), .d(FE_OCP_RBN3369_n_32436), .o(n_32740) );
oa22f80 FE_RC_383_0 ( .a(n_966), .b(n_44659), .c(n_897), .d(n_44637), .o(n_1327) );
in01f80 FE_RC_4145_0 ( .a(n_44365), .o(FE_RN_1801_0) );
in01f80 newInst_1493 ( .a(newNet_1492), .o(newNet_1493) );
in01f80 newInst_167 ( .a(newNet_166), .o(newNet_167) );
no02f80 g774977 ( .a(n_6160), .b(n_5299), .o(n_6161) );
oa12f80 g745075 ( .a(n_34817), .b(n_34897), .c(n_34846), .o(n_34930) );
no02f80 g739418 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_10_), .o(n_40725) );
na02f80 FE_RC_2895_0 ( .a(n_39987), .b(FE_RN_1254_0), .o(n_40089) );
oa12f80 g736322 ( .a(n_316), .b(n_43878), .c(FE_OFN1_n_43918), .o(n_43904) );
in01f80 newInst_717 ( .a(newNet_119), .o(newNet_717) );
no02f80 g776841 ( .a(n_4173), .b(n_4058), .o(n_4230) );
na02f80 g744466 ( .a(n_35536), .b(n_35446), .o(n_35522) );
na02f80 g759758 ( .a(n_21299), .b(n_21253), .o(n_21756) );
in01f80 g737633 ( .a(n_42764), .o(n_42765) );
in01f80 g753160 ( .a(n_27544), .o(n_27545) );
no02f80 g744794 ( .a(n_35132), .b(n_47233), .o(n_35173) );
na02f80 FE_RC_4143_0 ( .a(FE_RN_1799_0), .b(n_16829), .o(n_16857) );
na02f80 g753503 ( .a(n_27540), .b(n_26771), .o(n_27559) );
in01f80 newInst_2095 ( .a(newNet_2094), .o(newNet_2095) );
in01f80 newInst_576 ( .a(newNet_575), .o(newNet_576) );
oa12f80 g746690 ( .a(n_34331), .b(n_34330), .c(n_34329), .o(n_34802) );
no02f80 g742990 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_10_), .o(n_36968) );
in01f80 g781113 ( .a(n_241), .o(n_235) );
in01f80 g748038 ( .a(n_31974), .o(n_31975) );
no02f80 g776908 ( .a(FE_OCP_RBN2610_n_3718), .b(n_2913), .o(n_3785) );
in01f80 FE_OCP_DRV_C1589_n_21343 ( .a(n_21343), .o(FE_OCP_DRV_N1589_n_21343) );
in01f80 g744229 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_4_), .o(n_35506) );
no02f80 g784754 ( .a(n_47239), .b(n_7743), .o(n_47240) );
no02f80 g744067 ( .a(n_44223), .b(n_34954), .o(n_35950) );
oa22f80 g739714 ( .a(n_40528), .b(n_40172), .c(n_40529), .d(n_40171), .o(n_40559) );
in01f80 FE_OCP_RBC3836_n_19241 ( .a(FE_OCP_RBN3834_n_19241), .o(FE_OCP_RBN3836_n_19241) );
in01f80 g758111 ( .a(n_22099), .o(n_22131) );
no02f80 g774869 ( .a(n_6196), .b(FE_OCP_RBN2943_n_5454), .o(n_6213) );
in01f80 g746904 ( .a(n_33055), .o(n_33056) );
in01f80 FE_OCP_RBC2799_n_15434 ( .a(n_15434), .o(FE_OCP_RBN2799_n_15434) );
in01f80 g753783 ( .a(n_26493), .o(n_26494) );
no02f80 g750639 ( .a(n_29477), .b(n_29561), .o(n_29351) );
no02f80 g784791 ( .a(n_11556), .b(n_10916), .o(n_47279) );
in01f80 g759923 ( .a(n_21247), .o(n_21248) );
no02f80 g771746 ( .a(n_8879), .b(n_8189), .o(n_8919) );
na02f80 FE_RC_3084_0 ( .a(FE_RN_1360_0), .b(FE_RN_1359_0), .o(FE_RN_1361_0) );
na02f80 g769233 ( .a(FE_OCP_RBN3094_n_11475), .b(n_10369), .o(n_11675) );
na02f80 g777144 ( .a(n_3668), .b(n_3631), .o(n_3669) );
in01f80 g741822 ( .a(n_38930), .o(n_38507) );
na02f80 g740748 ( .a(n_39489), .b(n_39451), .o(n_39518) );
in01f80 g761496 ( .a(n_20220), .o(n_19899) );
in01f80 g741739 ( .a(n_38530), .o(n_38529) );
no02f80 g756904 ( .a(n_23329), .b(n_23288), .o(n_23428) );
na02f80 g762332 ( .a(n_18009), .b(FE_OCP_RBN2149_FE_OCPN861_n_45450), .o(n_18025) );
in01f80 g769214 ( .a(n_11520), .o(n_11518) );
in01f80 newInst_1216 ( .a(newNet_1215), .o(newNet_1216) );
no02f80 g778707 ( .a(n_2414), .b(n_3039), .o(n_2498) );
oa12f80 g778550 ( .a(n_2331), .b(n_2533), .c(n_2330), .o(n_2374) );
in01f80 FE_RC_4252_0 ( .a(n_20295), .o(FE_RN_1871_0) );
no02f80 g766120 ( .a(n_14628), .b(FE_OCP_RBN3529_n_13765), .o(n_14631) );
na02f80 g771358 ( .a(n_8951), .b(FE_OCP_RBN3472_n_7886), .o(n_9016) );
in01f80 g742181 ( .a(n_38301), .o(n_38302) );
na02f80 g768334 ( .a(n_12584), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_14_), .o(n_12618) );
no02f80 g744325 ( .a(n_44174), .b(n_34895), .o(n_36075) );
oa22f80 g749052 ( .a(n_32207), .b(n_31615), .c(n_32206), .d(n_31616), .o(n_32258) );
in01f80 g761343 ( .a(n_19002), .o(n_19003) );
in01f80 g762867 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_26_), .o(n_17722) );
no02f80 g781334 ( .a(n_7), .b(beta_18), .o(n_122) );
na02f80 g743725 ( .a(n_37342), .b(n_36818), .o(n_37362) );
in01f80 g739479 ( .a(n_40713), .o(n_40867) );
na02f80 g776835 ( .a(n_3864), .b(n_3863), .o(n_3913) );
in01f80 g770746 ( .a(n_10116), .o(n_10186) );
na02f80 g740162 ( .a(FE_OCP_RBN3721_n_39913), .b(n_46950), .o(n_40182) );
in01f80 g752111 ( .a(n_28749), .o(n_28782) );
in01f80 newInst_786 ( .a(newNet_174), .o(newNet_786) );
oa12f80 g741741 ( .a(n_38463), .b(n_38462), .c(n_38461), .o(n_38955) );
no02f80 g748281 ( .a(FE_OCP_RBN3735_n_31819), .b(n_46957), .o(n_32046) );
in01f80 newInst_3499 ( .a(newNet_3498), .o(newNet_3499) );
in01f80 g778054 ( .a(n_3056), .o(n_3057) );
in01f80 newInst_729 ( .a(newNet_728), .o(newNet_729) );
oa12f80 FE_RC_2017_0 ( .a(FE_RN_666_0), .b(FE_RN_667_0), .c(n_14021), .o(n_14157) );
na02f80 g736566 ( .a(n_43531), .b(n_43287), .o(n_43638) );
na02f80 g773050 ( .a(n_7717), .b(n_7743), .o(n_7860) );
in01f80 g776667 ( .a(n_47012), .o(n_4289) );
na02f80 g778980 ( .a(n_2188), .b(n_1037), .o(n_2231) );
no02f80 g747790 ( .a(n_33392), .b(n_33438), .o(n_33671) );
ms00f80 cos_out_reg_8_ ( .ck(newNet_3668), .d(n_43738), .o(cos_out_8) );
in01f80 g741333 ( .a(n_38974), .o(n_38975) );
in01f80 newInst_2635 ( .a(newNet_1704), .o(newNet_2635) );
no02f80 g779608 ( .a(n_1518), .b(n_1543), .o(n_1858) );
in01f80 g758203 ( .a(n_22494), .o(n_22495) );
oa22f80 g748615 ( .a(n_31438), .b(n_31419), .c(n_31437), .d(n_31420), .o(n_31514) );
no02f80 FE_RC_2284_0 ( .a(FE_RN_854_0), .b(n_34174), .o(n_34212) );
in01f80 newInst_139 ( .a(newNet_138), .o(newNet_139) );
no02f80 g778586 ( .a(n_2591), .b(n_2651), .o(n_2712) );
no02f80 g773237 ( .a(n_7572), .b(n_7547), .o(n_7596) );
in01f80 g754095 ( .a(n_26120), .o(n_26179) );
no02f80 g754168 ( .a(n_26795), .b(n_26453), .o(n_26818) );
na02f80 FE_RC_2313_0 ( .a(FE_RN_878_0), .b(n_35241), .o(n_35277) );
in01f80 g774571 ( .a(n_6556), .o(n_6789) );
no02f80 g779119 ( .a(n_1955), .b(delay_add_ln22_unr2_stage2_stallmux_q_12_), .o(n_1976) );
no02f80 g771759 ( .a(n_9002), .b(n_44563), .o(n_9169) );
in01f80 g775842 ( .a(n_5028), .o(n_5029) );
in01f80 g770388 ( .a(FE_OCP_RBN2887_n_10570), .o(n_10613) );
no02f80 g759587 ( .a(cordic_combinational_sub_ln23_0_unr20_z_0_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_1_), .o(n_21484) );
no02f80 g768880 ( .a(n_45685), .b(delay_xor_ln21_unr9_stage4_stallmux_q_12_), .o(n_12056) );
na02f80 g768037 ( .a(n_12914), .b(n_12985), .o(n_13075) );
in01f80 newInst_1221 ( .a(newNet_1220), .o(newNet_1221) );
in01f80 g781227 ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_0_), .o(n_167) );
na02f80 g784782 ( .a(n_16241), .b(n_14805), .o(n_47268) );
na02f80 g779640 ( .a(n_1442), .b(n_1441), .o(n_1927) );
no02f80 g742075 ( .a(FE_OCP_RBN3441_n_37945), .b(n_38315), .o(n_38378) );
ao22s80 FE_RC_2627_0 ( .a(n_22772), .b(n_44155), .c(n_22771), .d(n_22677), .o(n_22942) );
ao12f80 g739939 ( .a(n_39860), .b(n_40086), .c(n_39897), .o(n_40231) );
no02f80 g742706 ( .a(n_37396), .b(n_37276), .o(n_37486) );
no02f80 g774316 ( .a(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .b(delay_xor_ln21_unr6_stage3_stallmux_q_9_), .o(n_6772) );
na02f80 g742312 ( .a(n_37822), .b(n_37821), .o(n_37866) );
in01f80 newInst_2489 ( .a(newNet_91), .o(newNet_2489) );
in01f80 newInst_1985 ( .a(newNet_1984), .o(newNet_1985) );
in01f80 g772487 ( .a(n_8525), .o(n_8526) );
na02f80 g781043 ( .a(cos_out_30), .b(FE_OFN1_n_43918), .o(n_308) );
oa12f80 g762808 ( .a(n_17323), .b(n_17659), .c(n_16996), .o(n_17660) );
na02f80 g776985 ( .a(n_3958), .b(n_3957), .o(n_4044) );
in01f80 newInst_1976 ( .a(newNet_1760), .o(newNet_1976) );
no02f80 g740672 ( .a(n_39554), .b(n_39540), .o(n_39992) );
na02f80 g770467 ( .a(n_10559), .b(FE_OCP_RBN3592_n_8902), .o(n_10579) );
no02f80 g742975 ( .a(n_46254), .b(delay_add_ln22_unr23_stage9_stallmux_q_19_), .o(n_37004) );
no02f80 g769037 ( .a(FE_OCP_RBN2113_n_45224), .b(delay_xor_ln21_unr9_stage4_stallmux_q_7_), .o(n_11780) );
na02f80 FE_RC_4054_0 ( .a(FE_RN_1762_0), .b(n_16474), .o(FE_RN_1763_0) );
in01f80 g739885 ( .a(n_40232), .o(n_40233) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_5_ ( .ck(newNet_1799), .d(n_16412), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_5_) );
na02f80 g757217 ( .a(n_23112), .b(n_23111), .o(n_23140) );
in01f80 newInst_3436 ( .a(newNet_1831), .o(newNet_3436) );
na02f80 g780825 ( .a(n_460), .b(n_432), .o(n_602) );
ao22s80 g736540 ( .a(n_43573), .b(n_43146), .c(n_43574), .d(n_43145), .o(n_43653) );
na02f80 g750136 ( .a(n_29815), .b(n_29814), .o(n_29904) );
oa12f80 g766098 ( .a(n_14415), .b(n_14556), .c(n_14555), .o(n_14584) );
oa12f80 g750160 ( .a(FE_OCP_RBN2572_n_29922), .b(n_29260), .c(n_30136), .o(n_30210) );
in01f80 FE_RC_2310_0 ( .a(n_34733), .o(FE_RN_876_0) );
oa22f80 FE_RC_332_0 ( .a(n_22379), .b(n_22618), .c(n_22380), .d(n_22636), .o(n_22806) );
no02f80 g738828 ( .a(n_41327), .b(n_41314), .o(n_41372) );
ao22s80 FE_RC_763_0 ( .a(n_7587), .b(n_8434), .c(n_7586), .d(n_8435), .o(n_8548) );
in01f80 newInst_430 ( .a(newNet_222), .o(newNet_430) );
no02f80 g774825 ( .a(n_6290), .b(n_5754), .o(n_6415) );
ao12f80 g777010 ( .a(n_3592), .b(n_3593), .c(n_3594), .o(n_3600) );
na02f80 g770310 ( .a(n_10720), .b(n_9955), .o(n_10776) );
no02f80 g775582 ( .a(n_5473), .b(n_5512), .o(n_5559) );
na02f80 g744318 ( .a(n_35488), .b(n_35495), .o(n_35489) );
in01f80 g771329 ( .a(n_9111), .o(n_9173) );
no02f80 g751950 ( .a(n_28751), .b(n_28750), .o(n_28752) );
na02f80 g761036 ( .a(n_19315), .b(FE_OCP_DRV_N1554_n_19314), .o(n_19344) );
in01f80 g760699 ( .a(n_19770), .o(n_19771) );
no02f80 g746215 ( .a(n_33820), .b(n_33917), .o(n_33821) );
in01f80 FE_OFC816_n_19885 ( .a(FE_OFN833_n_19885), .o(FE_OFN816_n_19885) );
in01f80 FE_OCP_RBC2204_n_18242 ( .a(n_18242), .o(FE_OCP_RBN2204_n_18242) );
ao22s80 FE_RC_3876_0 ( .a(n_28738), .b(n_29350), .c(n_28737), .d(n_29349), .o(n_29450) );
in01f80 g741155 ( .a(n_38834), .o(n_38835) );
in01f80 g773049 ( .a(n_7860), .o(n_7775) );
na02f80 g739516 ( .a(n_40685), .b(n_40684), .o(n_40709) );
in01f80 g767258 ( .a(n_13497), .o(n_13562) );
in01f80 newInst_774 ( .a(newNet_450), .o(newNet_774) );
ao12f80 g780746 ( .a(n_588), .b(n_590), .c(n_587), .o(n_731) );
na02f80 g780841 ( .a(n_461), .b(n_482), .o(n_624) );
na02f80 g779217 ( .a(n_1863), .b(n_1624), .o(n_1869) );
no02f80 g773173 ( .a(FE_OCPN940_n_7712), .b(n_7700), .o(n_7858) );
in01f80 FE_OCP_RBC3101_n_22504 ( .a(n_22504), .o(FE_OCP_RBN3101_n_22504) );
in01f80 g768699 ( .a(n_12292), .o(n_12225) );
in01f80 newInst_1461 ( .a(newNet_1460), .o(newNet_1461) );
oa12f80 g745162 ( .a(n_36231), .b(n_36230), .c(n_36229), .o(n_36285) );
in01f80 g774355 ( .a(n_6747), .o(n_6748) );
na02f80 g776450 ( .a(n_4708), .b(n_4710), .o(n_4709) );
in01f80 newInst_1663 ( .a(newNet_1662), .o(newNet_1663) );
na02f80 g772412 ( .a(n_8508), .b(n_8561), .o(n_8670) );
in01f80 g762659 ( .a(n_17950), .o(n_17951) );
in01f80 FE_OCP_RBC2748_n_9584 ( .a(n_9584), .o(FE_OCP_RBN2748_n_9584) );
in01f80 g757873 ( .a(n_22359), .o(n_22317) );
in01f80 newInst_468 ( .a(newNet_467), .o(newNet_468) );
in01f80 newInst_2466 ( .a(newNet_1757), .o(newNet_2466) );
na02f80 g776236 ( .a(n_4626), .b(n_4617), .o(n_4723) );
na02f80 g780787 ( .a(n_425), .b(n_370), .o(n_429) );
in01f80 FE_OCPC880_n_31944 ( .a(FE_OCPN879_n_31944), .o(FE_OCPN880_n_31944) );
no02f80 g764363 ( .a(n_16236), .b(n_16233), .o(n_16204) );
no02f80 g773411 ( .a(n_7553), .b(n_6681), .o(n_7572) );
in01f80 g761799 ( .a(n_18678), .o(n_18676) );
oa22f80 g744709 ( .a(n_36479), .b(n_35967), .c(n_36480), .d(n_35966), .o(n_36527) );
in01f80 FE_OCPC1505_n_17680 ( .a(n_17680), .o(FE_OCPN1505_n_17680) );
no02f80 FE_RC_2953_0 ( .a(n_44498), .b(n_10944), .o(FE_RN_1289_0) );
in01f80 g736576 ( .a(n_43567), .o(n_43568) );
na02f80 g772923 ( .a(n_7835), .b(n_7851), .o(n_7852) );
no02f80 g751939 ( .a(n_28149), .b(n_28040), .o(n_28150) );
ao12f80 g742889 ( .a(n_37082), .b(n_37079), .c(n_36466), .o(n_37080) );
na02f80 g743216 ( .a(n_35497), .b(n_36834), .o(n_36887) );
in01f80 g778297 ( .a(n_2973), .o(n_2974) );
in01f80 newInst_1544 ( .a(newNet_1457), .o(newNet_1544) );
no02f80 g741112 ( .a(n_38940), .b(n_38997), .o(n_39048) );
in01f80 g764304 ( .a(n_16432), .o(n_16433) );
in01f80 g750735 ( .a(n_29236), .o(n_29237) );
in01f80 FE_OCP_RBC2392_n_19434 ( .a(FE_OCP_RBN2391_n_19434), .o(FE_OCP_RBN2392_n_19434) );
in01f80 g751692 ( .a(n_28437), .o(n_28447) );
no02f80 FE_RC_4095_0 ( .a(FE_RN_1790_0), .b(FE_OCPN3795_FE_RN_1789_0), .o(n_22326) );
na02f80 g766649 ( .a(n_13818), .b(FE_OCP_RBN2249_n_13017), .o(n_13842) );
no02f80 g773532 ( .a(n_7470), .b(n_7469), .o(n_7471) );
na02f80 g751429 ( .a(n_28458), .b(n_28525), .o(n_28580) );
in01f80 g764099 ( .a(delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(n_17054) );
na02f80 g743090 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_18_), .o(n_37106) );
in01f80 g755796 ( .a(n_24344), .o(n_24345) );
in01f80 FE_OFC798_n_46285 ( .a(n_46285), .o(FE_OFN798_n_46285) );
in01f80 g768718 ( .a(n_12067), .o(n_12143) );
no02f80 g736715 ( .a(n_43346), .b(FE_OCP_RBN3067_n_43230), .o(n_43431) );
in01f80 newInst_43 ( .a(newNet_42), .o(newNet_43) );
ao12f80 g772674 ( .a(n_8481), .b(n_8480), .c(n_8479), .o(n_9321) );
na02f80 g750517 ( .a(n_29474), .b(n_29429), .o(n_29524) );
no02f80 g760772 ( .a(n_20088), .b(n_20087), .o(n_20089) );
no02f80 g745544 ( .a(n_34311), .b(n_34376), .o(n_34438) );
oa12f80 g760890 ( .a(n_19500), .b(n_19499), .c(n_19498), .o(n_21229) );
no02f80 g766052 ( .a(n_14607), .b(n_14505), .o(n_14648) );
in01f80 g754289 ( .a(n_26037), .o(n_26009) );
na02f80 g755560 ( .a(n_24452), .b(n_24477), .o(n_24602) );
na02f80 g751963 ( .a(n_28897), .b(n_28879), .o(n_29006) );
na02f80 g772933 ( .a(n_7897), .b(n_7896), .o(n_7898) );
in01f80 g747361 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_8_), .o(n_32529) );
in01f80 g768644 ( .a(n_12191), .o(n_12192) );
oa12f80 g763957 ( .a(n_16399), .b(n_16532), .c(n_16431), .o(n_16609) );
in01f80 FE_OCP_RBC2804_n_30534 ( .a(n_30534), .o(FE_OCP_RBN2804_n_30534) );
in01f80 newInst_296 ( .a(newNet_92), .o(newNet_296) );
no02f80 g766642 ( .a(n_14308), .b(n_14307), .o(n_14309) );
no02f80 g749711 ( .a(n_31349), .b(n_31291), .o(n_31350) );
no02f80 g747732 ( .a(n_33884), .b(n_33353), .o(n_33933) );
na02f80 g767078 ( .a(n_13597), .b(n_12585), .o(n_13642) );
no02f80 g778983 ( .a(n_2209), .b(n_2208), .o(n_2226) );
in01f80 g775238 ( .a(n_5917), .o(n_5918) );
in01f80 g745221 ( .a(delay_sub_ln23_0_unr28_stage9_stallmux_q_1_), .o(n_35854) );
in01f80 g744871 ( .a(n_35192), .o(n_35249) );
in01f80 g757454 ( .a(n_22869), .o(n_22944) );
no02f80 g756544 ( .a(n_23551), .b(delay_add_ln22_unr14_stage6_stallmux_q_18_), .o(n_23585) );
na02f80 g777913 ( .a(n_3083), .b(n_2968), .o(n_3117) );
in01f80 g759282 ( .a(n_20976), .o(n_20977) );
in01f80 FE_OCPC970_n_14716 ( .a(n_14716), .o(FE_OCPN970_n_14716) );
oa22f80 g752602 ( .a(n_27565), .b(n_27348), .c(n_27566), .d(n_27349), .o(n_27622) );
in01f80 newInst_1578 ( .a(newNet_1577), .o(newNet_1578) );
no02f80 g741505 ( .a(n_38754), .b(n_38741), .o(n_38775) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_29_ ( .ck(newNet_3293), .d(n_32339), .o(delay_add_ln22_unr20_stage8_stallmux_q_29_) );
no02f80 g747162 ( .a(n_32741), .b(n_32740), .o(n_32742) );
in01f80 newInst_1454 ( .a(newNet_573), .o(newNet_1454) );
in01f80 newInst_1945 ( .a(newNet_298), .o(newNet_1945) );
no02f80 g747783 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_13_), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_12_), .o(n_32319) );
na02f80 g746130 ( .a(n_33757), .b(n_33756), .o(n_33778) );
no02f80 g757550 ( .a(n_44084), .b(delay_xor_ln21_unr15_stage6_stallmux_q_9_), .o(n_23322) );
in01f80 g764377 ( .a(n_16321), .o(n_16400) );
in01f80 g778299 ( .a(n_3361), .o(n_2679) );
in01f80 fopt784013 ( .a(n_27582), .o(n_45745) );
no02f80 g774153 ( .a(n_6872), .b(delay_xor_ln21_unr6_stage3_stallmux_q_20_), .o(n_7123) );
ao12f80 g742359 ( .a(n_37704), .b(n_37782), .c(FE_OCP_RBN2187_n_37686), .o(n_37850) );
no02f80 g740221 ( .a(n_39966), .b(FE_OCP_RBN3021_n_39942), .o(n_40034) );
ao12f80 g784614 ( .a(n_42704), .b(n_42687), .c(n_42681), .o(n_46942) );
ms00f80 delay_add_ln22_unr2_stage2_stallmux_q_reg_31_ ( .ck(newNet_3008), .d(n_1118), .o(delay_add_ln22_unr2_stage2_stallmux_q_31_) );
na02f80 g757776 ( .a(n_23092), .b(n_23091), .o(n_23093) );
na02f80 g774158 ( .a(n_6674), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_0_), .o(n_6675) );
ao22s80 g770916 ( .a(n_9890), .b(n_9745), .c(n_9901), .d(FE_OCP_RBN2768_n_9745), .o(n_10138) );
in01f80 newInst_1020 ( .a(newNet_1019), .o(newNet_1020) );
in01f80 g756454 ( .a(n_23997), .o(n_23998) );
in01f80 newInst_1400 ( .a(newNet_1388), .o(newNet_1400) );
in01f80 FE_OCP_RBC2941_FE_RN_473_0 ( .a(FE_RN_473_0), .o(FE_OCP_RBN2941_FE_RN_473_0) );
in01f80 g745053 ( .a(n_35861), .o(n_35906) );
oa22f80 FE_RC_1437_0 ( .a(n_31831), .b(n_32196), .c(n_31832), .d(n_32218), .o(n_32311) );
oa12f80 g753362 ( .a(n_26819), .b(n_26883), .c(n_26774), .o(n_26993) );
no02f80 g746969 ( .a(FE_OCP_RBN2168_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_28_), .o(n_33075) );
in01f80 FE_RC_1943_0 ( .a(n_46415), .o(FE_RN_620_0) );
no02f80 g775150 ( .a(n_5995), .b(n_4972), .o(n_6051) );
na02f80 g745845 ( .a(n_44112), .b(n_34427), .o(n_34428) );
in01f80 FE_RC_1106_0 ( .a(n_44059), .o(FE_RN_331_0) );
no02f80 g772863 ( .a(n_8040), .b(n_8084), .o(n_8141) );
na02f80 FE_RC_751_0 ( .a(delay_xor_ln22_unr18_stage7_stallmux_q_6_), .b(FE_OCPN877_n_44734), .o(FE_RN_234_0) );
no02f80 g776557 ( .a(n_4306), .b(n_4044), .o(n_4421) );
in01f80 newInst_3146 ( .a(newNet_3145), .o(newNet_3146) );
na02f80 g738925 ( .a(n_41190), .b(n_41198), .o(n_41199) );
no02f80 g751542 ( .a(n_28467), .b(delay_add_ln22_unr17_stage7_stallmux_q_19_), .o(n_28571) );
no02f80 g780562 ( .a(n_923), .b(n_660), .o(n_1026) );
ao22s80 g737226 ( .a(n_42900), .b(n_42356), .c(n_42888), .d(n_42355), .o(n_43134) );
in01f80 g777240 ( .a(n_3805), .o(n_3806) );
in01f80 g773186 ( .a(n_7854), .o(n_7855) );
no02f80 g764399 ( .a(n_16093), .b(n_16057), .o(n_16241) );
na02f80 g775707 ( .a(n_5432), .b(n_5413), .o(n_5414) );
in01f80 g744588 ( .a(n_36644), .o(n_36645) );
oa22f80 g777221 ( .a(FE_OCP_RBN2580_n_3734), .b(n_47019), .c(n_3734), .d(n_3439), .o(n_3824) );
in01f80 newInst_809 ( .a(newNet_808), .o(newNet_809) );
in01f80 g775835 ( .a(n_5463), .o(n_5464) );
in01f80 g745773 ( .a(n_34304), .o(n_34305) );
no02f80 g755046 ( .a(n_25415), .b(n_25416), .o(n_25446) );
no02f80 g779530 ( .a(n_1620), .b(n_1619), .o(n_1646) );
in01f80 g747942 ( .a(n_33208), .o(n_33226) );
na02f80 g751476 ( .a(n_28548), .b(n_27654), .o(n_28525) );
oa22f80 FE_RC_614_0 ( .a(n_40921), .b(n_41256), .c(n_40922), .d(FE_OCP_RBN2198_n_41256), .o(n_41312) );
na02f80 g774472 ( .a(n_6586), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_9_), .o(n_6630) );
no02f80 g740050 ( .a(n_40043), .b(n_40015), .o(n_40078) );
no02f80 g739086 ( .a(n_41051), .b(n_40749), .o(n_41064) );
ao22s80 FE_RC_3789_0 ( .a(n_20540), .b(n_20679), .c(n_20500), .d(n_20678), .o(n_20877) );
no02f80 g756303 ( .a(n_23949), .b(n_23612), .o(n_23976) );
ao22s80 g771414 ( .a(n_9083), .b(n_8967), .c(n_9084), .d(n_8966), .o(n_9292) );
oa12f80 g743604 ( .a(n_36102), .b(n_36416), .c(n_36192), .o(n_36444) );
oa12f80 g767590 ( .a(n_12923), .b(n_13100), .c(n_12776), .o(n_13216) );
ao12f80 g780304 ( .a(n_965), .b(n_964), .c(n_1079), .o(n_1050) );
in01f80 g779258 ( .a(n_1838), .o(n_1811) );
oa12f80 g749000 ( .a(n_30946), .b(n_30945), .c(n_30944), .o(n_31008) );
in01f80 newInst_1817 ( .a(newNet_1816), .o(newNet_1817) );
oa12f80 g772369 ( .a(n_7955), .b(n_8519), .c(n_7997), .o(n_8725) );
in01f80 FE_OCP_RBC3667_n_20812 ( .a(n_20812), .o(FE_OCP_RBN3667_n_20812) );
in01f80 g741325 ( .a(n_39120), .o(n_39121) );
no02f80 g754701 ( .a(n_26231), .b(n_26307), .o(n_26232) );
in01f80 g779456 ( .a(n_2145), .o(n_2146) );
in01f80 g754198 ( .a(n_26040), .o(n_26041) );
in01f80 g762128 ( .a(n_18244), .o(n_18245) );
na02f80 g763930 ( .a(n_17101), .b(delay_sub_ln23_0_unr12_stage5_stallmux_q_18_), .o(n_17261) );
ao22s80 g780244 ( .a(n_995), .b(n_798), .c(n_849), .d(n_45809), .o(n_1069) );
in01f80 g768602 ( .a(n_12363), .o(n_12364) );
na02f80 g756248 ( .a(n_24072), .b(n_23665), .o(n_24058) );
in01f80 g755697 ( .a(n_24592), .o(n_24593) );
na02f80 g769979 ( .a(n_11037), .b(n_10925), .o(n_11071) );
in01f80 FE_OCPC1513_FE_OFN738_n_22641 ( .a(FE_OFN738_n_22641), .o(FE_OCPN1513_FE_OFN738_n_22641) );
oa12f80 g752734 ( .a(n_27011), .b(n_27193), .c(n_27192), .o(n_27194) );
in01f80 g771035 ( .a(n_9682), .o(n_9756) );
in01f80 FE_RC_1316_0 ( .a(n_43171), .o(FE_RN_387_0) );
oa22f80 FE_RC_3358_0 ( .a(n_27520), .b(n_27674), .c(n_27519), .d(n_27696), .o(n_27784) );
in01f80 g772510 ( .a(n_8489), .o(n_8490) );
no02f80 g764426 ( .a(n_16052), .b(n_14452), .o(n_16128) );
in01f80 g776575 ( .a(n_4480), .o(n_4481) );
na02f80 g737687 ( .a(n_42367), .b(n_42366), .o(n_42397) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_27_ ( .ck(newNet_2636), .d(n_22914), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_27_) );
na02f80 FE_RC_1569_0 ( .a(FE_RN_446_0), .b(n_28333), .o(n_28405) );
in01f80 g751029 ( .a(n_30166), .o(n_29883) );
ao12f80 g761623 ( .a(n_18818), .b(n_19540), .c(n_18816), .o(n_19611) );
na02f80 g764413 ( .a(n_16172), .b(n_16171), .o(n_16234) );
no02f80 g746964 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_23_), .o(n_32995) );
in01f80 g768352 ( .a(n_12579), .o(n_12580) );
oa12f80 g748101 ( .a(n_32825), .b(n_32824), .c(n_32823), .o(n_33371) );
no02f80 g763270 ( .a(n_17087), .b(FE_OCP_RBN1210_n_16814), .o(n_17283) );
in01f80 FE_OCP_DRV_C1593_n_34494 ( .a(n_34494), .o(FE_OCP_DRV_N1593_n_34494) );
ao12f80 g773659 ( .a(n_7304), .b(n_7303), .c(n_7302), .o(n_7771) );
na02f80 g773708 ( .a(n_7244), .b(delay_add_ln22_unr5_stage3_stallmux_q_16_), .o(n_7268) );
oa12f80 g760382 ( .a(n_20147), .b(FE_OCP_DRV_N1610_n_20146), .c(n_20145), .o(n_20205) );
na02f80 g777309 ( .a(n_4675), .b(n_3470), .o(n_5297) );
in01f80 g737936 ( .a(n_42298), .o(n_42299) );
in01f80 g749666 ( .a(n_30154), .o(n_30121) );
oa22f80 g763869 ( .a(n_16928), .b(n_16310), .c(n_16929), .d(n_16311), .o(n_17058) );
no02f80 g766793 ( .a(n_13661), .b(FE_OCPN860_n_12880), .o(n_13662) );
na02f80 g746035 ( .a(n_33781), .b(n_32986), .o(n_33881) );
in01f80 newInst_496 ( .a(newNet_354), .o(newNet_496) );
in01f80 FE_OCP_RBC2179_FE_RN_526_0 ( .a(FE_RN_526_0), .o(FE_OCP_RBN2179_FE_RN_526_0) );
oa12f80 g750566 ( .a(n_29884), .b(n_30440), .c(n_30332), .o(n_30477) );
no02f80 g771927 ( .a(n_8741), .b(n_8749), .o(n_8835) );
in01f80 g776170 ( .a(n_4843), .o(n_4802) );
oa12f80 g736470 ( .a(n_43245), .b(n_43722), .c(n_43311), .o(n_43754) );
no02f80 g741569 ( .a(n_38660), .b(n_38663), .o(n_38689) );
in01f80 FE_OCPC974_n_46956 ( .a(n_46956), .o(FE_OCPN974_n_46956) );
na02f80 g754225 ( .a(n_26037), .b(n_23466), .o(n_26036) );
in01f80 g773160 ( .a(n_7849), .o(n_7811) );
in01f80 g770704 ( .a(n_10390), .o(n_10391) );
in01f80 newInst_1874 ( .a(newNet_492), .o(newNet_1874) );
oa12f80 g751202 ( .a(n_29334), .b(n_29783), .c(n_29310), .o(n_29824) );
no02f80 g741593 ( .a(n_38622), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38645) );
no02f80 g768588 ( .a(n_12265), .b(n_12264), .o(n_12266) );
in01f80 g754952 ( .a(n_25383), .o(n_25418) );
in01f80 FE_OFC809_n_36594 ( .a(n_36594), .o(FE_OFN809_n_36594) );
no02f80 g751735 ( .a(n_44143), .b(n_28090), .o(n_28346) );
ao12f80 g761625 ( .a(n_18934), .b(n_19494), .c(n_18664), .o(n_19573) );
in01f80 FE_OCP_DRV_C1570_n_29777 ( .a(FE_OCP_DRV_N1569_n_29777), .o(FE_OCP_DRV_N1570_n_29777) );
in01f80 newInst_206 ( .a(newNet_205), .o(newNet_206) );
oa22f80 g747677 ( .a(n_32111), .b(n_31769), .c(n_32112), .d(n_31768), .o(n_32192) );
in01f80 newInst_969 ( .a(newNet_968), .o(newNet_969) );
na02f80 g752930 ( .a(n_27765), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_22_), .o(n_28053) );
no02f80 g744774 ( .a(n_35196), .b(n_35170), .o(n_35262) );
in01f80 g756079 ( .a(n_24264), .o(n_24265) );
in01f80 g778040 ( .a(n_3130), .o(n_3131) );
na02f80 g755127 ( .a(n_25373), .b(n_24529), .o(n_25502) );
in01f80 g738282 ( .a(n_42232), .o(n_41911) );
no02f80 FE_RC_2398_0 ( .a(n_42526), .b(n_42527), .o(FE_RN_944_0) );
no02f80 g737350 ( .a(n_42822), .b(n_42762), .o(n_42841) );
in01f80 g754118 ( .a(n_26142), .o(n_26143) );
in01f80 newInst_650 ( .a(newNet_649), .o(newNet_650) );
in01f80 FE_OCP_RBC3282_n_44365 ( .a(n_44365), .o(FE_OCP_RBN3282_n_44365) );
in01f80 g778507 ( .a(n_3127), .o(n_2393) );
in01f80 g738461 ( .a(n_41764), .o(n_41765) );
in01f80 g778147 ( .a(n_2850), .o(n_2851) );
in01f80 g770057 ( .a(n_11019), .o(n_11037) );
in01f80 g742263 ( .a(n_37861), .o(n_37862) );
no02f80 g748396 ( .a(FE_OCPN1052_n_31674), .b(n_30637), .o(n_31764) );
na02f80 g748011 ( .a(n_33001), .b(n_32455), .o(n_33085) );
oa12f80 g758378 ( .a(n_21871), .b(n_21950), .c(n_21807), .o(n_21999) );
na02f80 g759519 ( .a(n_20821), .b(n_20496), .o(n_20822) );
na02f80 g773686 ( .a(n_7311), .b(n_7788), .o(n_7325) );
ao22s80 g749899 ( .a(n_30922), .b(n_30412), .c(n_30921), .d(n_30413), .o(n_31281) );
na02f80 g773146 ( .a(n_7599), .b(n_7676), .o(n_7677) );
in01f80 g739974 ( .a(n_39959), .o(n_39960) );
no02f80 g763796 ( .a(FE_OCP_RBN3286_n_44365), .b(n_44847), .o(n_16936) );
no02f80 g771119 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_4_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_), .o(n_9993) );
oa22f80 FE_RC_275_0 ( .a(n_14658), .b(n_14714), .c(n_14657), .d(n_14715), .o(n_14814) );
oa12f80 g750933 ( .a(n_28975), .b(n_28974), .c(n_28973), .o(n_29031) );
in01f80 g739439 ( .a(n_40720), .o(n_40812) );
in01f80 g771953 ( .a(n_9480), .o(n_9434) );
in01f80 g769478 ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11707) );
na02f80 g777073 ( .a(n_3824), .b(n_3690), .o(n_3941) );
in01f80 g748197 ( .a(n_32182), .o(n_32183) );
no02f80 g749363 ( .a(n_30602), .b(n_30369), .o(n_30649) );
in01f80 g753081 ( .a(n_27270), .o(n_27271) );
no02f80 g766012 ( .a(n_14613), .b(n_14396), .o(n_14649) );
in01f80 newInst_1044 ( .a(newNet_1043), .o(newNet_1044) );
na02f80 g776199 ( .a(n_4917), .b(n_4826), .o(n_4938) );
in01f80 g743445 ( .a(n_36592), .o(n_36565) );
na02f80 g749886 ( .a(n_30078), .b(FE_OCP_RBN3566_n_29857), .o(n_30176) );
in01f80 g765160 ( .a(n_15308), .o(n_15309) );
in01f80 fopt782967 ( .a(n_44430), .o(n_44429) );
na02f80 g737384 ( .a(n_42783), .b(n_42791), .o(n_43135) );
in01f80 FE_OCP_RBC3024_n_39942 ( .a(FE_OCP_RBN3021_n_39942), .o(FE_OCP_RBN3024_n_39942) );
in01f80 FE_RC_2531_0 ( .a(n_17510), .o(FE_RN_1032_0) );
no02f80 g751357 ( .a(n_29487), .b(n_29047), .o(n_29511) );
no02f80 g767095 ( .a(n_13414), .b(n_12634), .o(n_13459) );
no02f80 g769842 ( .a(n_11178), .b(n_11131), .o(n_11215) );
ao12f80 g747853 ( .a(n_33194), .b(n_33193), .c(n_33192), .o(n_33762) );
na02f80 g775052 ( .a(n_6107), .b(n_6188), .o(n_6171) );
na02f80 g736664 ( .a(n_43164), .b(n_43190), .o(n_43374) );
in01f80 g763354 ( .a(n_17126), .o(n_17127) );
in01f80 newInst_1177 ( .a(newNet_537), .o(newNet_1177) );
in01f80 g774780 ( .a(n_6453), .o(n_6454) );
ao12f80 g743175 ( .a(n_36709), .b(n_36889), .c(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36891) );
na02f80 g740410 ( .a(n_39942), .b(n_39581), .o(n_40030) );
in01f80 newInst_1129 ( .a(newNet_455), .o(newNet_1129) );
in01f80 g776329 ( .a(n_4931), .o(n_4932) );
oa12f80 g752604 ( .a(n_27511), .b(FE_OCP_RBN3736_n_27535), .c(n_27213), .o(n_27582) );
in01f80 g750786 ( .a(n_29193), .o(n_29194) );
na02f80 g762316 ( .a(n_18056), .b(n_18055), .o(n_18114) );
in01f80 g771336 ( .a(n_9354), .o(n_9374) );
in01f80 FE_OCP_RBC3034_n_26842 ( .a(n_26842), .o(FE_OCP_RBN3034_n_26842) );
in01f80 newInst_418 ( .a(newNet_417), .o(newNet_418) );
in01f80 g777782 ( .a(n_3425), .o(n_3426) );
ao12f80 g743140 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_8_), .c(delay_sub_ln21_0_unr23_stage9_stallmux_q_9_), .o(n_37034) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_2_ ( .ck(newNet_3389), .d(n_26477), .o(delay_add_ln22_unr17_stage7_stallmux_q_2_) );
na02f80 g770132 ( .a(n_10787), .b(n_44463), .o(n_10849) );
ao12f80 g756756 ( .a(n_23410), .b(n_23409), .c(n_23408), .o(n_24747) );
in01f80 g743233 ( .a(delay_sub_ln22_unr24_stage9_stallmux_q_2_), .o(n_36834) );
na02f80 g771860 ( .a(n_9692), .b(n_9870), .o(n_10657) );
no02f80 g738391 ( .a(n_41707), .b(n_41671), .o(n_41751) );
in01f80 newInst_3567 ( .a(newNet_2684), .o(newNet_3567) );
no02f80 g776358 ( .a(n_4549), .b(n_4428), .o(n_4496) );
oa12f80 g752597 ( .a(n_27438), .b(n_27568), .c(n_27229), .o(n_27630) );
na02f80 g758882 ( .a(n_21358), .b(n_45070), .o(n_21398) );
in01f80 newInst_1785 ( .a(newNet_1784), .o(newNet_1785) );
oa12f80 g761952 ( .a(n_18136), .b(n_18248), .c(n_18091), .o(n_18269) );
ao12f80 g766810 ( .a(n_13657), .b(n_13705), .c(n_13747), .o(n_13853) );
na02f80 g765931 ( .a(n_14798), .b(FE_OCP_RBN3529_n_13765), .o(n_14799) );
no02f80 g762615 ( .a(n_17971), .b(n_17970), .o(n_17972) );
na02f80 g779041 ( .a(n_2118), .b(n_1879), .o(n_2172) );
na02f80 g769344 ( .a(FE_OCP_RBN2005_delay_sub_ln23_unr9_stage4_stallmux_q_3_), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_5_), .o(n_11544) );
no02f80 g757401 ( .a(n_44084), .b(delay_xor_ln22_unr15_stage6_stallmux_q_7_), .o(n_22972) );
na02f80 g765330 ( .a(n_13785), .b(n_15048), .o(n_15113) );
no02f80 g743363 ( .a(n_36616), .b(n_36634), .o(n_36690) );
in01f80 g757580 ( .a(n_22903), .o(n_22860) );
in01f80 newInst_745 ( .a(newNet_22), .o(newNet_745) );
ao12f80 g757428 ( .a(n_22991), .b(n_22990), .c(n_22989), .o(n_23105) );
in01f80 g755279 ( .a(n_25013), .o(n_25014) );
in01f80 g743705 ( .a(n_36373), .o(n_36374) );
na02f80 g746403 ( .a(n_33388), .b(n_33386), .o(n_33387) );
in01f80 FE_OCP_RBC2169_n_32892 ( .a(FE_OCP_RBN2166_n_32892), .o(FE_OCP_RBN2169_n_32892) );
no02f80 g761271 ( .a(n_19875), .b(n_20014), .o(n_20901) );
in01f80 g745988 ( .a(n_46955), .o(n_34039) );
na02f80 g739291 ( .a(n_40754), .b(n_40848), .o(n_40923) );
na02f80 g753646 ( .a(n_26624), .b(n_26623), .o(n_26625) );
in01f80 newInst_988 ( .a(newNet_668), .o(newNet_988) );
in01f80 newInst_594 ( .a(newNet_203), .o(newNet_594) );
no02f80 g751051 ( .a(n_30097), .b(n_30033), .o(n_30161) );
in01f80 FE_OCP_RBC3574_n_44563 ( .a(FE_OCP_RBN3572_n_44563), .o(FE_OCP_RBN3574_n_44563) );
in01f80 g779153 ( .a(n_1967), .o(n_1999) );
na02f80 g780216 ( .a(n_1114), .b(n_1113), .o(n_1115) );
no02f80 g778477 ( .a(n_2374), .b(n_2449), .o(n_2435) );
in01f80 g762962 ( .a(delay_sub_ln21_0_unr11_stage5_stallmux_q_24_), .o(n_17772) );
in01f80 FE_OCP_RBC2356_n_13858 ( .a(FE_OCP_RBN2355_n_13858), .o(FE_OCP_RBN2356_n_13858) );
in01f80 newInst_3524 ( .a(newNet_3523), .o(newNet_3524) );
no02f80 g765270 ( .a(n_15116), .b(n_14340), .o(n_15119) );
oa12f80 g764551 ( .a(n_16110), .b(n_16154), .c(n_16109), .o(n_16183) );
na02f80 g774865 ( .a(n_6181), .b(n_6032), .o(n_6202) );
na02f80 g780507 ( .a(n_868), .b(n_945), .o(n_987) );
in01f80 g771261 ( .a(n_9552), .o(n_9415) );
no02f80 g761547 ( .a(n_18890), .b(FE_OCP_RBN1329_n_18866), .o(n_18921) );
in01f80 g780128 ( .a(delay_add_ln22_unr2_stage2_stallmux_q_14_), .o(n_1173) );
oa12f80 g773118 ( .a(n_7919), .b(n_8362), .c(n_7908), .o(n_8721) );
oa22f80 g737337 ( .a(n_42823), .b(n_42348), .c(n_42812), .d(n_42349), .o(n_43102) );
na02f80 g765812 ( .a(n_14954), .b(n_14974), .o(n_15066) );
na02f80 g742018 ( .a(n_44035), .b(n_38004), .o(n_38055) );
in01f80 g737679 ( .a(n_42505), .o(n_42486) );
no02f80 g749448 ( .a(n_30510), .b(n_27014), .o(n_30539) );
in01f80 g752234 ( .a(n_27916), .o(n_27917) );
in01f80 newInst_2860 ( .a(newNet_2859), .o(newNet_2860) );
oa22f80 FE_RC_616_0 ( .a(n_40598), .b(n_40578), .c(delay_sub_ln23_0_unr27_stage10_stallmux_z), .d(n_44687), .o(n_40588) );
ao22s80 FE_RC_1150_0 ( .a(n_37087), .b(n_37594), .c(n_37086), .d(n_37593), .o(n_37686) );
na02f80 g775444 ( .a(n_5651), .b(n_4556), .o(n_5712) );
no02f80 g773437 ( .a(n_7553), .b(n_6707), .o(n_7571) );
no02f80 g775276 ( .a(n_5911), .b(n_5677), .o(n_5920) );
na02f80 g747875 ( .a(n_32003), .b(n_31548), .o(n_32032) );
ao12f80 g754497 ( .a(n_26868), .b(n_26740), .c(n_26856), .o(n_26905) );
na02f80 g777602 ( .a(n_3395), .b(n_3387), .o(n_5242) );
oa12f80 g748644 ( .a(n_32590), .b(n_32610), .c(n_32589), .o(n_33362) );
na02f80 g773828 ( .a(n_7093), .b(n_7092), .o(n_7455) );
in01f80 g753387 ( .a(n_27083), .o(n_27098) );
na02f80 g758265 ( .a(n_22208), .b(FE_OFN735_n_22641), .o(n_22951) );
no02f80 g761150 ( .a(n_19078), .b(n_18944), .o(n_19113) );
na02f80 g747084 ( .a(n_32929), .b(n_32908), .o(n_33014) );
in01f80 g777888 ( .a(n_47341), .o(n_3240) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_22_ ( .ck(newNet_3615), .d(n_17594), .o(delay_add_ln22_unr11_stage5_stallmux_q_22_) );
no02f80 g759712 ( .a(FE_OCP_RBN1910_n_20545), .b(n_45066), .o(n_20611) );
no02f80 g754930 ( .a(n_25327), .b(n_24332), .o(n_25328) );
in01f80 g746007 ( .a(n_33923), .o(n_33924) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_26_ ( .ck(newNet_2639), .d(n_22829), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_26_) );
no02f80 g749848 ( .a(n_31040), .b(n_30102), .o(n_31088) );
no02f80 g740632 ( .a(n_39604), .b(n_39611), .o(n_39635) );
in01f80 g737291 ( .a(n_42894), .o(n_42895) );
in01f80 g759049 ( .a(n_21496), .o(n_21533) );
no02f80 g741602 ( .a(n_38583), .b(n_38778), .o(n_38590) );
in01f80 newInst_3583 ( .a(newNet_3582), .o(newNet_3583) );
na02f80 g769364 ( .a(FE_OCPN867_n_45697), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_25_), .o(n_12084) );
na02f80 g740254 ( .a(n_40207), .b(n_39994), .o(n_40311) );
in01f80 g769782 ( .a(n_11240), .o(n_11241) );
in01f80 newInst_2441 ( .a(newNet_2440), .o(newNet_2441) );
in01f80 g767478 ( .a(n_13494), .o(n_13472) );
in01f80 g771480 ( .a(n_9288), .o(n_9289) );
no02f80 g780383 ( .a(n_860), .b(n_1098), .o(n_850) );
na03f80 g761707 ( .a(n_18582), .b(n_19369), .c(n_19400), .o(n_19521) );
na02f80 g766684 ( .a(n_14220), .b(n_14219), .o(n_14221) );
no02f80 g743332 ( .a(n_37828), .b(n_46226), .o(n_37855) );
na02f80 g779079 ( .a(n_2049), .b(n_2018), .o(n_2068) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_21_ ( .ck(newNet_2852), .d(n_11759), .o(delay_add_ln22_unr8_stage4_stallmux_q_21_) );
na02f80 g758801 ( .a(n_21548), .b(n_21506), .o(n_21956) );
ao22s80 g778513 ( .a(n_2516), .b(n_2116), .c(n_2465), .d(n_2117), .o(n_2616) );
in01f80 g738440 ( .a(n_41902), .o(n_41903) );
in01f80 g763327 ( .a(n_17001), .o(n_17002) );
no02f80 g760712 ( .a(n_20182), .b(n_20181), .o(n_20277) );
in01f80 newInst_2478 ( .a(newNet_2477), .o(newNet_2478) );
in01f80 newInst_2224 ( .a(newNet_2223), .o(newNet_2224) );
no02f80 g761253 ( .a(FE_OCP_RBN3827_n_18951), .b(n_19014), .o(n_19015) );
no02f80 g737962 ( .a(n_42169), .b(n_42196), .o(n_42178) );
na02f80 g752723 ( .a(n_27960), .b(n_27813), .o(n_28027) );
no02f80 g765868 ( .a(n_14792), .b(n_14225), .o(n_14827) );
no02f80 g750601 ( .a(n_30440), .b(n_30433), .o(n_30434) );
no02f80 g777305 ( .a(n_3938), .b(n_4136), .o(n_4200) );
in01f80 g737858 ( .a(n_42618), .o(n_42619) );
na02f80 g758199 ( .a(FE_OCPN979_n_21973), .b(n_20724), .o(n_22041) );
na02f80 g749239 ( .a(n_32156), .b(n_31374), .o(n_32174) );
no02f80 g772399 ( .a(n_8573), .b(n_8015), .o(n_8656) );
in01f80 newInst_1717 ( .a(newNet_361), .o(newNet_1717) );
na02f80 g750538 ( .a(n_29453), .b(n_29476), .o(n_29572) );
no02f80 g752041 ( .a(n_28143), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_4_), .o(n_28166) );
na02f80 g771706 ( .a(n_9053), .b(n_9040), .o(n_9234) );
na02f80 g767473 ( .a(n_13226), .b(n_12322), .o(n_13360) );
na02f80 g766413 ( .a(n_14094), .b(n_13132), .o(n_14156) );
no02f80 g741882 ( .a(n_38244), .b(n_38055), .o(n_38286) );
na02f80 g781024 ( .a(cos_out_27), .b(FE_OFN1_n_43918), .o(n_297) );
oa22f80 g739275 ( .a(n_45153), .b(n_40341), .c(n_45155), .d(delay_add_ln22_unr27_stage10_stallmux_q_5_), .o(n_40998) );
in01f80 g779426 ( .a(n_1688), .o(n_1689) );
oa12f80 g761719 ( .a(n_18992), .b(n_19401), .c(n_18964), .o(n_19526) );
no02f80 g775874 ( .a(n_47003), .b(n_47016), .o(n_5372) );
in01f80 g742979 ( .a(n_37006), .o(n_36972) );
no02f80 g748240 ( .a(FE_OCP_RBN3731_n_31819), .b(n_31871), .o(n_32118) );
na02f80 g745459 ( .a(n_34349), .b(FE_OCP_RBN2471_n_34285), .o(n_34463) );
no02f80 g773001 ( .a(n_7965), .b(n_7964), .o(n_7999) );
in01f80 newInst_1352 ( .a(newNet_26), .o(newNet_1352) );
na02f80 g778486 ( .a(n_3058), .b(n_2438), .o(n_2543) );
no02f80 g746794 ( .a(n_33104), .b(n_33098), .o(n_33105) );
oa12f80 g763037 ( .a(n_17233), .b(n_17452), .c(n_17449), .o(n_17487) );
oa12f80 g778996 ( .a(n_2096), .b(n_2106), .c(n_2095), .o(n_2394) );
oa12f80 g747099 ( .a(n_32550), .b(n_32714), .c(n_32554), .o(n_32762) );
na02f80 g756873 ( .a(n_23989), .b(n_23803), .o(n_24034) );
in01f80 g774908 ( .a(n_6228), .o(n_6290) );
in01f80 newInst_2736 ( .a(newNet_2409), .o(newNet_2736) );
no02f80 g775661 ( .a(n_5546), .b(n_5212), .o(n_5591) );
in01f80 g746324 ( .a(n_34350), .o(n_33564) );
na02f80 g744689 ( .a(n_35287), .b(FE_OCPN1794_n_30612), .o(n_35342) );
na03f80 FE_RC_623_0 ( .a(n_39640), .b(n_39743), .c(n_39744), .o(n_39749) );
ao12f80 g755911 ( .a(n_25167), .b(n_25188), .c(n_25122), .o(n_25716) );
no02f80 g746381 ( .a(n_33559), .b(n_33219), .o(n_33607) );
no02f80 g768461 ( .a(n_12457), .b(n_12456), .o(n_12458) );
no02f80 g742791 ( .a(n_37272), .b(n_37126), .o(n_37273) );
in01f80 FE_OCP_RBC2339_n_29385 ( .a(n_29385), .o(FE_OCP_RBN2339_n_29385) );
na03f80 g783816 ( .a(n_15392), .b(n_15353), .c(FE_OCPN1007_n_13962), .o(n_45501) );
na02f80 g760794 ( .a(n_19591), .b(FE_OCP_DRV_N1558_n_19590), .o(n_19623) );
in01f80 newInst_1190 ( .a(newNet_1189), .o(newNet_1190) );
na02f80 g746025 ( .a(n_33964), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33836) );
oa22f80 FE_RC_3231_0 ( .a(n_11745), .b(n_11964), .c(n_11987), .d(n_11746), .o(n_12197) );
no02f80 g754970 ( .a(n_25182), .b(n_25155), .o(n_25212) );
oa12f80 g741344 ( .a(n_38802), .b(n_38843), .c(n_38813), .o(n_38828) );
in01f80 FE_RC_14_0 ( .a(n_2269), .o(FE_RN_4_0) );
in01f80 newInst_434 ( .a(newNet_433), .o(newNet_434) );
na02f80 g768962 ( .a(n_11786), .b(n_11774), .o(n_11788) );
in01f80 g777287 ( .a(n_3815), .o(n_3816) );
no02f80 g737249 ( .a(n_42899), .b(n_42764), .o(n_42931) );
no02f80 g771405 ( .a(n_9609), .b(n_9563), .o(n_9688) );
in01f80 FE_OCP_DRV_C3160_n_31303 ( .a(FE_OCP_DRV_N3159_n_31303), .o(FE_OCP_DRV_N3160_n_31303) );
no02f80 g766291 ( .a(n_14534), .b(n_14568), .o(n_14677) );
na02f80 g745519 ( .a(n_34650), .b(n_34648), .o(n_34649) );
na02f80 g754155 ( .a(n_26947), .b(n_26452), .o(n_26834) );
na02f80 g757493 ( .a(n_22899), .b(n_22898), .o(n_22933) );
na02f80 g739562 ( .a(n_40616), .b(delay_add_ln22_unr27_stage10_stallmux_q_0_), .o(n_40739) );
in01f80 g764130 ( .a(n_16699), .o(n_16681) );
no02f80 g755707 ( .a(n_25171), .b(n_25083), .o(n_25223) );
na02f80 g770176 ( .a(n_10727), .b(n_10664), .o(n_10875) );
na02f80 g758991 ( .a(n_21537), .b(FE_OCPN1524_n_45072), .o(n_21644) );
no02f80 g762409 ( .a(FE_OCP_RBN3409_n_45120), .b(n_18487), .o(n_18584) );
in01f80 g747353 ( .a(n_33544), .o(n_32728) );
no02f80 g778627 ( .a(n_2620), .b(FE_OCP_RBN2294_n_2438), .o(n_2617) );
no02f80 g771996 ( .a(n_44498), .b(n_8810), .o(n_10081) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_7_ ( .ck(newNet_1279), .d(n_854), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_7_) );
no02f80 g743221 ( .a(n_36803), .b(n_36847), .o(n_36876) );
no02f80 g773698 ( .a(n_7244), .b(delay_add_ln22_unr5_stage3_stallmux_q_16_), .o(n_7291) );
no02f80 g746091 ( .a(n_33779), .b(n_33829), .o(n_33878) );
ao12f80 g747965 ( .a(n_32776), .b(n_33048), .c(n_32452), .o(n_33131) );
no03m80 g756251 ( .a(n_24047), .b(n_24671), .c(n_24063), .o(n_24816) );
ao12f80 g772032 ( .a(n_8773), .b(n_8824), .c(n_8772), .o(n_10078) );
in01f80 FE_RC_3075_0 ( .a(n_27125), .o(FE_RN_1354_0) );
na02f80 g765585 ( .a(n_15044), .b(n_15045), .o(n_15136) );
no02f80 g776103 ( .a(n_4906), .b(n_4905), .o(n_4975) );
oa22f80 g744716 ( .a(FE_OCP_RBN2665_n_35207), .b(n_30614), .c(n_35207), .d(n_30633), .o(n_35231) );
no02f80 FE_RC_1741_0 ( .a(n_11707), .b(FE_RN_487_0), .o(FE_RN_488_0) );
oa12f80 g768241 ( .a(n_12676), .b(n_12675), .c(n_12674), .o(n_12729) );
na02f80 g741530 ( .a(n_38732), .b(n_38731), .o(n_38740) );
in01f80 g777943 ( .a(n_3159), .o(n_3160) );
no02f80 g746861 ( .a(n_34081), .b(n_33951), .o(n_34132) );
in01f80 g743326 ( .a(n_36722), .o(n_36723) );
na02f80 g768468 ( .a(n_12424), .b(n_12385), .o(n_12587) );
oa12f80 g770535 ( .a(n_10432), .b(n_10431), .c(n_10430), .o(n_10496) );
in01f80 FE_RC_1234_0 ( .a(FE_RN_371_0), .o(n_6554) );
in01f80 g759503 ( .a(delay_sub_ln23_0_unr16_stage6_stallmux_q_3_), .o(n_22658) );
in01f80 g780032 ( .a(n_1255), .o(n_1256) );
in01f80 FE_OCPC1765_n_33447 ( .a(n_33447), .o(FE_OCPN1765_n_33447) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_21_ ( .ck(newNet_1511), .d(n_32258), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_21_) );
in01f80 g780435 ( .a(n_822), .o(n_886) );
no02f80 g760003 ( .a(n_20667), .b(n_20778), .o(n_20786) );
in01f80 FE_OCPC1416_FE_OCP_RBN1362_n_20504 ( .a(FE_OCPN1415_FE_OCP_RBN1362_n_20504), .o(FE_OCPN1416_FE_OCP_RBN1362_n_20504) );
no02f80 g746582 ( .a(n_34473), .b(n_34580), .o(n_34615) );
no02f80 g757561 ( .a(n_23298), .b(n_23296), .o(n_23297) );
in01f80 newInst_3576 ( .a(newNet_3575), .o(newNet_3576) );
ao12f80 g749758 ( .a(n_30072), .b(n_30119), .c(n_29869), .o(n_30203) );
in01f80 g740695 ( .a(n_39477), .o(n_39478) );
in01f80 FE_OCP_RBC2657_FE_RN_1288_0 ( .a(FE_RN_1288_0), .o(FE_OCP_RBN2657_FE_RN_1288_0) );
in01f80 newInst_1356 ( .a(newNet_1355), .o(newNet_1356) );
na02f80 g743146 ( .a(n_36982), .b(n_37084), .o(n_37236) );
oa22f80 g742825 ( .a(n_37286), .b(n_37177), .c(n_37266), .d(n_37176), .o(n_37392) );
oa12f80 g755665 ( .a(n_24551), .b(n_24550), .c(n_24549), .o(n_26296) );
oa22f80 g768442 ( .a(n_12366), .b(n_12287), .c(n_12412), .d(n_12288), .o(n_12436) );
no02f80 g749302 ( .a(n_30646), .b(n_30708), .o(n_30709) );
oa12f80 g736300 ( .a(n_297), .b(n_43879), .c(FE_OFN1_n_43918), .o(n_43909) );
oa22f80 g764228 ( .a(n_16742), .b(n_16253), .c(n_16743), .d(n_16254), .o(n_16815) );
in01f80 g769961 ( .a(n_10998), .o(n_11024) );
oa12f80 g774275 ( .a(n_6390), .b(n_6514), .c(n_6371), .o(n_6572) );
na02f80 g743036 ( .a(n_37150), .b(n_37041), .o(n_37180) );
na02f80 g760435 ( .a(n_20033), .b(n_19968), .o(n_20030) );
na02f80 g765822 ( .a(n_15289), .b(n_14561), .o(n_15362) );
na02f80 g764450 ( .a(n_16615), .b(n_15965), .o(n_16674) );
in01f80 FE_OCPC1731_n_34369 ( .a(n_34369), .o(FE_OCPN1731_n_34369) );
in01f80 g775826 ( .a(n_5136), .o(n_5137) );
in01f80 g772530 ( .a(n_8642), .o(n_8591) );
na02f80 g744679 ( .a(n_35253), .b(n_35200), .o(n_35272) );
in01f80 g743388 ( .a(n_36733), .o(n_36734) );
oa12f80 g778212 ( .a(n_2673), .b(n_2674), .c(n_2438), .o(n_2774) );
na02f80 g770961 ( .a(n_9625), .b(n_9670), .o(n_9723) );
no02f80 g751996 ( .a(n_28919), .b(n_28937), .o(n_29004) );
na02f80 g778135 ( .a(n_2899), .b(n_2898), .o(n_2977) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_21_ ( .ck(newNet_1315), .d(n_1249), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_21_) );
no02f80 g777765 ( .a(n_3454), .b(n_3453), .o(n_3455) );
na02f80 g762321 ( .a(n_18160), .b(n_18159), .o(n_18213) );
no02f80 g741509 ( .a(n_38709), .b(n_38656), .o(n_38710) );
no02f80 FE_RC_3495_0 ( .a(n_30526), .b(n_30527), .o(FE_RN_1507_0) );
ao12f80 g760841 ( .a(n_20058), .b(n_20057), .c(n_19731), .o(n_20088) );
na02f80 g740177 ( .a(FE_OCP_RBN3715_n_39913), .b(n_39947), .o(n_40036) );
in01f80 FE_OCP_RBC2536_n_3645 ( .a(n_3645), .o(FE_OCP_RBN2536_n_3645) );
in01f80 newInst_2502 ( .a(newNet_671), .o(newNet_2502) );
in01f80 g775775 ( .a(n_5606), .o(n_5607) );
na02f80 g737216 ( .a(n_42907), .b(n_42797), .o(n_42920) );
in01f80 g774896 ( .a(n_6311), .o(n_6312) );
no02f80 g739101 ( .a(n_41058), .b(n_41057), .o(n_41059) );
na02f80 g780142 ( .a(n_948), .b(n_1006), .o(n_1085) );
in01f80 g779589 ( .a(n_1972), .o(n_1973) );
na02f80 g762363 ( .a(n_45002), .b(n_18531), .o(n_18616) );
na02f80 g760494 ( .a(n_19974), .b(n_18230), .o(n_20027) );
na02f80 g766995 ( .a(n_13737), .b(n_13736), .o(n_13738) );
ao22s80 g756516 ( .a(n_23821), .b(n_23773), .c(n_23783), .d(delay_sub_ln21_0_unr14_stage6_stallmux_q_23_), .o(n_23844) );
ao22s80 g768322 ( .a(n_12519), .b(n_12329), .c(n_12482), .d(n_12328), .o(n_13625) );
na02f80 g777161 ( .a(n_4675), .b(n_5166), .o(n_5328) );
na02f80 g751899 ( .a(n_28991), .b(n_28907), .o(n_29456) );
no02f80 g756203 ( .a(FE_OCP_RBN2278_n_24173), .b(FE_OCPN3164_n_24117), .o(n_24221) );
in01f80 newInst_3654 ( .a(newNet_3653), .o(newNet_3654) );
ao12f80 g749100 ( .a(n_30833), .b(n_30862), .c(n_30832), .o(n_30945) );
in01f80 fopt783560 ( .a(n_45149), .o(n_45153) );
in01f80 FE_OCPC1048_n_24819 ( .a(FE_OCPN1047_n_24819), .o(FE_OCPN1048_n_24819) );
in01f80 g762891 ( .a(n_17630), .o(n_17628) );
oa12f80 g776260 ( .a(n_4696), .b(n_4697), .c(n_4695), .o(n_4775) );
in01f80 newInst_2827 ( .a(newNet_815), .o(newNet_2827) );
na02f80 FE_RC_2703_0 ( .a(FE_RN_1132_0), .b(FE_RN_1135_0), .o(FE_RN_1136_0) );
no02f80 g745443 ( .a(FE_OCP_RBN2988_n_35539), .b(n_35108), .o(n_36126) );
no02f80 g746484 ( .a(n_34777), .b(n_34741), .o(n_34844) );
ao12f80 g744447 ( .a(n_35385), .b(n_35460), .c(n_35410), .o(n_35495) );
oa12f80 g773120 ( .a(n_7840), .b(n_8362), .c(n_7296), .o(n_8644) );
in01f80 g777296 ( .a(n_4864), .o(n_4817) );
in01f80 newInst_2438 ( .a(newNet_163), .o(newNet_2438) );
na02f80 g737888 ( .a(n_42201), .b(n_42131), .o(n_42417) );
oa12f80 g751498 ( .a(n_28286), .b(n_28372), .c(n_28294), .o(n_28477) );
no02f80 g746271 ( .a(n_44814), .b(FE_OCP_RBN1681_n_33491), .o(n_33618) );
no02f80 g773142 ( .a(FE_OCP_RBN2228_n_7598), .b(n_7630), .o(n_7667) );
in01f80 g769688 ( .a(n_11333), .o(n_11342) );
in01f80 g758552 ( .a(FE_OCP_RBN1848_n_22068), .o(n_22187) );
in01f80 g740665 ( .a(n_40011), .o(n_39627) );
in01f80 g774501 ( .a(n_6591), .o(n_6592) );
no02f80 g751384 ( .a(n_28535), .b(n_28512), .o(n_28513) );
in01f80 g756762 ( .a(n_23443), .o(n_23444) );
oa12f80 g742788 ( .a(n_37315), .b(n_37314), .c(n_37313), .o(n_37393) );
no02f80 g767829 ( .a(n_12796), .b(n_12942), .o(n_12797) );
in01f80 FE_OCP_RBC3634_n_47260 ( .a(n_47260), .o(FE_OCP_RBN3634_n_47260) );
na02f80 g736364 ( .a(n_43814), .b(n_43440), .o(n_43809) );
in01f80 g751555 ( .a(n_28522), .o(n_28574) );
in01f80 g771393 ( .a(n_9527), .o(n_9528) );
no02f80 g746958 ( .a(n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_), .o(n_33246) );
na02f80 g769254 ( .a(FE_OCP_RBN3093_n_11475), .b(FE_OCP_RBN2999_n_11004), .o(n_11649) );
in01f80 g749007 ( .a(n_31177), .o(n_31261) );
no02f80 g747112 ( .a(n_33995), .b(n_33994), .o(n_33996) );
na02f80 g771751 ( .a(n_10159), .b(n_10158), .o(n_10160) );
na02f80 g743383 ( .a(n_36565), .b(delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36617) );
in01f80 g748349 ( .a(n_31858), .o(n_31859) );
in01f80 g742304 ( .a(n_37842), .o(n_37843) );
na02f80 g748145 ( .a(n_31805), .b(n_32139), .o(n_32163) );
na02f80 g770180 ( .a(n_10710), .b(n_10756), .o(n_10845) );
no02f80 g767058 ( .a(FE_OCP_RBN2459_n_13765), .b(n_13934), .o(n_13970) );
ao12f80 g738122 ( .a(n_41809), .b(n_42030), .c(n_41830), .o(n_42041) );
no02f80 g771618 ( .a(n_10341), .b(n_10284), .o(n_10343) );
na02f80 g774366 ( .a(n_6510), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(n_6656) );
in01f80 newInst_1034 ( .a(newNet_905), .o(newNet_1034) );
no02f80 g766187 ( .a(n_14998), .b(n_14733), .o(n_14735) );
in01f80 newInst_2312 ( .a(newNet_2311), .o(newNet_2312) );
no02f80 g754966 ( .a(n_25155), .b(n_25154), .o(n_25156) );
ao22s80 FE_RC_2940_0 ( .a(n_11809), .b(n_12024), .c(n_11808), .d(n_11989), .o(n_12067) );
in01f80 g769655 ( .a(n_11364), .o(n_11365) );
in01f80 FE_OCP_RBC3136_n_32380 ( .a(n_32380), .o(FE_OCP_RBN3136_n_32380) );
in01f80 g763768 ( .a(n_17266), .o(n_17306) );
in01f80 g757727 ( .a(n_22709), .o(n_22666) );
in01f80 g736992 ( .a(n_43266), .o(n_43247) );
oa12f80 g762755 ( .a(n_17766), .b(n_17846), .c(n_17718), .o(n_17928) );
no02f80 g767705 ( .a(n_12870), .b(n_12869), .o(n_12898) );
na02f80 g777627 ( .a(n_3372), .b(n_3211), .o(n_3387) );
na02f80 g761761 ( .a(n_18678), .b(FE_OFN778_n_17093), .o(n_18679) );
in01f80 fopt783672 ( .a(n_5272), .o(n_45323) );
ao12f80 g762796 ( .a(n_17758), .b(n_45450), .c(delay_xor_ln21_unr12_stage5_stallmux_q_9_), .o(n_17778) );
na02f80 g774755 ( .a(n_6355), .b(n_6262), .o(n_6485) );
in01f80 FE_OCPC1771_n_26801 ( .a(n_26801), .o(FE_OCPN1771_n_26801) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_27_ ( .ck(newNet_3130), .d(n_40567), .o(delay_add_ln22_unr27_stage10_stallmux_q_27_) );
no02f80 g772999 ( .a(n_7724), .b(n_7458), .o(n_7774) );
na02f80 g749916 ( .a(n_30120), .b(n_30011), .o(n_30147) );
in01f80 g777812 ( .a(n_3388), .o(n_3406) );
in01f80 FE_OCP_RBC1674_n_36492 ( .a(n_36492), .o(FE_OCP_RBN1674_n_36492) );
na02f80 g745526 ( .a(n_34405), .b(n_34320), .o(n_34630) );
ao12f80 g772030 ( .a(n_8085), .b(n_8824), .c(n_8031), .o(n_8868) );
in01f80 FE_OCPC930_n_44083 ( .a(FE_OCPN929_n_44083), .o(FE_OCPN930_n_44083) );
oa12f80 g757175 ( .a(n_23528), .b(n_23527), .c(n_23526), .o(n_23670) );
ao12f80 g746503 ( .a(n_34528), .b(n_34527), .c(n_35542), .o(n_35559) );
ao12f80 g745141 ( .a(n_34710), .b(n_34725), .c(n_34709), .o(n_34765) );
in01f80 FE_OCPC1499_n_26125 ( .a(n_26125), .o(FE_OCPN1499_n_26125) );
na02f80 FE_RC_2863_0 ( .a(FE_RN_1233_0), .b(n_14329), .o(n_14447) );
no02f80 g751600 ( .a(FE_OCP_RBN3403_n_28597), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_26_), .o(n_28736) );
in01f80 FE_OCP_RBC2346_n_29448 ( .a(n_29448), .o(FE_OCP_RBN2346_n_29448) );
no02f80 g742598 ( .a(n_37569), .b(n_37453), .o(n_37570) );
in01f80 g757365 ( .a(n_23416), .o(n_23417) );
no02f80 g740589 ( .a(n_39671), .b(n_39664), .o(n_39704) );
na02f80 FE_RC_669_0 ( .a(FE_RN_212_0), .b(n_36945), .o(n_37144) );
na02f80 g752559 ( .a(n_27598), .b(n_27427), .o(n_27599) );
in01f80 g757868 ( .a(n_22389), .o(n_22421) );
na02f80 g763019 ( .a(n_17937), .b(n_17430), .o(n_17981) );
oa12f80 g779374 ( .a(n_1840), .b(n_1466), .c(FE_OCPN946_n_1780), .o(n_1841) );
oa12f80 g738210 ( .a(n_41674), .b(n_41946), .c(n_41510), .o(n_41969) );
in01f80 FE_RC_3111_0 ( .a(n_31652), .o(FE_RN_1377_0) );
ao12f80 g775057 ( .a(n_5969), .b(n_6038), .c(n_5963), .o(n_6054) );
no02f80 g773434 ( .a(n_7608), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_29_), .o(n_7638) );
no02f80 g779226 ( .a(n_1818), .b(n_1817), .o(n_1819) );
in01f80 g781268 ( .a(n_89), .o(n_90) );
na02f80 g766632 ( .a(n_13917), .b(n_13888), .o(n_14059) );
na02f80 g760625 ( .a(n_19808), .b(FE_OFN815_n_19807), .o(n_19835) );
no02f80 FE_RC_3688_0 ( .a(FE_RN_1619_0), .b(FE_RN_1620_0), .o(FE_RN_1621_0) );
na02f80 g775508 ( .a(n_5375), .b(n_5301), .o(n_5433) );
no02f80 FE_RC_2204_0 ( .a(FE_RN_792_0), .b(n_26338), .o(n_26506) );
na02f80 g751577 ( .a(n_28447), .b(n_28466), .o(n_28489) );
in01f80 g740246 ( .a(n_40314), .o(n_40315) );
in01f80 newInst_2648 ( .a(newNet_2647), .o(newNet_2648) );
no02f80 g766424 ( .a(n_14233), .b(FE_OCP_RBN2249_n_13017), .o(n_14270) );
oa22f80 FE_RC_1700_0 ( .a(n_23447), .b(n_26081), .c(FE_OCPN1494_n_23398), .d(FE_OCP_RBN2832_n_26081), .o(n_26198) );
no02f80 g778379 ( .a(n_2510), .b(n_2404), .o(n_2561) );
in01f80 FE_OCP_RBC1211_n_31515 ( .a(n_31515), .o(FE_OCP_RBN1211_n_31515) );
na02f80 g771822 ( .a(n_9281), .b(n_9380), .o(n_9311) );
oa12f80 g739756 ( .a(n_40197), .b(n_40456), .c(n_40042), .o(n_40473) );
ao12f80 g746186 ( .a(n_35088), .b(n_35087), .c(n_35086), .o(n_35653) );
na02f80 g741751 ( .a(n_38873), .b(n_38495), .o(n_38496) );
in01f80 FE_RC_2023_0 ( .a(n_13514), .o(FE_RN_672_0) );
na02f80 g748330 ( .a(n_31783), .b(n_30328), .o(n_31836) );
in01f80 g746780 ( .a(n_32976), .o(n_32977) );
in01f80 newInst_1881 ( .a(newNet_1880), .o(newNet_1881) );
na02f80 g740636 ( .a(n_39545), .b(n_39556), .o(n_39989) );
na02f80 g764578 ( .a(n_16509), .b(n_16508), .o(n_16510) );
ao12f80 g759371 ( .a(n_20539), .b(n_20693), .c(n_20492), .o(n_20802) );
ao12f80 g776744 ( .a(n_3856), .b(n_4028), .c(n_3862), .o(n_4039) );
no02f80 g740073 ( .a(n_39977), .b(n_40007), .o(n_40008) );
na02f80 FE_RC_2990_0 ( .a(FE_RN_1305_0), .b(n_9849), .o(FE_RN_1306_0) );
no02f80 g781092 ( .a(n_275), .b(n_264), .o(n_282) );
oa22f80 FE_RC_809_0 ( .a(n_7498), .b(n_8376), .c(n_7499), .d(n_8386), .o(n_8474) );
in01f80 g750573 ( .a(n_29450), .o(n_29449) );
oa12f80 g763029 ( .a(n_17482), .b(n_17588), .c(n_17406), .o(n_17678) );
in01f80 FE_OCP_RBC3220_n_21358 ( .a(FE_OCP_RBN3219_n_21358), .o(FE_OCP_RBN3220_n_21358) );
na02f80 g736937 ( .a(n_43038), .b(n_46941), .o(n_43213) );
na02f80 g751486 ( .a(n_28798), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_30_), .o(n_28799) );
in01f80 g751512 ( .a(n_28865), .o(n_28866) );
no02f80 FE_RC_2789_0 ( .a(n_34037), .b(FE_RN_1191_0), .o(FE_RN_1192_0) );
in01f80 FE_OCP_RBC1682_n_33491 ( .a(FE_OCP_RBN1680_n_33491), .o(FE_OCP_RBN1682_n_33491) );
na02f80 g760388 ( .a(n_20098), .b(FE_OCP_RBN2511_n_19884), .o(n_20129) );
no02f80 g763113 ( .a(n_17545), .b(n_17544), .o(n_17546) );
oa12f80 g760345 ( .a(n_20783), .b(n_20782), .c(n_20781), .o(n_20871) );
in01f80 g778104 ( .a(n_3026), .o(n_3027) );
no02f80 g753642 ( .a(n_26659), .b(n_26691), .o(n_26718) );
in01f80 newInst_3515 ( .a(newNet_3514), .o(newNet_3515) );
no02f80 g757441 ( .a(n_22990), .b(n_22989), .o(n_22991) );
in01f80 newInst_1870 ( .a(newNet_1869), .o(newNet_1870) );
in01f80 FE_OCP_RBC2400_n_2885 ( .a(n_2885), .o(FE_OCP_RBN2400_n_2885) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_29_ ( .ck(newNet_1376), .d(n_36728), .o(delay_sub_ln23_unr29_stage9_stallmux_q_2_) );
in01f80 g772747 ( .a(n_45828), .o(n_8254) );
na02f80 g781077 ( .a(n_262), .b(n_48), .o(n_269) );
in01f80 newInst_3108 ( .a(newNet_3107), .o(newNet_3108) );
no02f80 g738066 ( .a(n_42116), .b(n_42115), .o(n_42114) );
no02f80 g749784 ( .a(n_31249), .b(n_31324), .o(n_31283) );
in01f80 newInst_123 ( .a(newNet_122), .o(newNet_123) );
in01f80 newInst_3416 ( .a(newNet_1854), .o(newNet_3416) );
in01f80 newInst_898 ( .a(newNet_603), .o(newNet_898) );
ao22s80 FE_RC_231_0 ( .a(n_13956), .b(n_13045), .c(n_13046), .d(n_13955), .o(n_14099) );
in01f80 FE_OCP_RBC3668_n_20812 ( .a(FE_OCP_RBN3667_n_20812), .o(FE_OCP_RBN3668_n_20812) );
no02f80 g774468 ( .a(n_6676), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_16_), .o(n_6836) );
oa22f80 FE_RC_3839_0 ( .a(n_32754), .b(n_32659), .c(n_32715), .d(n_32660), .o(n_32784) );
in01f80 FE_RC_1634_0 ( .a(n_11991), .o(FE_RN_453_0) );
ao12f80 g778940 ( .a(n_2254), .b(n_2260), .c(n_2253), .o(n_2327) );
no02f80 g770425 ( .a(n_10525), .b(n_10563), .o(n_10600) );
oa12f80 g739245 ( .a(n_40889), .b(n_45153), .c(n_40891), .o(n_40921) );
ms00f80 delay_xor_ln22_unr6_stage3_stallmux_q_reg_9_ ( .ck(newNet_203), .d(n_46173), .o(delay_xor_ln22_unr6_stage3_stallmux_q_9_) );
no02f80 g749186 ( .a(n_30714), .b(FE_OCP_RBN3674_FE_RN_1581_0), .o(n_30750) );
no02f80 FE_RC_997_0 ( .a(FE_RN_285_0), .b(FE_OCP_RBN3820_n_44061), .o(FE_RN_287_0) );
in01f80 newInst_2759 ( .a(newNet_2758), .o(newNet_2759) );
oa12f80 g753802 ( .a(n_26278), .b(n_26425), .c(n_26362), .o(n_26525) );
in01f80 g764232 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_11_), .o(n_17995) );
in01f80 g765047 ( .a(n_15497), .o(n_15611) );
na02f80 g772720 ( .a(n_8107), .b(n_7817), .o(n_8162) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_20_ ( .ck(newNet_1850), .d(n_16846), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_20_) );
na02f80 g740279 ( .a(n_40310), .b(n_39807), .o(n_40363) );
no02f80 FE_RC_3196_0 ( .a(FE_RN_1420_0), .b(n_7247), .o(n_7320) );
ao12f80 g749661 ( .a(n_31258), .b(n_31295), .c(FE_OCP_RBN3013_n_31117), .o(n_31396) );
na02f80 g773870 ( .a(n_6953), .b(delay_add_ln22_unr5_stage3_stallmux_q_9_), .o(n_7049) );
oa12f80 g747136 ( .a(n_32854), .b(n_32856), .c(n_32853), .o(n_32927) );
na02f80 g768753 ( .a(n_12122), .b(n_12121), .o(n_12123) );
no02f80 g741688 ( .a(FE_OCP_RBN2352_n_38534), .b(n_38778), .o(n_38567) );
na02f80 g772977 ( .a(n_7756), .b(n_7677), .o(n_7799) );
in01f80 FE_OCP_RBC3219_n_21358 ( .a(FE_OCP_RBN3218_n_21358), .o(FE_OCP_RBN3219_n_21358) );
in01f80 g778018 ( .a(n_3673), .o(n_3155) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_6_ ( .ck(newNet_3477), .d(n_21602), .o(delay_add_ln22_unr14_stage6_stallmux_q_6_) );
oa12f80 g757610 ( .a(n_22643), .b(n_23221), .c(n_22729), .o(n_23260) );
no02f80 g773711 ( .a(n_7335), .b(n_7333), .o(n_7334) );
in01f80 g760534 ( .a(n_19969), .o(n_20044) );
in01f80 g738326 ( .a(n_41915), .o(n_41884) );
oa12f80 g738178 ( .a(n_41987), .b(n_41995), .c(n_41986), .o(n_42013) );
in01f80 g750885 ( .a(n_29034), .o(n_29035) );
in01f80 g746984 ( .a(n_32936), .o(n_33276) );
na02f80 g753725 ( .a(n_26479), .b(n_26506), .o(n_26480) );
in01f80 newInst_974 ( .a(newNet_973), .o(newNet_974) );
na02f80 g746339 ( .a(n_33525), .b(n_33524), .o(n_33526) );
na02f80 g740000 ( .a(n_39956), .b(n_39858), .o(n_40021) );
no02f80 g759674 ( .a(n_20350), .b(n_20282), .o(n_20421) );
na02f80 g754550 ( .a(n_26865), .b(n_26864), .o(n_26903) );
na02f80 g755131 ( .a(n_25373), .b(n_24451), .o(n_25500) );
ao22s80 g736290 ( .a(n_43877), .b(n_43428), .c(n_43876), .d(n_43427), .o(n_43901) );
oa12f80 g739047 ( .a(n_41088), .b(n_41087), .c(n_41086), .o(n_41121) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_1_ ( .ck(newNet_962), .d(n_22535), .o(delay_xor_ln21_unr15_stage6_stallmux_q_1_) );
no02f80 g752346 ( .a(n_27829), .b(delay_add_ln22_unr17_stage7_stallmux_q_0_), .o(n_27830) );
oa22f80 FE_RC_957_0 ( .a(n_28336), .b(n_32429), .c(n_32566), .d(n_32471), .o(n_32545) );
in01f80 FE_OCP_RBC2504_n_13896 ( .a(FE_OCP_RBN2500_n_13896), .o(FE_OCP_RBN2504_n_13896) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_8_ ( .ck(newNet_141), .d(n_46388), .o(delay_xor_ln22_unr9_stage4_stallmux_q_8_) );
na02f80 g765164 ( .a(n_15929), .b(n_15841), .o(n_15972) );
in01f80 g759790 ( .a(n_21859), .o(n_21860) );
in01f80 g761543 ( .a(n_18897), .o(n_18898) );
in01f80 g777867 ( .a(n_3250), .o(n_3251) );
na02f80 g737023 ( .a(n_43103), .b(n_42772), .o(n_43133) );
in01f80 newInst_1808 ( .a(newNet_1807), .o(newNet_1808) );
in01f80 newInst_2701 ( .a(newNet_2700), .o(newNet_2701) );
no02f80 g773973 ( .a(n_7217), .b(delay_xor_ln22_unr6_stage3_stallmux_q_24_), .o(n_7271) );
in01f80 FE_RC_4176_0 ( .a(n_33870), .o(FE_RN_1823_0) );
in01f80 g757437 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .o(n_23034) );
in01f80 g762051 ( .a(n_18631), .o(n_18632) );
no02f80 g742830 ( .a(n_37286), .b(n_37034), .o(n_37297) );
in01f80 g736681 ( .a(n_43116), .o(n_43117) );
in01f80 newInst_2614 ( .a(newNet_2613), .o(newNet_2614) );
no02f80 g753101 ( .a(n_27384), .b(n_27667), .o(n_27465) );
in01f80 g759846 ( .a(n_22393), .o(n_22484) );
in01f80 g745642 ( .a(n_35525), .o(n_36022) );
no02f80 g743340 ( .a(n_36703), .b(n_36750), .o(n_36755) );
oa22f80 FE_RC_1522_0 ( .a(n_24350), .b(n_27772), .c(n_27796), .d(n_27745), .o(n_27818) );
in01f80 newInst_1266 ( .a(newNet_611), .o(newNet_1266) );
no02f80 g776430 ( .a(n_4538), .b(n_4176), .o(n_4634) );
in01f80 g746750 ( .a(n_32980), .o(n_32951) );
in01f80 newInst_1469 ( .a(newNet_1468), .o(newNet_1469) );
oa12f80 g746362 ( .a(n_33487), .b(n_33486), .c(n_33485), .o(n_33539) );
in01f80 newInst_3748 ( .a(newNet_3747), .o(newNet_3748) );
na02f80 g738165 ( .a(n_42003), .b(n_41706), .o(n_42004) );
no02f80 g757014 ( .a(n_23803), .b(n_24087), .o(n_24045) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_4_ ( .ck(newNet_2617), .d(n_21276), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_4_) );
no02f80 g762972 ( .a(n_17962), .b(n_17961), .o(n_17963) );
in01f80 g769267 ( .a(n_11752), .o(n_11712) );
na02f80 g771303 ( .a(n_9782), .b(n_9781), .o(n_9783) );
na02f80 g772631 ( .a(n_8225), .b(n_8145), .o(n_8359) );
no02f80 g740186 ( .a(n_39812), .b(n_39546), .o(n_40111) );
na02f80 FE_RC_2478_0 ( .a(FE_RN_999_0), .b(n_40453), .o(n_40468) );
no02f80 g756770 ( .a(n_23439), .b(n_23462), .o(n_23500) );
ao12f80 g777608 ( .a(n_3449), .b(n_3456), .c(n_3448), .o(n_5165) );
na02f80 g743120 ( .a(FE_OCP_RBN3355_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_10_), .o(n_37102) );
in01f80 g748357 ( .a(n_33279), .o(n_32777) );
na02f80 g779146 ( .a(n_1935), .b(n_1904), .o(n_1956) );
in01f80 g745008 ( .a(n_34903), .o(n_34932) );
in01f80 g783842 ( .a(n_17533), .o(n_45525) );
in01f80 g743835 ( .a(n_35876), .o(n_35877) );
no03m80 FE_RC_3333_0 ( .a(n_33717), .b(n_33828), .c(n_33786), .o(n_33962) );
no02f80 g778729 ( .a(n_2277), .b(n_2270), .o(n_2330) );
na02f80 g771290 ( .a(n_9834), .b(n_9833), .o(n_9835) );
in01f80 g779433 ( .a(n_1534), .o(n_1535) );
in01f80 g739038 ( .a(n_41133), .o(n_41158) );
in01f80 g737927 ( .a(n_42302), .o(n_42274) );
oa22f80 g762766 ( .a(n_17799), .b(n_17794), .c(n_17846), .d(n_17795), .o(n_19314) );
no02f80 g749275 ( .a(n_30682), .b(n_30709), .o(n_30829) );
no02f80 g760824 ( .a(FE_OCP_RBN3493_n_19390), .b(n_18010), .o(n_19473) );
ao22s80 g746568 ( .a(n_34666), .b(n_34579), .c(n_34810), .d(n_34614), .o(n_35110) );
na02f80 g739228 ( .a(n_40890), .b(n_40888), .o(n_40906) );
ao22s80 FE_RC_3904_0 ( .a(n_30466), .b(n_30427), .c(n_27014), .d(n_30428), .o(n_30500) );
na02f80 g739268 ( .a(n_40762), .b(n_44769), .o(n_40853) );
ao12f80 g738608 ( .a(n_41571), .b(n_41716), .c(n_41492), .o(n_41965) );
no02f80 g755062 ( .a(n_25077), .b(n_24972), .o(n_25152) );
na03f80 g774149 ( .a(n_6607), .b(n_6642), .c(n_6577), .o(n_6745) );
in01f80 g753565 ( .a(n_26835), .o(n_26836) );
in01f80 newInst_1286 ( .a(newNet_1285), .o(newNet_1286) );
no02f80 g740355 ( .a(n_39721), .b(n_39674), .o(n_39733) );
no02f80 g738338 ( .a(n_41732), .b(n_41668), .o(n_41775) );
na02f80 g775141 ( .a(n_6187), .b(n_6066), .o(n_6140) );
oa12f80 g780428 ( .a(n_675), .b(n_707), .c(n_687), .o(n_715) );
na02f80 g773036 ( .a(n_8014), .b(n_8013), .o(n_8079) );
na02f80 g776488 ( .a(n_4430), .b(n_4143), .o(n_4509) );
in01f80 FE_RC_3676_0 ( .a(FE_OCPN1403_n_21007), .o(FE_RN_1615_0) );
in01f80 newInst_1612 ( .a(newNet_1611), .o(newNet_1612) );
ao12f80 g776809 ( .a(n_3815), .b(n_4139), .c(n_3940), .o(n_4297) );
no02f80 g747745 ( .a(n_33792), .b(n_33743), .o(n_33682) );
na02f80 FE_RC_2606_0 ( .a(FE_RN_1084_0), .b(n_17954), .o(FE_RN_1083_0) );
in01f80 g750096 ( .a(n_29918), .o(n_29919) );
na02f80 FE_RC_2301_0 ( .a(FE_RN_868_0), .b(n_25288), .o(FE_RN_869_0) );
na02f80 g750823 ( .a(FE_OCP_RBN2281_n_29111), .b(FE_OCP_RBN2264_n_29033), .o(n_29211) );
in01f80 newInst_3055 ( .a(newNet_3054), .o(newNet_3055) );
no02f80 FE_RC_153_0 ( .a(FE_RN_46_0), .b(FE_RN_45_0), .o(FE_RN_47_0) );
in01f80 g748317 ( .a(n_31800), .o(n_31801) );
no02f80 g770562 ( .a(n_10455), .b(n_10523), .o(n_10640) );
no02f80 g764695 ( .a(n_15981), .b(n_16067), .o(n_16140) );
no02f80 g777700 ( .a(n_3303), .b(n_3172), .o(n_3304) );
no02f80 g762118 ( .a(n_18775), .b(n_18666), .o(n_18910) );
na02f80 g765395 ( .a(n_15330), .b(n_15252), .o(n_15369) );
na02f80 g762283 ( .a(n_18617), .b(n_18729), .o(n_19231) );
in01f80 FE_RC_626_0 ( .a(n_32579), .o(FE_RN_193_0) );
ms00f80 delay_sub_ln23_0_unr15_stage6_stallmux_q_reg ( .ck(newNet_1777), .d(n_21691), .o(delay_sub_ln23_0_unr15_stage6_stallmux_q) );
in01f80 g771852 ( .a(n_9435), .o(n_9436) );
na02f80 g737587 ( .a(n_42746), .b(n_42445), .o(n_42767) );
oa12f80 g778753 ( .a(n_2223), .b(n_2222), .c(n_2221), .o(n_2473) );
in01f80 newInst_237 ( .a(newNet_235), .o(newNet_237) );
in01f80 g738012 ( .a(n_42179), .o(n_42180) );
in01f80 newInst_2881 ( .a(newNet_1784), .o(newNet_2881) );
in01f80 newInst_956 ( .a(newNet_112), .o(newNet_956) );
no02f80 g780888 ( .a(n_374), .b(n_385), .o(n_391) );
na02f80 g742867 ( .a(n_37249), .b(n_37248), .o(n_37250) );
in01f80 g748320 ( .a(n_31840), .o(n_31841) );
in01f80 g766151 ( .a(n_14554), .o(n_14577) );
in01f80 newInst_1637 ( .a(newNet_1636), .o(newNet_1637) );
in01f80 g772304 ( .a(n_8548), .o(n_8562) );
in01f80 g780170 ( .a(n_1142), .o(n_1130) );
in01f80 g746604 ( .a(n_34635), .o(n_34693) );
oa22f80 g777836 ( .a(n_3186), .b(n_2733), .c(n_3228), .d(n_2732), .o(n_3264) );
oa12f80 g757678 ( .a(n_22417), .b(n_22625), .c(n_22415), .o(n_22703) );
na02f80 g745379 ( .a(FE_OCP_RBN2992_n_35539), .b(n_35845), .o(n_35929) );
in01f80 FE_RC_3593_0 ( .a(FE_OCPN1429_n_23792), .o(FE_RN_1568_0) );
in01f80 g765101 ( .a(n_15382), .o(n_15420) );
na02f80 g767547 ( .a(n_13322), .b(n_13193), .o(n_13323) );
in01f80 g763704 ( .a(n_17537), .o(n_17607) );
in01f80 FE_RC_1303_0 ( .a(FE_OCP_RBN1342_n_19077), .o(FE_RN_381_0) );
no02f80 g751867 ( .a(n_28217), .b(n_28056), .o(n_28218) );
oa22f80 g784543 ( .a(n_11655), .b(FE_OFN802_n_46285), .c(n_11527), .d(FE_OCP_RBN3043_n_46337), .o(n_46364) );
na02f80 g776441 ( .a(n_4529), .b(FE_OCP_RBN3577_n_4528), .o(n_4659) );
no02f80 g746639 ( .a(n_33340), .b(n_33269), .o(n_33368) );
in01f80 g752775 ( .a(n_27193), .o(n_27158) );
in01f80 newInst_739 ( .a(newNet_738), .o(newNet_739) );
in01f80 FE_OCP_RBC2297_n_2438 ( .a(FE_OCP_RBN2292_n_2438), .o(FE_OCP_RBN2297_n_2438) );
ms00f80 delay_sub_ln23_0_unr22_stage8_stallmux_q_reg ( .ck(newNet_1554), .d(n_30156), .o(delay_sub_ln23_0_unr22_stage8_stallmux_q) );
in01f80 newInst_1382 ( .a(newNet_1319), .o(newNet_1382) );
in01f80 g780327 ( .a(n_1046), .o(n_974) );
na02f80 g737714 ( .a(n_42392), .b(n_42124), .o(n_42445) );
in01f80 FE_OCP_RBC2631_n_29947 ( .a(n_29947), .o(FE_OCP_RBN2631_n_29947) );
no02f80 g775914 ( .a(n_4925), .b(FE_OCP_RBN2728_n_4219), .o(n_4952) );
in01f80 g764583 ( .a(n_16181), .o(n_16182) );
in01f80 g772843 ( .a(n_8154), .o(n_8155) );
na02f80 g778175 ( .a(n_2864), .b(n_2863), .o(n_2956) );
in01f80 FE_OCP_RBC2806_n_30643 ( .a(n_30643), .o(FE_OCP_RBN2806_n_30643) );
oa12f80 g736319 ( .a(n_337), .b(n_43853), .c(n_43918), .o(n_43891) );
in01f80 newInst_696 ( .a(newNet_695), .o(newNet_696) );
na02f80 g746883 ( .a(FE_OCP_RBN3387_n_33108), .b(delay_add_ln22_unr20_stage8_stallmux_q_30_), .o(n_33377) );
na02f80 g776422 ( .a(n_4366), .b(n_4457), .o(n_4494) );
na02f80 FE_RC_2822_0 ( .a(n_34412), .b(FE_RN_1210_0), .o(FE_RN_1211_0) );
no02f80 g751596 ( .a(n_28458), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_22_), .o(n_28627) );
in01f80 g756553 ( .a(n_23818), .o(n_23819) );
in01f80 newInst_3733 ( .a(newNet_3732), .o(newNet_3733) );
no02f80 g750328 ( .a(n_29730), .b(n_29533), .o(n_29731) );
in01f80 newInst_3467 ( .a(newNet_3466), .o(newNet_3467) );
in01f80 newInst_1587 ( .a(newNet_1120), .o(newNet_1587) );
no02f80 g755686 ( .a(n_24370), .b(n_24322), .o(n_24435) );
in01f80 g741269 ( .a(n_39068), .o(n_39069) );
in01f80 g739900 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_6_), .o(n_40696) );
in01f80 newInst_1236 ( .a(newNet_1235), .o(newNet_1236) );
oa12f80 g736426 ( .a(n_344), .b(n_43761), .c(FE_OFN2_n_43918), .o(n_43818) );
no02f80 g754579 ( .a(n_25464), .b(n_25463), .o(n_25465) );
na02f80 g781014 ( .a(sin_out_12), .b(FE_OFN3_n_43918), .o(n_325) );
in01f80 newInst_912 ( .a(newNet_911), .o(newNet_912) );
in01f80 FE_OCPC940_n_7712 ( .a(FE_OCPN939_n_7712), .o(FE_OCPN940_n_7712) );
in01f80 newInst_2026 ( .a(newNet_2025), .o(newNet_2026) );
in01f80 g741889 ( .a(n_39232), .o(n_38429) );
in01f80 fopt ( .a(n_47187), .o(n_47186) );
na02f80 g739188 ( .a(n_40796), .b(n_40706), .o(n_40797) );
na02f80 g741024 ( .a(n_38915), .b(n_38860), .o(n_38967) );
na02f80 g754147 ( .a(n_25937), .b(n_23317), .o(n_26001) );
oa12f80 g773652 ( .a(n_6864), .b(n_7332), .c(n_6940), .o(n_7351) );
in01f80 g765519 ( .a(n_15714), .o(n_15715) );
in01f80 FE_OFC766_n_15670 ( .a(FE_OFN763_n_15670), .o(FE_OFN766_n_15670) );
oa22f80 FE_RC_3239_0 ( .a(FE_OCP_RBN1167_n_18949), .b(n_18950), .c(n_18949), .d(n_18859), .o(n_19011) );
in01f80 g759491 ( .a(n_20935), .o(n_20965) );
na02f80 g780891 ( .a(n_403), .b(n_437), .o(n_444) );
na02f80 g744729 ( .a(n_35154), .b(n_30614), .o(n_35235) );
na02f80 g748081 ( .a(n_31875), .b(n_31836), .o(n_31934) );
in01f80 g745285 ( .a(n_36174), .o(n_36175) );
na02f80 g741655 ( .a(n_38537), .b(n_38778), .o(n_38557) );
in01f80 g762229 ( .a(n_18149), .o(n_18150) );
na02f80 g771050 ( .a(n_9362), .b(n_9421), .o(n_9456) );
in01f80 g773934 ( .a(n_7020), .o(n_7021) );
in01f80 g738934 ( .a(n_41320), .o(n_41292) );
in01f80 g740440 ( .a(n_39967), .o(n_39931) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_3_ ( .ck(newNet_913), .d(n_27750), .o(delay_xor_ln21_unr18_stage7_stallmux_q_3_) );
in01f80 g737327 ( .a(n_42857), .o(n_42871) );
no02f80 g770879 ( .a(n_10006), .b(n_9899), .o(n_10111) );
in01f80 g771961 ( .a(n_9651), .o(n_9728) );
no02f80 FE_RC_2725_0 ( .a(FE_RN_1150_0), .b(FE_RN_1152_0), .o(n_8448) );
in01f80 FE_RC_4191_0 ( .a(n_24158), .o(FE_RN_1836_0) );
na02f80 g748636 ( .a(n_31308), .b(n_31271), .o(n_31272) );
no02f80 g762261 ( .a(n_18726), .b(n_18725), .o(n_18767) );
no02f80 g737579 ( .a(n_42288), .b(n_42287), .o(n_42314) );
ao12f80 g740839 ( .a(n_39076), .b(n_39380), .c(n_39045), .o(n_39431) );
in01f80 newInst_1689 ( .a(newNet_1688), .o(newNet_1689) );
in01f80 newInst_640 ( .a(newNet_189), .o(newNet_640) );
na02f80 g773924 ( .a(n_7013), .b(n_7012), .o(n_7014) );
no02f80 g755592 ( .a(n_24469), .b(FE_OCP_RBN2366_n_24372), .o(n_24570) );
in01f80 g765982 ( .a(n_14697), .o(n_14724) );
in01f80 g770319 ( .a(n_10692), .o(n_10693) );
oa22f80 FE_RC_3205_0 ( .a(FE_RN_1424_0), .b(FE_OCPN875_n_44672), .c(n_1064), .d(n_44637), .o(n_1343) );
na02f80 g748583 ( .a(n_31336), .b(n_31245), .o(n_31365) );
in01f80 g766950 ( .a(n_14297), .o(n_14389) );
no02f80 g751000 ( .a(n_30161), .b(n_30129), .o(n_30902) );
na02f80 g744510 ( .a(n_36745), .b(n_36744), .o(n_36746) );
oa12f80 g749701 ( .a(n_31311), .b(n_31417), .c(n_31416), .o(n_31458) );
ao22s80 g773487 ( .a(n_7525), .b(n_6963), .c(n_7493), .d(n_6962), .o(n_7982) );
na02f80 g778332 ( .a(n_3178), .b(n_2438), .o(n_2649) );
in01f80 newInst_215 ( .a(newNet_66), .o(newNet_215) );
oa12f80 g737259 ( .a(n_42657), .b(n_42918), .c(n_42608), .o(n_42928) );
na02f80 g758814 ( .a(n_22117), .b(n_21592), .o(n_22210) );
no02f80 g748834 ( .a(n_31265), .b(n_31264), .o(n_31297) );
in01f80 newInst_3533 ( .a(newNet_3532), .o(newNet_3533) );
oa22f80 g784373 ( .a(FE_OFN806_n_46196), .b(n_6435), .c(FE_OFN84_n_46137), .d(n_6407), .o(n_46179) );
no02f80 g754717 ( .a(FE_OCP_RBN2959_n_26231), .b(n_26546), .o(n_26609) );
no02f80 g738518 ( .a(FE_OCP_RBN2312_n_41420), .b(n_41626), .o(n_41667) );
in01f80 g778673 ( .a(FE_OCPN850_n_2306), .o(n_2274) );
na02f80 g748941 ( .a(n_31054), .b(n_31053), .o(n_31055) );
in01f80 g762782 ( .a(n_17914), .o(n_17998) );
in01f80 newInst_2121 ( .a(newNet_2120), .o(newNet_2121) );
ao12f80 g742363 ( .a(n_37798), .b(n_37797), .c(n_37796), .o(n_38713) );
oa12f80 g759607 ( .a(n_21698), .b(n_21601), .c(n_21374), .o(n_21724) );
no02f80 g781314 ( .a(beta_31), .b(beta_17), .o(n_53) );
no02f80 g763742 ( .a(n_16685), .b(n_16600), .o(n_16755) );
in01f80 g739781 ( .a(n_40496), .o(n_40497) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_24_ ( .ck(newNet_2380), .d(FE_OCP_RBN1328_n_36489), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_24_) );
na02f80 g752905 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_28_), .o(n_28132) );
no02f80 g760415 ( .a(n_20064), .b(n_19943), .o(n_20080) );
no02f80 g752955 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .o(n_28050) );
in01f80 newInst_3617 ( .a(newNet_3616), .o(newNet_3617) );
in01f80 g779594 ( .a(n_1494), .o(n_1401) );
in01f80 g778926 ( .a(n_2169), .o(n_2200) );
oa22f80 g776880 ( .a(n_3875), .b(n_3743), .c(n_3876), .d(n_3799), .o(n_4099) );
no02f80 g758055 ( .a(n_23058), .b(n_22807), .o(n_23529) );
no02f80 g754456 ( .a(n_25545), .b(n_25272), .o(n_25635) );
in01f80 newInst_2542 ( .a(newNet_1617), .o(newNet_2542) );
ao12f80 g774169 ( .a(n_7141), .b(n_6872), .c(delay_xor_ln22_unr6_stage3_stallmux_q_19_), .o(n_7265) );
no02f80 g767885 ( .a(n_12728), .b(delay_add_ln22_unr8_stage4_stallmux_q_21_), .o(n_12766) );
no02f80 g775418 ( .a(n_5541), .b(n_5499), .o(n_5605) );
in01f80 g770742 ( .a(n_10145), .o(n_10188) );
in01f80 g739261 ( .a(n_40952), .o(n_40953) );
in01f80 newInst_3500 ( .a(newNet_3499), .o(newNet_3500) );
in01f80 newInst_370 ( .a(newNet_360), .o(newNet_370) );
na02f80 g740541 ( .a(n_39643), .b(n_39657), .o(n_39658) );
in01f80 g757353 ( .a(n_23064), .o(n_23101) );
in01f80 g752223 ( .a(delay_xor_ln21_unr18_stage7_stallmux_q_12_), .o(n_27944) );
ao12f80 g745258 ( .a(n_34747), .b(n_34675), .c(n_34369), .o(n_34748) );
no02f80 FE_RC_4161_0 ( .a(FE_RN_1812_0), .b(n_33484), .o(n_33501) );
in01f80 g754619 ( .a(n_27131), .o(FE_RN_1481_0) );
in01f80 FE_RC_1144_0 ( .a(n_47240), .o(FE_RN_346_0) );
no02f80 g745740 ( .a(n_34149), .b(n_34100), .o(n_34264) );
in01f80 g741635 ( .a(n_38635), .o(n_38636) );
in01f80 FE_RC_3351_0 ( .a(n_20744), .o(FE_RN_1461_0) );
in01f80 g780140 ( .a(n_1194), .o(n_1185) );
na02f80 g743398 ( .a(n_36653), .b(n_36633), .o(n_36703) );
na02f80 g777403 ( .a(n_3627), .b(n_3626), .o(n_3651) );
na02f80 FE_RC_2279_0 ( .a(FE_RN_850_0), .b(n_28079), .o(FE_RN_851_0) );
in01f80 g746927 ( .a(n_32897), .o(n_32916) );
na02f80 g765004 ( .a(n_15497), .b(n_15609), .o(n_15536) );
na02f80 g778590 ( .a(n_2639), .b(n_2710), .o(n_2732) );
in01f80 g747977 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_12_), .o(n_32082) );
na02f80 g756046 ( .a(n_25026), .b(n_25133), .o(n_25163) );
in01f80 g769209 ( .a(n_11680), .o(n_11681) );
in01f80 g772560 ( .a(n_8400), .o(n_8401) );
ao12f80 g745271 ( .a(FE_OCP_RBN2987_n_35539), .b(n_36171), .c(n_36022), .o(n_36023) );
no02f80 g780629 ( .a(n_779), .b(n_839), .o(n_900) );
in01f80 g744751 ( .a(n_35178), .o(n_35179) );
no02f80 g769331 ( .a(n_10708), .b(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(n_11795) );
no02f80 g740329 ( .a(n_40245), .b(n_39937), .o(n_40357) );
oa22f80 g750974 ( .a(n_28872), .b(n_28865), .c(n_28873), .d(n_28866), .o(n_29898) );
no02f80 g747156 ( .a(n_32906), .b(delay_add_ln22_unr20_stage8_stallmux_q_6_), .o(n_32967) );
na02f80 g746828 ( .a(n_33157), .b(n_33156), .o(n_33182) );
na02f80 g745851 ( .a(n_34097), .b(n_34096), .o(n_34148) );
na02f80 g742237 ( .a(FE_OCP_RBN3425_n_44881), .b(n_38047), .o(n_38135) );
ao12f80 g741890 ( .a(n_38354), .b(n_38358), .c(n_38353), .o(n_39232) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_0_ ( .ck(newNet_2694), .d(n_20378), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_0_) );
in01f80 FE_OCP_RBC3013_n_31117 ( .a(FE_OCP_RBN3702_n_31064), .o(FE_OCP_RBN3013_n_31117) );
na02f80 g769396 ( .a(n_44336), .b(n_10293), .o(n_11538) );
in01f80 FE_RC_3539_0 ( .a(n_18866), .o(FE_RN_1532_0) );
ao12f80 g748021 ( .a(n_31823), .b(n_31777), .c(n_31897), .o(n_31936) );
na02f80 g769091 ( .a(n_11509), .b(n_11485), .o(n_11555) );
na02f80 g755808 ( .a(n_24291), .b(n_23278), .o(n_24373) );
in01f80 newInst_1580 ( .a(newNet_1579), .o(newNet_1580) );
no02f80 g745430 ( .a(FE_OCP_RBN2987_n_35539), .b(n_35392), .o(n_35839) );
in01f80 g757483 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_4_), .o(n_22939) );
in01f80 FE_OCP_RBC3842_n_19555 ( .a(n_19555), .o(FE_OCP_RBN3842_n_19555) );
no02f80 g747534 ( .a(n_33814), .b(n_33793), .o(n_35542) );
in01f80 FE_OCP_RBC3333_n_44962 ( .a(n_44962), .o(FE_OCP_RBN3333_n_44962) );
in01f80 newInst_1674 ( .a(newNet_1673), .o(newNet_1674) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_11_ ( .ck(newNet_928), .d(n_27863), .o(delay_xor_ln21_unr18_stage7_stallmux_q_11_) );
na02f80 g769580 ( .a(n_11408), .b(n_11390), .o(n_11494) );
in01f80 newInst_3454 ( .a(newNet_970), .o(newNet_3454) );
oa12f80 g759259 ( .a(n_21758), .b(n_21757), .c(n_21756), .o(n_21802) );
oa22f80 FE_RC_4263_0 ( .a(n_32678), .b(FE_OCP_RBN2153_n_32772), .c(n_32679), .d(n_32772), .o(n_32827) );
ao12f80 g745180 ( .a(n_34467), .b(FE_OCP_DRV_N1594_n_34494), .c(n_34466), .o(n_34540) );
in01f80 g772317 ( .a(n_8684), .o(n_8760) );
ao12f80 g766674 ( .a(n_13855), .b(n_13854), .c(n_13853), .o(n_15791) );
in01f80 g740318 ( .a(n_39781), .o(n_39816) );
no02f80 g750998 ( .a(n_28868), .b(n_28609), .o(n_28918) );
no02f80 FE_RC_3556_0 ( .a(FE_RN_1543_0), .b(n_13229), .o(n_13310) );
no02f80 g746741 ( .a(n_34172), .b(n_34171), .o(n_34173) );
na02f80 FE_RC_3085_0 ( .a(n_20926), .b(FE_RN_1361_0), .o(n_20947) );
na02f80 g745548 ( .a(n_34342), .b(n_34260), .o(n_34375) );
in01f80 g751757 ( .a(n_28320), .o(n_28321) );
no02f80 g761821 ( .a(n_18375), .b(n_17423), .o(n_18437) );
in01f80 g767278 ( .a(n_13698), .o(n_13699) );
na02f80 g780735 ( .a(n_605), .b(n_604), .o(n_606) );
na02f80 g768413 ( .a(n_12361), .b(n_12208), .o(n_12376) );
oa12f80 g784656 ( .a(n_11361), .b(n_11316), .c(n_11187), .o(n_46986) );
in01f80 g773059 ( .a(n_7745), .o(n_7789) );
no02f80 g744302 ( .a(FE_OCP_RBN2903_n_44174), .b(FE_OCP_RBN2712_n_35075), .o(n_36000) );
no02f80 FE_RC_378_0 ( .a(FE_RN_113_0), .b(n_12458), .o(n_12528) );
in01f80 g752560 ( .a(n_27686), .o(n_27662) );
na02f80 FE_RC_2346_0 ( .a(FE_RN_899_0), .b(n_32505), .o(FE_RN_900_0) );
no02f80 g761859 ( .a(n_18321), .b(n_18346), .o(n_18718) );
in01f80 g767924 ( .a(n_12921), .o(n_12922) );
in01f80 g749685 ( .a(n_31259), .o(n_31638) );
oa12f80 g750170 ( .a(n_30901), .b(n_30923), .c(n_30900), .o(n_31371) );
in01f80 g754247 ( .a(FE_OFN507_n_25938), .o(n_25962) );
oa22f80 FE_RC_3268_0 ( .a(n_11804), .b(n_11990), .c(n_11803), .d(n_12025), .o(n_12212) );
in01f80 g745982 ( .a(n_35763), .o(n_35298) );
no02f80 g765568 ( .a(n_15103), .b(n_14396), .o(n_15293) );
no02f80 g746818 ( .a(n_32914), .b(n_32920), .o(n_33350) );
oa22f80 g745328 ( .a(n_36049), .b(n_35804), .c(FE_OCP_RBN2995_n_35539), .d(n_35259), .o(n_36217) );
no02f80 g756264 ( .a(n_24096), .b(n_24081), .o(n_24157) );
oa12f80 g770342 ( .a(n_10688), .b(n_10687), .c(n_10686), .o(n_10744) );
in01f80 g776583 ( .a(n_4451), .o(n_4452) );
no02f80 g778949 ( .a(n_2143), .b(n_2134), .o(n_2135) );
in01f80 FE_OCP_RBC2219_n_12698 ( .a(n_12698), .o(FE_OCP_RBN2219_n_12698) );
in01f80 FE_RC_3135_0 ( .a(n_15656), .o(FE_RN_1390_0) );
in01f80 FE_RC_509_0 ( .a(n_28191), .o(FE_RN_157_0) );
in01f80 g764206 ( .a(n_16820), .o(n_16821) );
ms00f80 cos_out_reg_16_ ( .ck(newNet_3741), .d(n_43817), .o(cos_out_16) );
na02f80 g770998 ( .a(n_9888), .b(n_9845), .o(n_9927) );
in01f80 FE_OCP_RBC3707_n_16649 ( .a(n_16649), .o(FE_OCP_RBN3707_n_16649) );
ms00f80 delay_xor_ln21_unr18_stage7_stallmux_q_reg_6_ ( .ck(newNet_903), .d(n_27815), .o(delay_xor_ln21_unr18_stage7_stallmux_q_6_) );
in01f80 g748709 ( .a(n_44042), .o(n_32605) );
in01f80 FE_OCP_RBC2582_n_3734 ( .a(FE_OCP_RBN2579_n_3734), .o(FE_OCP_RBN2582_n_3734) );
in01f80 newInst_829 ( .a(newNet_828), .o(newNet_829) );
ao12f80 g779801 ( .a(n_1686), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_23_), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_24_), .o(n_1722) );
no02f80 g753452 ( .a(n_26844), .b(n_25363), .o(n_26918) );
in01f80 g747511 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_25_), .o(n_32991) );
na02f80 g764968 ( .a(n_15242), .b(n_15157), .o(n_15357) );
in01f80 newInst_366 ( .a(newNet_365), .o(newNet_366) );
in01f80 g755091 ( .a(n_25076), .o(n_25077) );
no02f80 g756583 ( .a(n_23599), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_19_), .o(n_23679) );
ao12f80 g779263 ( .a(n_1737), .b(n_1736), .c(n_1735), .o(n_2250) );
oa12f80 g747637 ( .a(n_31788), .b(n_32169), .c(n_32168), .o(n_32196) );
no02f80 g749903 ( .a(n_30019), .b(n_30018), .o(n_30020) );
no02f80 g774332 ( .a(n_6806), .b(delay_xor_ln21_unr6_stage3_stallmux_q_14_), .o(n_6924) );
in01f80 FE_OCP_RBC3653_n_10100 ( .a(FE_OCP_RBN3652_n_10100), .o(FE_OCP_RBN3653_n_10100) );
na02f80 g760853 ( .a(n_19363), .b(n_18675), .o(n_19470) );
in01f80 FE_OCP_RBC2649_n_3840 ( .a(n_3840), .o(FE_OCP_RBN2649_n_3840) );
no02f80 g741449 ( .a(n_38770), .b(n_38778), .o(n_38771) );
in01f80 FE_RC_508_0 ( .a(n_28189), .o(FE_RN_156_0) );
in01f80 g768070 ( .a(n_12748), .o(n_12717) );
in01f80 newInst_2170 ( .a(newNet_1124), .o(newNet_2170) );
na02f80 g742901 ( .a(n_37135), .b(n_37010), .o(n_37011) );
in01f80 FE_OCPC902_n_44581 ( .a(FE_OCP_RBN2556_n_44576), .o(FE_OCPN902_n_44581) );
na02f80 g738523 ( .a(n_41582), .b(n_41176), .o(n_41674) );
in01f80 g751907 ( .a(n_29100), .o(n_29150) );
na02f80 g755619 ( .a(n_24499), .b(n_23944), .o(n_24565) );
na02f80 g745416 ( .a(FE_OCP_RBN2986_n_35539), .b(n_35631), .o(n_35679) );
in01f80 newInst_3020 ( .a(newNet_3019), .o(newNet_3020) );
no02f80 g760421 ( .a(n_20655), .b(n_19988), .o(n_20742) );
ms00f80 delay_sub_ln23_0_unr24_stage8_stallmux_q_reg_20_ ( .ck(newNet_1515), .d(n_32228), .o(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_) );
in01f80 newInst_1591 ( .a(newNet_1590), .o(newNet_1591) );
in01f80 g738860 ( .a(n_41322), .o(n_41421) );
na02f80 g771361 ( .a(FE_RN_1125_0), .b(n_9210), .o(n_9350) );
no02f80 g760939 ( .a(n_19254), .b(n_19277), .o(n_19358) );
in01f80 newInst_526 ( .a(newNet_293), .o(newNet_526) );
in01f80 newInst_3061 ( .a(newNet_3060), .o(newNet_3061) );
no02f80 g760975 ( .a(n_19349), .b(n_19319), .o(n_19457) );
in01f80 g748700 ( .a(n_31360), .o(n_31361) );
no02f80 g772883 ( .a(n_7992), .b(n_7991), .o(n_8084) );
no02f80 g743562 ( .a(n_36533), .b(n_36149), .o(n_36560) );
na02f80 g777349 ( .a(n_4759), .b(n_4970), .o(n_5069) );
no02f80 g775182 ( .a(n_5802), .b(n_4875), .o(n_5839) );
na03f80 g762215 ( .a(n_18568), .b(n_18665), .c(n_18664), .o(n_18666) );
na02f80 g767305 ( .a(n_13652), .b(n_13651), .o(n_13653) );
na02f80 g769307 ( .a(n_11455), .b(n_10977), .o(n_11509) );
in01f80 g740901 ( .a(n_39342), .o(n_39399) );
no02f80 g776529 ( .a(n_4421), .b(n_4357), .o(n_4588) );
in01f80 newInst_1560 ( .a(newNet_1559), .o(newNet_1560) );
no02f80 g737607 ( .a(n_42222), .b(n_42241), .o(n_42242) );
in01f80 g771217 ( .a(n_9556), .o(n_9557) );
in01f80 g757533 ( .a(delay_sub_ln21_0_unr14_stage6_stallmux_q_21_), .o(n_22717) );
in01f80 newInst_220 ( .a(newNet_219), .o(newNet_220) );
in01f80 g750020 ( .a(n_30316), .o(n_30317) );
in01f80 newInst_3068 ( .a(newNet_881), .o(newNet_3068) );
in01f80 g762904 ( .a(n_17697), .o(n_17681) );
na02f80 g749612 ( .a(n_30299), .b(n_32076), .o(n_30300) );
na02f80 g765966 ( .a(n_45520), .b(FE_OCP_RBN3528_n_13765), .o(n_14726) );
no03m80 g742434 ( .a(n_37608), .b(n_37609), .c(n_37116), .o(n_37630) );
no02f80 FE_RC_4159_0 ( .a(FE_RN_1809_0), .b(FE_RN_1810_0), .o(FE_RN_1811_0) );
na02f80 g759074 ( .a(n_21488), .b(n_21569), .o(n_21641) );
na02f80 g778418 ( .a(n_2672), .b(delay_add_ln22_unr2_stage2_stallmux_q_26_), .o(n_2790) );
ao12f80 g761782 ( .a(n_18185), .b(n_18376), .c(n_18213), .o(n_18518) );
na02f80 g741233 ( .a(n_39175), .b(n_39123), .o(n_39201) );
no02f80 g738289 ( .a(n_41839), .b(n_41838), .o(n_41840) );
in01f80 FE_OCP_RBC2275_n_24077 ( .a(n_24077), .o(FE_OCP_RBN2275_n_24077) );
no02f80 g757209 ( .a(n_44068), .b(delay_xor_ln22_unr15_stage6_stallmux_q_14_), .o(n_23079) );
no02f80 g776502 ( .a(n_4481), .b(n_4582), .o(n_4756) );
na02f80 g737522 ( .a(n_42550), .b(n_42491), .o(n_42594) );
in01f80 g762924 ( .a(n_17842), .o(n_17884) );
in01f80 FE_RC_2020_0 ( .a(n_20264), .o(FE_RN_670_0) );
oa22f80 g749443 ( .a(n_31941), .b(n_31631), .c(n_31911), .d(n_31632), .o(n_32004) );
no02f80 g779007 ( .a(n_2173), .b(n_1083), .o(n_2208) );
in01f80 FE_OCP_RBC3717_n_39913 ( .a(FE_OCP_RBN3716_n_39913), .o(FE_OCP_RBN3717_n_39913) );
in01f80 g770665 ( .a(n_10192), .o(n_10193) );
no02f80 g766901 ( .a(n_13647), .b(FE_OCPN1764_n_13646), .o(n_13657) );
na02f80 g779277 ( .a(n_1753), .b(n_959), .o(n_1834) );
in01f80 g771014 ( .a(n_9749), .o(n_9750) );
na02f80 g762968 ( .a(n_17742), .b(n_17741), .o(n_17743) );
na02f80 g740366 ( .a(FE_OCP_RBN3020_n_39942), .b(n_39810), .o(n_40310) );
na02f80 g776640 ( .a(n_4009), .b(n_3922), .o(n_4078) );
oa12f80 g757375 ( .a(n_22996), .b(n_22995), .c(n_22994), .o(n_24158) );
ao12f80 g746422 ( .a(n_33425), .b(n_33424), .c(n_33423), .o(n_34098) );
in01f80 FE_OCP_RBC2952_n_21489 ( .a(FE_OCP_RBN2951_n_21489), .o(FE_OCP_RBN2952_n_21489) );
na02f80 g776692 ( .a(n_4297), .b(n_4269), .o(n_4270) );
na02f80 g760301 ( .a(n_20834), .b(n_20927), .o(n_20928) );
in01f80 g737848 ( .a(n_42622), .o(n_42623) );
na02f80 g762167 ( .a(n_18192), .b(n_17921), .o(n_18242) );
no02f80 g777060 ( .a(n_4819), .b(n_4818), .o(n_4820) );
na02f80 g763835 ( .a(n_16640), .b(n_16637), .o(n_16684) );
in01f80 newInst_3473 ( .a(newNet_3472), .o(newNet_3473) );
ao22s80 g742037 ( .a(FE_OCP_RBN3445_n_37945), .b(n_37518), .c(FE_OCP_RBN3449_n_37945), .d(n_37545), .o(n_38393) );
ao12f80 g757764 ( .a(n_22432), .b(n_22590), .c(n_22465), .o(n_22624) );
na02f80 g775053 ( .a(n_6092), .b(n_5967), .o(n_6136) );
no02f80 g736989 ( .a(FE_OCPN1247_n_43120), .b(n_43005), .o(n_43503) );
no02f80 g737717 ( .a(n_42285), .b(n_42076), .o(n_42389) );
in01f80 g753422 ( .a(n_26989), .o(n_26990) );
in01f80 g755379 ( .a(n_24932), .o(n_24933) );
no02f80 g770248 ( .a(n_10745), .b(n_10725), .o(n_10726) );
na02f80 g752636 ( .a(n_27476), .b(n_27206), .o(n_27565) );
ao12f80 g743268 ( .a(n_37960), .b(n_37959), .c(n_37958), .o(n_38093) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_20_ ( .ck(newNet_3420), .d(n_27714), .o(delay_add_ln22_unr17_stage7_stallmux_q_20_) );
in01f80 FE_OCP_RBC2484_n_38601 ( .a(n_38601), .o(FE_OCP_RBN2484_n_38601) );
no02f80 g777099 ( .a(n_3733), .b(n_3604), .o(n_3809) );
oa12f80 g742557 ( .a(n_37273), .b(n_37421), .c(n_37471), .o(n_37509) );
in01f80 g756499 ( .a(n_23995), .o(n_23996) );
in01f80 g765906 ( .a(n_14917), .o(n_14918) );
no02f80 g769088 ( .a(n_11478), .b(n_11437), .o(n_11498) );
in01f80 FE_OCP_DRV_C1545_n_18860 ( .a(n_18860), .o(FE_OCP_DRV_N1545_n_18860) );
oa12f80 g756752 ( .a(n_23938), .b(n_23866), .c(n_23803), .o(n_24036) );
na02f80 g737730 ( .a(n_42352), .b(n_42270), .o(n_42412) );
no02f80 g755989 ( .a(n_24179), .b(n_21852), .o(n_24210) );
ao12f80 g768511 ( .a(n_12368), .b(n_45659), .c(delay_xor_ln22_unr9_stage4_stallmux_q_17_), .o(n_12387) );
no02f80 g779789 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_6_), .o(n_1451) );
oa22f80 FE_RC_3736_0 ( .a(n_36720), .b(n_36734), .c(n_36721), .d(n_36733), .o(n_36776) );
in01f80 g755321 ( .a(n_25470), .o(n_25638) );
in01f80 g776248 ( .a(n_4825), .o(n_4826) );
no02f80 FE_RC_3616_0 ( .a(n_20440), .b(n_20422), .o(n_20511) );
no02f80 g739176 ( .a(n_40881), .b(n_41120), .o(n_40958) );
oa22f80 FE_RC_2637_0 ( .a(n_8393), .b(FE_OCP_RBN3500_n_8187), .c(FE_OCP_RBN3501_n_8187), .d(FE_OCP_RBN2466_n_8393), .o(n_8569) );
na02f80 g757395 ( .a(n_44068), .b(delay_xor_ln21_unr15_stage6_stallmux_q_16_), .o(n_23161) );
na02f80 g769176 ( .a(n_11590), .b(n_11547), .o(n_11636) );
oa12f80 g770297 ( .a(n_10454), .b(n_10650), .c(n_10523), .o(n_10745) );
no02f80 g773107 ( .a(n_7997), .b(n_7954), .o(n_8605) );
no02f80 g756646 ( .a(n_23576), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_15_), .o(n_23600) );
na02f80 g755859 ( .a(n_24305), .b(delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24339) );
oa12f80 g749549 ( .a(n_30051), .b(n_45631), .c(n_30356), .o(n_30379) );
no02f80 g780501 ( .a(n_691), .b(n_706), .o(n_717) );
in01f80 FE_RC_2285_0 ( .a(n_17665), .o(FE_RN_855_0) );
in01f80 g777270 ( .a(n_3670), .o(n_3671) );
in01f80 g780584 ( .a(n_829), .o(n_884) );
na02f80 FE_RC_917_0 ( .a(FE_RN_271_0), .b(FE_RN_270_0), .o(FE_RN_272_0) );
na02f80 g739475 ( .a(n_40686), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_2_), .o(n_40820) );
na02f80 g745627 ( .a(n_34369), .b(n_33964), .o(n_34674) );
in01f80 FE_OCP_RBC1331_n_18866 ( .a(FE_OCP_RBN1330_n_18866), .o(FE_OCP_RBN1331_n_18866) );
no02f80 g755898 ( .a(n_24390), .b(n_24389), .o(n_24391) );
no02f80 g765122 ( .a(n_15125), .b(n_15162), .o(n_15281) );
in01f80 newInst_2834 ( .a(newNet_2833), .o(newNet_2834) );
na02f80 g751314 ( .a(n_29636), .b(n_29045), .o(n_29649) );
ao12f80 g766842 ( .a(n_12722), .b(n_13560), .c(FE_OCP_DRV_N3150_n_12773), .o(n_13601) );
no02f80 g773792 ( .a(n_7182), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_13_), .o(n_7204) );
in01f80 g762787 ( .a(n_17912), .o(n_17913) );
no02f80 g764287 ( .a(FE_OCP_RBN2907_n_16230), .b(n_14618), .o(n_16336) );
in01f80 g777859 ( .a(n_3224), .o(n_3225) );
ao12f80 g761773 ( .a(n_19195), .b(n_19194), .c(n_19193), .o(n_19735) );
no02f80 g746263 ( .a(n_33674), .b(n_33328), .o(n_33687) );
no02f80 g753820 ( .a(n_26358), .b(FE_OCPN1488_n_23447), .o(n_26406) );
in01f80 g755013 ( .a(FE_OCP_RBN2596_n_25181), .o(n_25270) );
na02f80 g770989 ( .a(n_9504), .b(n_9503), .o(n_9550) );
na02f80 g749861 ( .a(FE_OCP_RBN3012_n_31117), .b(n_31288), .o(n_31340) );
na02f80 g765962 ( .a(n_14670), .b(n_14633), .o(n_14727) );
na02f80 g776296 ( .a(n_4592), .b(n_4397), .o(n_4630) );
no02f80 g769700 ( .a(n_11285), .b(n_11284), .o(n_11357) );
in01f80 FE_RC_2124_0 ( .a(n_20836), .o(FE_RN_740_0) );
no02f80 g758794 ( .a(n_21587), .b(n_45081), .o(n_21617) );
ao12f80 g751364 ( .a(n_29010), .b(n_29388), .c(n_29006), .o(n_29460) );
no02f80 g752800 ( .a(n_27810), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_7_), .o(n_27880) );
ao12f80 g777027 ( .a(n_3556), .b(n_3557), .c(n_3388), .o(n_3583) );
in01f80 FE_RC_2051_0 ( .a(FE_RN_693_0), .o(n_26112) );
in01f80 newInst_3422 ( .a(newNet_2444), .o(newNet_3422) );
na02f80 g738596 ( .a(n_41499), .b(n_41462), .o(n_41500) );
in01f80 g752571 ( .a(n_27643), .o(n_27619) );
no02f80 g754523 ( .a(n_26511), .b(FE_OCPN928_n_26231), .o(n_26577) );
na02f80 g768491 ( .a(n_12336), .b(delay_add_ln22_unr8_stage4_stallmux_q_9_), .o(n_12398) );
no02f80 g765990 ( .a(n_14745), .b(n_14761), .o(n_14898) );
in01f80 FE_RC_2216_0 ( .a(n_32603), .o(FE_RN_800_0) );
oa22f80 g784425 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_2_), .c(n_36353), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_46237) );
no02f80 g780423 ( .a(n_847), .b(n_821), .o(n_1079) );
ao22s80 g781207 ( .a(n_90), .b(n_158), .c(n_85), .d(beta_26), .o(n_163) );
no02f80 g743914 ( .a(n_35916), .b(n_35783), .o(n_35954) );
no02f80 g775919 ( .a(n_6030), .b(FE_OCP_RBN2727_n_4219), .o(n_4991) );
in01f80 g775271 ( .a(delay_add_ln22_unr5_stage3_stallmux_q_13_), .o(n_7135) );
na02f80 g770570 ( .a(n_10102), .b(n_10016), .o(n_10277) );
ao22s80 FE_RC_1292_0 ( .a(n_9017), .b(n_8930), .c(n_8929), .d(n_9018), .o(n_9198) );
na02f80 g763682 ( .a(FE_OCP_RBN3707_n_16649), .b(n_16396), .o(n_16714) );
na02f80 g778202 ( .a(n_2795), .b(n_2794), .o(n_2906) );
in01f80 g756501 ( .a(n_23731), .o(n_23732) );
ao22s80 FE_RC_4269_0 ( .a(n_21745), .b(n_21709), .c(n_21685), .d(n_21768), .o(n_21874) );
in01f80 g767400 ( .a(n_13385), .o(n_14543) );
ao12f80 g754802 ( .a(n_26073), .b(n_26106), .c(n_26072), .o(n_26634) );
in01f80 g742742 ( .a(n_37407), .o(n_37408) );
na02f80 g750947 ( .a(n_28974), .b(n_28973), .o(n_28975) );
in01f80 g739771 ( .a(n_40509), .o(n_40510) );
in01f80 g762995 ( .a(n_17762), .o(n_17763) );
na02f80 FE_RC_2145_0 ( .a(FE_RN_550_0), .b(n_15142), .o(FE_RN_755_0) );
oa22f80 FE_RC_10_0 ( .a(FE_OCP_RBN2294_n_2438), .b(FE_OCP_RBN2379_n_3502), .c(FE_OCP_RBN2297_n_2438), .d(n_3502), .o(n_3018) );
in01f80 newInst_263 ( .a(newNet_262), .o(newNet_263) );
ao12f80 g746774 ( .a(FE_OCP_RBN2167_n_32892), .b(n_32959), .c(n_32991), .o(n_32997) );
in01f80 g755136 ( .a(n_25613), .o(n_25614) );
no03m80 FE_RC_1034_0 ( .a(n_33146), .b(n_32629), .c(n_33087), .o(n_33191) );
in01f80 newInst_482 ( .a(newNet_146), .o(newNet_482) );
no02f80 g746704 ( .a(n_33270), .b(n_33153), .o(n_33271) );
in01f80 FE_OFC738_n_22641 ( .a(FE_OFN734_n_22641), .o(FE_OFN738_n_22641) );
ao22s80 g778409 ( .a(n_2458), .b(n_2492), .c(n_2520), .d(n_2463), .o(n_2599) );
in01f80 g743303 ( .a(n_36739), .o(n_36740) );
no02f80 g765307 ( .a(n_15719), .b(n_15870), .o(n_16020) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_22_ ( .ck(newNet_2385), .d(n_36432), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_) );
in01f80 newInst_2118 ( .a(newNet_2117), .o(newNet_2118) );
na02f80 g749768 ( .a(n_31221), .b(n_31189), .o(n_31190) );
in01f80 newInst_3301 ( .a(newNet_1246), .o(newNet_3301) );
ao12f80 g779654 ( .a(n_1748), .b(n_1686), .c(delay_sub_ln23_0_unr2_stage2_stallmux_q_22_), .o(n_1798) );
oa12f80 g767510 ( .a(n_13223), .b(n_13222), .c(n_13221), .o(n_14733) );
na02f80 g771839 ( .a(n_9648), .b(n_9811), .o(n_9813) );
in01f80 g768591 ( .a(n_12314), .o(n_12315) );
in01f80 FE_OCP_RBC3732_n_31819 ( .a(FE_OCP_RBN3085_n_31819), .o(FE_OCP_RBN3732_n_31819) );
na02f80 g738331 ( .a(n_41818), .b(n_41817), .o(n_41819) );
oa12f80 g752972 ( .a(n_27762), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_5_), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_4_), .o(n_28204) );
in01f80 newInst_2514 ( .a(newNet_2513), .o(newNet_2514) );
na02f80 g737371 ( .a(n_42838), .b(n_42770), .o(n_42846) );
no02f80 g745405 ( .a(n_36049), .b(n_35240), .o(n_36123) );
na02f80 g760866 ( .a(n_19365), .b(n_18455), .o(n_19363) );
no02f80 g750806 ( .a(n_29118), .b(n_28645), .o(n_29164) );
in01f80 g746939 ( .a(n_32879), .o(n_32918) );
na02f80 g775061 ( .a(n_6070), .b(n_6111), .o(n_6159) );
in01f80 newInst_2068 ( .a(newNet_2067), .o(newNet_2068) );
no02f80 FE_RC_2427_0 ( .a(FE_RN_962_0), .b(FE_RN_963_0), .o(FE_RN_964_0) );
na02f80 g739450 ( .a(n_44775), .b(n_40581), .o(n_40928) );
oa12f80 g760519 ( .a(n_20133), .b(n_20450), .c(n_20178), .o(n_20516) );
in01f80 g772372 ( .a(n_8601), .o(n_8602) );
na02f80 g768090 ( .a(FE_OCPN860_n_12880), .b(n_12838), .o(n_13031) );
in01f80 FE_RC_2865_0 ( .a(n_33834), .o(FE_RN_1235_0) );
in01f80 g760177 ( .a(n_20660), .o(n_20661) );
oa12f80 g759438 ( .a(n_20916), .b(n_20915), .c(n_20914), .o(n_20970) );
no02f80 g778312 ( .a(n_2947), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_29_), .o(n_2835) );
in01f80 g763789 ( .a(n_18483), .o(n_16968) );
no02f80 g774832 ( .a(n_6251), .b(n_6304), .o(n_6305) );
in01f80 drc784748 ( .a(n_30633), .o(n_47233) );
in01f80 g760168 ( .a(n_21562), .o(n_21597) );
na02f80 g760353 ( .a(n_20835), .b(n_20810), .o(n_20811) );
in01f80 FE_OCP_RBC2628_n_14590 ( .a(FE_OCP_RBN2627_n_14590), .o(FE_OCP_RBN2628_n_14590) );
no02f80 g772784 ( .a(n_8154), .b(FE_OCP_RBN3453_FE_OCPN1240_n_7721), .o(n_8177) );
in01f80 g764830 ( .a(n_15625), .o(n_15626) );
in01f80 g741131 ( .a(n_39074), .o(n_39075) );
in01f80 g736941 ( .a(n_43256), .o(n_43257) );
in01f80 g772251 ( .a(n_8770), .o(n_8813) );
ao12f80 g747702 ( .a(n_33392), .b(n_33391), .c(n_33552), .o(n_33420) );
in01f80 g743543 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_22_), .o(n_36950) );
na02f80 g769754 ( .a(n_11196), .b(n_11228), .o(n_11312) );
na02f80 g773815 ( .a(n_7209), .b(n_7208), .o(n_7210) );
no02f80 g738573 ( .a(n_41687), .b(n_41527), .o(n_41568) );
ao12f80 g774387 ( .a(n_6742), .b(n_6789), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_12_), .o(n_6892) );
na02f80 g769670 ( .a(n_11245), .b(n_11210), .o(n_11320) );
in01f80 g773553 ( .a(n_7430), .o(n_7431) );
in01f80 newInst_3699 ( .a(newNet_3698), .o(newNet_3699) );
na02f80 g756537 ( .a(n_23563), .b(n_23562), .o(n_23586) );
no02f80 g754811 ( .a(n_26007), .b(n_25369), .o(n_26034) );
in01f80 newInst_3684 ( .a(newNet_3683), .o(newNet_3684) );
na02f80 g761436 ( .a(n_18799), .b(n_18710), .o(n_18832) );
in01f80 g754641 ( .a(n_27131), .o(n_27246) );
ao12f80 g772342 ( .a(n_8589), .b(n_8613), .c(n_8588), .o(n_9767) );
in01f80 newInst_3327 ( .a(newNet_2982), .o(newNet_3327) );
oa12f80 g766567 ( .a(n_13967), .b(n_14435), .c(n_14039), .o(n_14494) );
no02f80 g755055 ( .a(n_25556), .b(n_25535), .o(n_25585) );
na02f80 g777092 ( .a(n_3890), .b(n_3604), .o(n_3926) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_5_ ( .ck(newNet_2614), .d(n_21426), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_5_) );
oa22f80 FE_RC_1481_0 ( .a(n_32287), .b(FE_OCP_RBN3136_n_32380), .c(n_28336), .d(n_32380), .o(n_32467) );
in01f80 g750541 ( .a(n_29429), .o(n_29430) );
na02f80 g752123 ( .a(n_28061), .b(n_27965), .o(n_28119) );
in01f80 newInst_303 ( .a(newNet_145), .o(newNet_303) );
no02f80 g770125 ( .a(n_10755), .b(n_10803), .o(n_10898) );
no02f80 g736692 ( .a(n_43465), .b(n_43451), .o(n_43522) );
no02f80 g765356 ( .a(n_15039), .b(n_15109), .o(n_15191) );
no02f80 g770143 ( .a(n_44853), .b(n_10413), .o(n_10674) );
ao12f80 g784608 ( .a(n_42950), .b(n_42928), .c(n_42673), .o(n_46936) );
na02f80 FE_RC_2925_0 ( .a(n_27157), .b(FE_RN_565_0), .o(FE_RN_1274_0) );
na02f80 g771609 ( .a(n_10210), .b(n_11266), .o(n_10296) );
in01f80 g773517 ( .a(n_8303), .o(n_7484) );
in01f80 g763363 ( .a(n_17083), .o(n_17123) );
na02f80 g772626 ( .a(n_8319), .b(n_8364), .o(n_8437) );
in01f80 FE_OFC0_n_43918 ( .a(n_43918), .o(FE_OFN0_n_43918) );
no02f80 g745336 ( .a(n_35882), .b(n_35844), .o(n_35959) );
in01f80 g770549 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_6_), .o(n_10493) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_8_ ( .ck(newNet_539), .d(n_17476), .o(delay_xor_ln22_unr12_stage5_stallmux_q_8_) );
in01f80 g760730 ( .a(n_19658), .o(n_19695) );
ao12f80 g746459 ( .a(n_33454), .b(n_33453), .c(n_33452), .o(n_34122) );
in01f80 g766965 ( .a(FE_OCP_RBN2324_n_13616), .o(n_13656) );
in01f80 g772270 ( .a(n_8810), .o(n_8811) );
na02f80 g777718 ( .a(n_3339), .b(n_3359), .o(n_3428) );
in01f80 FE_OCP_RBC2549_n_44944 ( .a(n_44944), .o(FE_OCP_RBN2549_n_44944) );
ao12f80 g767918 ( .a(n_12742), .b(n_12741), .c(n_12740), .o(n_13118) );
in01f80 g769200 ( .a(n_12165), .o(n_12166) );
in01f80 newInst_3039 ( .a(newNet_3038), .o(newNet_3039) );
ms00f80 delay_sub_ln23_0_unr11_stage5_stallmux_q_reg ( .ck(newNet_1888), .d(n_16338), .o(n_44365) );
in01f80 FE_RC_2772_0 ( .a(n_9012), .o(FE_RN_1181_0) );
in01f80 FE_OCPC857_n_45697 ( .a(FE_OCPN867_n_45697), .o(FE_OCPN857_n_45697) );
no02f80 g756241 ( .a(n_24676), .b(n_24675), .o(n_24677) );
na02f80 g771952 ( .a(FE_OCP_RBN3552_n_44575), .b(n_9151), .o(n_9206) );
na02f80 g744132 ( .a(n_35571), .b(n_35613), .o(n_35614) );
in01f80 newInst_1877 ( .a(newNet_1876), .o(newNet_1877) );
in01f80 g779101 ( .a(n_2059), .o(n_2060) );
no02f80 g776589 ( .a(n_4434), .b(n_4433), .o(n_4582) );
in01f80 g770540 ( .a(n_10494), .o(n_10495) );
in01f80 g780913 ( .a(n_467), .o(n_482) );
in01f80 g765887 ( .a(n_14927), .o(n_14878) );
na02f80 g784598 ( .a(n_16197), .b(n_14524), .o(n_46421) );
oa22f80 FE_RC_3265_0 ( .a(n_20874), .b(FE_RN_1397_0), .c(n_20904), .d(FE_RN_1398_0), .o(n_21059) );
no02f80 g753447 ( .a(n_26987), .b(n_26985), .o(n_26986) );
no02f80 g739360 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_21_), .o(n_40786) );
in01f80 fopt783061 ( .a(n_44464), .o(n_44490) );
na02f80 g756331 ( .a(n_24478), .b(n_24065), .o(n_24588) );
in01f80 FE_OCP_RBC3566_n_29857 ( .a(FE_OCP_RBN3564_n_29857), .o(FE_OCP_RBN3566_n_29857) );
in01f80 g759299 ( .a(n_21153), .o(n_21154) );
in01f80 newInst_1799 ( .a(newNet_1798), .o(newNet_1799) );
na03f80 FE_RC_2250_0 ( .a(n_37251), .b(FE_RN_828_0), .c(FE_RN_823_0), .o(FE_RN_829_0) );
in01f80 g743201 ( .a(n_36928), .o(n_36929) );
na02f80 g772817 ( .a(n_8115), .b(n_8114), .o(n_8251) );
ao12f80 g741798 ( .a(n_38445), .b(n_38444), .c(n_38443), .o(n_38964) );
na02f80 g759347 ( .a(n_21116), .b(n_21063), .o(n_21176) );
na02f80 g775245 ( .a(n_5883), .b(n_5736), .o(n_5959) );
in01f80 FE_OCP_RBC1364_n_20412 ( .a(n_20412), .o(FE_OCP_RBN1364_n_20412) );
na02f80 g753935 ( .a(n_26178), .b(n_26130), .o(n_26226) );
no02f80 g759407 ( .a(n_20829), .b(FE_OCP_RBN1728_FE_RN_1583_0), .o(n_20855) );
in01f80 g777002 ( .a(n_4096), .o(n_4097) );
na02f80 g747186 ( .a(n_32736), .b(n_32735), .o(n_32797) );
in01f80 g738491 ( .a(n_41671), .o(n_41731) );
na02f80 g738301 ( .a(n_41836), .b(n_41835), .o(n_41837) );
na03f80 g768914 ( .a(n_11774), .b(n_11786), .c(n_11697), .o(n_11927) );
na02f80 g764371 ( .a(n_16285), .b(FE_OCPN3775_n_14730), .o(n_16401) );
na02f80 g740603 ( .a(n_39593), .b(n_45841), .o(n_39615) );
in01f80 g741791 ( .a(n_38421), .o(n_38448) );
oa12f80 g738351 ( .a(n_41449), .b(n_41551), .c(n_41399), .o(n_41818) );
na02f80 g746314 ( .a(n_33503), .b(delay_sub_ln23_0_unr21_stage8_stallmux_q), .o(n_33547) );
na02f80 g753830 ( .a(n_26429), .b(n_26428), .o(n_26518) );
oa12f80 g763653 ( .a(n_16828), .b(n_16829), .c(delay_sub_ln21_0_unr11_stage5_stallmux_q_0_), .o(n_18404) );
no02f80 g740891 ( .a(n_39307), .b(n_39269), .o(n_39373) );
ao22s80 FE_RC_4058_0 ( .a(FE_RN_1764_0), .b(n_26390), .c(FE_RN_1765_0), .d(n_26401), .o(n_26588) );
in01f80 g762421 ( .a(n_18023), .o(n_18024) );
no02f80 g752844 ( .a(n_27304), .b(n_27354), .o(n_27429) );
in01f80 g739798 ( .a(n_40484), .o(n_40485) );
in01f80 g765835 ( .a(n_14909), .o(n_14929) );
in01f80 g776958 ( .a(n_3681), .o(n_3655) );
in01f80 fopt783478 ( .a(n_45070), .o(n_45073) );
in01f80 g767719 ( .a(n_12713), .o(n_12745) );
oa12f80 g749582 ( .a(n_30408), .b(n_30407), .c(n_30406), .o(n_31448) );
ao12f80 g757916 ( .a(n_21921), .b(n_22110), .c(n_21922), .o(n_22169) );
na02f80 g739129 ( .a(n_41026), .b(n_40823), .o(n_41027) );
in01f80 newInst_1304 ( .a(newNet_1303), .o(newNet_1304) );
na02f80 FE_RC_2339_0 ( .a(FE_RN_894_0), .b(FE_RN_895_0), .o(n_19097) );
no02f80 g771856 ( .a(n_9219), .b(n_9218), .o(n_9325) );
na02f80 g756474 ( .a(n_23768), .b(n_23767), .o(n_23790) );
na02f80 g753226 ( .a(n_27207), .b(FE_OCPN1864_n_26171), .o(n_27383) );
in01f80 FE_RC_1924_0 ( .a(n_35235), .o(FE_RN_608_0) );
ao12f80 g756227 ( .a(n_24738), .b(n_24737), .c(n_24736), .o(n_25135) );
na02f80 g778932 ( .a(n_2159), .b(n_1968), .o(n_2222) );
in01f80 g758781 ( .a(n_22242), .o(n_22243) );
in01f80 g763413 ( .a(n_17213), .o(n_17214) );
in01f80 fopt783205 ( .a(FE_OCP_RBN2126_n_44734), .o(n_44735) );
in01f80 g762224 ( .a(n_18188), .o(n_18189) );
na02f80 g744259 ( .a(n_44180), .b(n_35613), .o(n_36134) );
ao22s80 g740953 ( .a(n_39138), .b(n_39228), .c(n_39137), .d(n_39229), .o(n_39822) );
in01f80 g752370 ( .a(delay_add_ln22_unr17_stage7_stallmux_q_25_), .o(n_28630) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_6_ ( .ck(newNet_2806), .d(n_10392), .o(delay_add_ln22_unr8_stage4_stallmux_q_6_) );
na02f80 g744990 ( .a(n_34833), .b(n_34452), .o(n_34906) );
ao22s80 FE_RC_3441_0 ( .a(n_20401), .b(n_20728), .c(n_20400), .d(n_20686), .o(n_20848) );
na02f80 g759517 ( .a(n_20961), .b(n_20960), .o(n_20962) );
no02f80 g765197 ( .a(n_16099), .b(n_16098), .o(n_16131) );
in01f80 newInst_1537 ( .a(newNet_1536), .o(newNet_1537) );
oa12f80 g784434 ( .a(n_46208), .b(n_46204), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .o(n_46246) );
no02f80 g781162 ( .a(n_183), .b(n_180), .o(n_199) );
in01f80 newInst_1259 ( .a(newNet_1258), .o(newNet_1259) );
na02f80 g751969 ( .a(n_28793), .b(n_28899), .o(n_29049) );
no02f80 g766418 ( .a(n_14127), .b(n_13437), .o(n_14131) );
in01f80 FE_OCP_RBC2349_n_38515 ( .a(n_38515), .o(FE_OCP_RBN2349_n_38515) );
na02f80 g763408 ( .a(n_16941), .b(n_16902), .o(n_17033) );
na02f80 g738754 ( .a(n_41564), .b(n_41199), .o(n_41729) );
in01f80 g744742 ( .a(n_35264), .o(n_35265) );
ao12f80 g751927 ( .a(n_28924), .b(n_28919), .c(n_28901), .o(n_29462) );
no02f80 FE_RC_3719_0 ( .a(FE_RN_1636_0), .b(n_5920), .o(n_46996) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_23_ ( .ck(newNet_2940), .d(n_6376), .o(delay_add_ln22_unr5_stage3_stallmux_q_23_) );
in01f80 g742895 ( .a(n_37288), .o(n_37077) );
in01f80 FE_OCP_DRV_C1582_n_35500 ( .a(FE_OCP_DRV_N1581_n_35500), .o(FE_OCP_DRV_N1582_n_35500) );
in01f80 fopt783962 ( .a(FE_OCP_RBN2121_n_45224), .o(n_45659) );
in01f80 g763927 ( .a(n_17155), .o(n_17304) );
in01f80 drc784123 ( .a(n_45873), .o(n_45874) );
ao12f80 g755194 ( .a(n_25608), .b(n_25607), .c(n_25606), .o(n_25745) );
oa12f80 g768319 ( .a(n_12313), .b(n_12519), .c(n_12262), .o(n_12553) );
na02f80 g754106 ( .a(n_26165), .b(n_23486), .o(n_26166) );
in01f80 g737910 ( .a(n_42283), .o(n_42258) );
na02f80 g750860 ( .a(n_29113), .b(n_30364), .o(n_29114) );
ao22s80 FE_RC_3432_0 ( .a(n_26305), .b(n_26137), .c(n_26304), .d(n_26138), .o(n_26440) );
na02f80 g768067 ( .a(n_12721), .b(n_12671), .o(n_12765) );
in01f80 newInst_793 ( .a(newNet_792), .o(newNet_793) );
no02f80 g756011 ( .a(n_25032), .b(n_25124), .o(n_25140) );
no02f80 g752228 ( .a(n_28539), .b(n_44046), .o(n_28589) );
in01f80 g766342 ( .a(n_14328), .o(n_15250) );
oa22f80 g784564 ( .a(FE_OFN800_n_46285), .b(n_11098), .c(FE_OCP_RBN3709_n_46337), .d(n_11055), .o(n_46385) );
na02f80 g747410 ( .a(n_32578), .b(n_32582), .o(n_32601) );
na02f80 g749875 ( .a(n_31311), .b(n_31371), .o(n_31569) );
na02f80 g763399 ( .a(n_16191), .b(FE_OCP_RBN3725_n_16975), .o(n_17323) );
no02f80 g741835 ( .a(n_38340), .b(n_38164), .o(n_38341) );
ms00f80 delay_sub_ln23_0_unr28_stage10_stallmux_q_reg ( .ck(newNet_1438), .d(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(delay_sub_ln23_0_unr28_stage10_stallmux_q) );
na02f80 g753208 ( .a(n_27207), .b(n_26113), .o(n_27425) );
oa12f80 g756880 ( .a(n_23867), .b(n_24188), .c(n_23810), .o(n_24733) );
na02f80 g771570 ( .a(n_8979), .b(n_8946), .o(n_9080) );
no02f80 g752050 ( .a(n_28711), .b(n_28710), .o(n_28712) );
no02f80 g776724 ( .a(n_4304), .b(n_4277), .o(n_4401) );
in01f80 g784708 ( .a(n_11308), .o(n_47183) );
in01f80 g739216 ( .a(n_40827), .o(n_40828) );
no02f80 g743465 ( .a(n_36629), .b(n_36750), .o(n_36630) );
na02f80 g753083 ( .a(n_27208), .b(n_27232), .o(n_27269) );
in01f80 newInst_72 ( .a(newNet_71), .o(newNet_72) );
na02f80 g767892 ( .a(n_12905), .b(n_12910), .o(n_12925) );
in01f80 newInst_2812 ( .a(newNet_2811), .o(newNet_2812) );
na02f80 g743424 ( .a(n_36667), .b(FE_OCPN1770_delay_sub_ln23_0_unr23_stage8_stallmux_q), .o(n_36732) );
in01f80 g747478 ( .a(n_32687), .o(n_32612) );
oa22f80 g780071 ( .a(n_1218), .b(n_1057), .c(n_1220), .d(n_1058), .o(n_1224) );
in01f80 newInst_315 ( .a(newNet_171), .o(newNet_315) );
na02f80 g781213 ( .a(n_104), .b(n_84), .o(n_105) );
in01f80 FE_OCP_RBC3620_n_15135 ( .a(n_15135), .o(FE_OCP_RBN3620_n_15135) );
in01f80 g773535 ( .a(n_7452), .o(n_7453) );
in01f80 g747497 ( .a(delay_xor_ln21_unr21_stage8_stallmux_q_1_), .o(n_32367) );
no02f80 g750726 ( .a(n_29194), .b(n_28766), .o(n_29240) );
in01f80 newInst_1228 ( .a(newNet_1227), .o(newNet_1228) );
in01f80 g773416 ( .a(n_7593), .o(n_8634) );
in01f80 g774322 ( .a(n_6577), .o(n_6578) );
in01f80 FE_RC_1063_0 ( .a(n_37426), .o(FE_RN_312_0) );
in01f80 FE_OCP_RBC1167_n_18949 ( .a(n_18949), .o(FE_OCP_RBN1167_n_18949) );
in01f80 g776561 ( .a(n_4515), .o(n_4516) );
na02f80 g738505 ( .a(FE_OCP_RBN2314_n_41420), .b(n_41290), .o(n_41699) );
in01f80 g736813 ( .a(n_43177), .o(n_43178) );
na02f80 g773835 ( .a(n_7103), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_11_), .o(n_7165) );
in01f80 FE_OCP_RBC3103_n_32163 ( .a(n_32163), .o(FE_OCP_RBN3103_n_32163) );
no02f80 g741861 ( .a(n_38410), .b(n_38409), .o(n_38411) );
no02f80 g736654 ( .a(n_43369), .b(n_43283), .o(n_43477) );
na02f80 g749737 ( .a(n_31190), .b(FE_OCP_RBN3009_n_31117), .o(n_31257) );
no02f80 g768016 ( .a(n_12614), .b(n_12497), .o(n_12653) );
in01f80 newInst_3609 ( .a(newNet_2950), .o(newNet_3609) );
na02f80 g767808 ( .a(n_13118), .b(n_13017), .o(n_13192) );
in01f80 newInst_82 ( .a(newNet_45), .o(newNet_82) );
no02f80 g738587 ( .a(n_41760), .b(n_41418), .o(n_41817) );
in01f80 FE_OCP_RBC2376_n_29480 ( .a(n_29480), .o(FE_OCP_RBN2376_n_29480) );
no02f80 g780219 ( .a(n_45817), .b(n_763), .o(n_1077) );
no02f80 g775126 ( .a(n_5926), .b(n_5925), .o(n_5947) );
in01f80 g753955 ( .a(n_26218), .o(n_26283) );
in01f80 newInst_1914 ( .a(newNet_1913), .o(newNet_1914) );
in01f80 FE_OCPC1493_n_23398 ( .a(n_23398), .o(FE_OCPN1493_n_23398) );
ao12f80 g766285 ( .a(n_14181), .b(n_14199), .c(n_14243), .o(n_14244) );
na02f80 g779086 ( .a(n_1988), .b(n_1833), .o(n_2043) );
in01f80 g740453 ( .a(n_39790), .o(n_39791) );
no02f80 g757848 ( .a(n_22319), .b(n_22002), .o(n_22391) );
no02f80 g761447 ( .a(n_20086), .b(n_19986), .o(n_20218) );
no02f80 g748086 ( .a(n_31968), .b(n_31951), .o(n_32024) );
na02f80 g775046 ( .a(n_6157), .b(n_6086), .o(n_6169) );
in01f80 fopt783397 ( .a(n_44996), .o(n_44995) );
no02f80 g760391 ( .a(n_20742), .b(n_20741), .o(n_20743) );
no02f80 g741952 ( .a(n_38119), .b(n_38166), .o(n_38219) );
oa22f80 g748055 ( .a(n_31876), .b(n_31838), .c(n_31877), .d(n_31839), .o(n_31955) );
in01f80 g761632 ( .a(n_18893), .o(n_18918) );
oa22f80 FE_RC_1386_0 ( .a(FE_OCPN3781_n_16440), .b(n_16596), .c(FE_OCPN3783_n_16463), .d(FE_OCP_RBN3051_n_16596), .o(n_16702) );
na02f80 g752191 ( .a(n_28085), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_2_), .o(n_28160) );
in01f80 g758690 ( .a(n_21964), .o(n_21944) );
in01f80 FE_OCP_RBC3331_n_44962 ( .a(n_44962), .o(FE_OCP_RBN3331_n_44962) );
na02f80 g759620 ( .a(n_20726), .b(n_20683), .o(n_20846) );
na02f80 FE_RC_83_0 ( .a(delay_xor_ln22_unr12_stage5_stallmux_q_5_), .b(n_45450), .o(FE_RN_24_0) );
no02f80 g737183 ( .a(n_42985), .b(n_42708), .o(n_42996) );
no02f80 g784406 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_18_), .o(n_46218) );
na02f80 g746352 ( .a(n_33475), .b(n_33164), .o(n_33492) );
in01f80 g768137 ( .a(n_12790), .o(n_12881) );
no02f80 g780055 ( .a(n_1230), .b(n_894), .o(n_1238) );
in01f80 g776739 ( .a(n_4081), .o(n_4082) );
no02f80 g744786 ( .a(n_35057), .b(n_30588), .o(n_35122) );
oa12f80 g738250 ( .a(n_41693), .b(n_41919), .c(n_41666), .o(n_41924) );
na02f80 g756793 ( .a(n_23380), .b(n_23253), .o(n_23422) );
no02f80 g774487 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_13_), .o(n_6878) );
no02f80 g744085 ( .a(n_35595), .b(FE_OCP_DRV_N1586_n_35594), .o(n_35622) );
ms00f80 delay_sub_ln23_0_unr20_stage7_stallmux_q_reg_17_ ( .ck(newNet_1628), .d(n_27165), .o(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_) );
in01f80 newInst_1038 ( .a(newNet_1037), .o(newNet_1038) );
oa12f80 g746516 ( .a(n_34810), .b(n_34809), .c(n_34299), .o(n_34811) );
in01f80 FE_OCP_RBC2310_n_29298 ( .a(FE_OCP_RBN2309_n_29298), .o(FE_OCP_RBN2310_n_29298) );
in01f80 g744033 ( .a(n_35669), .o(n_35700) );
in01f80 g768243 ( .a(n_12612), .o(n_12613) );
oa12f80 g777976 ( .a(n_2324), .b(n_3031), .c(n_2301), .o(n_3096) );
in01f80 g773625 ( .a(n_7702), .o(n_7728) );
no02f80 g774993 ( .a(n_6090), .b(n_6089), .o(n_6091) );
no02f80 g737530 ( .a(n_42494), .b(n_42435), .o(n_42495) );
in01f80 g752351 ( .a(n_27825), .o(n_27826) );
no02f80 g759936 ( .a(n_21406), .b(n_21481), .o(n_21446) );
in01f80 g748207 ( .a(n_32178), .o(n_32179) );
ao22s80 FE_RC_3323_0 ( .a(n_23714), .b(n_24140), .c(n_23715), .d(n_24139), .o(n_24222) );
no02f80 g756362 ( .a(n_24415), .b(n_24414), .o(n_24416) );
no02f80 g764693 ( .a(n_15768), .b(n_15523), .o(n_15770) );
in01f80 g739232 ( .a(n_41070), .o(n_41071) );
in01f80 newInst_2560 ( .a(newNet_2559), .o(newNet_2560) );
no02f80 g762236 ( .a(n_18163), .b(delay_add_ln22_unr11_stage5_stallmux_q_16_), .o(n_18215) );
ao12f80 g756426 ( .a(n_24239), .b(n_24238), .c(n_24237), .o(n_24299) );
in01f80 FE_OCP_RBC2963_n_26231 ( .a(FE_OCP_RBN2959_n_26231), .o(FE_OCP_RBN2963_n_26231) );
in01f80 g772910 ( .a(n_7966), .o(n_8063) );
in01f80 FE_RC_33_0 ( .a(n_6157), .o(FE_RN_7_0) );
in01f80 newInst_2807 ( .a(newNet_2204), .o(newNet_2807) );
oa22f80 g753463 ( .a(n_26788), .b(n_26647), .c(n_26732), .d(n_26648), .o(n_26810) );
in01f80 g739949 ( .a(n_40257), .o(n_40336) );
na02f80 g737034 ( .a(n_43082), .b(n_42597), .o(n_43113) );
no02f80 g737547 ( .a(n_42508), .b(n_42507), .o(n_42509) );
in01f80 g743164 ( .a(n_37084), .o(n_36981) );
no02f80 g760466 ( .a(n_20072), .b(n_18803), .o(n_20090) );
oa22f80 g739897 ( .a(FE_OCP_RBN3046_n_40231), .b(n_40362), .c(n_40258), .d(n_40361), .o(n_40428) );
na02f80 g747205 ( .a(n_32699), .b(n_32698), .o(n_32700) );
na02f80 g741660 ( .a(n_38521), .b(n_38375), .o(n_38541) );
in01f80 newInst_1072 ( .a(newNet_362), .o(newNet_1072) );
no02f80 g776709 ( .a(n_4335), .b(n_4446), .o(n_4573) );
in01f80 g743441 ( .a(n_37784), .o(n_37785) );
in01f80 g779161 ( .a(n_1940), .o(n_2445) );
na02f80 g751183 ( .a(n_29818), .b(n_29851), .o(n_29945) );
no02f80 g757598 ( .a(n_23276), .b(n_22695), .o(n_23277) );
in01f80 g759948 ( .a(n_21692), .o(n_21749) );
no02f80 g780470 ( .a(n_671), .b(n_707), .o(n_688) );
na02f80 g755360 ( .a(n_24911), .b(FE_OCP_RBN2404_n_24638), .o(n_24936) );
na02f80 g777653 ( .a(n_3428), .b(n_2913), .o(n_3433) );
na02f80 FE_RC_818_0 ( .a(n_8985), .b(FE_OCP_RBN2468_n_8767), .o(FE_RN_246_0) );
in01f80 g759994 ( .a(n_20632), .o(n_20633) );
na02f80 g759166 ( .a(n_21147), .b(n_21188), .o(n_21277) );
no02f80 g754323 ( .a(FE_OCP_RBN1199_n_25763), .b(n_23354), .o(n_25830) );
in01f80 g740990 ( .a(n_39106), .o(n_39135) );
no02f80 g757548 ( .a(FE_OCP_RBN3823_n_44061), .b(delay_xor_ln21_unr15_stage6_stallmux_q_3_), .o(n_22932) );
ao12f80 g746520 ( .a(n_34666), .b(n_34740), .c(n_34739), .o(n_34741) );
in01f80 g768047 ( .a(n_12918), .o(n_12884) );
ao22s80 g773396 ( .a(n_7539), .b(n_6922), .c(n_7538), .d(n_6923), .o(n_7945) );
in01f80 newInst_2754 ( .a(newNet_2753), .o(newNet_2754) );
na02f80 g746107 ( .a(n_33737), .b(n_33718), .o(n_33964) );
in01f80 g774208 ( .a(n_6598), .o(n_6599) );
no02f80 g740037 ( .a(n_39907), .b(n_39867), .o(n_39908) );
na02f80 g748920 ( .a(n_46101), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_20_), .o(n_32450) );
in01f80 g778691 ( .a(n_2590), .o(n_2591) );
na02f80 g764917 ( .a(n_16066), .b(n_15633), .o(n_16137) );
no02f80 g736621 ( .a(n_43565), .b(n_43316), .o(n_43566) );
in01f80 g743805 ( .a(n_36322), .o(n_36323) );
no02f80 g760199 ( .a(FE_OCPN1261_n_20242), .b(n_19414), .o(n_20567) );
in01f80 g740508 ( .a(n_39724), .o(n_39725) );
na02f80 g738985 ( .a(n_41205), .b(n_40856), .o(n_41220) );
na02f80 g763380 ( .a(FE_OCP_RBN3726_FE_RN_1787_0), .b(FE_OCPN3789_n_15708), .o(n_17329) );
no02f80 g770808 ( .a(n_10134), .b(n_10054), .o(n_10178) );
in01f80 FE_OCPC1433_n_30614 ( .a(n_30614), .o(FE_OCPN1433_n_30614) );
na02f80 g753481 ( .a(FE_OCP_RBN3034_n_26842), .b(n_26498), .o(n_26917) );
na02f80 g762197 ( .a(n_18167), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_14_), .o(n_18216) );
in01f80 g766080 ( .a(n_14664), .o(n_14610) );
ao12f80 g768482 ( .a(n_12358), .b(n_12357), .c(n_12356), .o(n_13074) );
na02f80 g740628 ( .a(n_39637), .b(n_39618), .o(n_39648) );
na02f80 g748902 ( .a(n_32393), .b(delay_sub_ln23_0_unr24_stage8_stallmux_q_2_), .o(n_32446) );
no02f80 g751586 ( .a(n_28447), .b(n_27669), .o(n_28577) );
no02f80 g747721 ( .a(n_32088), .b(n_32086), .o(n_32150) );
no04s80 g747177 ( .a(n_32706), .b(FE_OCP_RBN3369_n_32436), .c(n_32643), .d(n_32704), .o(n_32707) );
na02f80 g740385 ( .a(n_39803), .b(n_39878), .o(n_39851) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_19_ ( .ck(newNet_2957), .d(n_6297), .o(delay_add_ln22_unr5_stage3_stallmux_q_19_) );
in01f80 newInst_3371 ( .a(newNet_317), .o(newNet_3371) );
in01f80 newInst_2636 ( .a(newNet_2635), .o(newNet_2636) );
na02f80 g757898 ( .a(n_23083), .b(n_23117), .o(n_23118) );
ms00f80 delay_sub_ln23_0_unr8_stage4_stallmux_q_reg_3_ ( .ck(newNet_1076), .d(n_9653), .o(delay_sub_ln23_0_unr8_stage4_stallmux_q_3_) );
in01f80 g768428 ( .a(n_12497), .o(n_12498) );
in01f80 newInst_1059 ( .a(newNet_1058), .o(newNet_1059) );
in01f80 newInst_2770 ( .a(newNet_2769), .o(newNet_2770) );
na02f80 g775663 ( .a(n_47000), .b(n_5629), .o(n_5736) );
oa12f80 g762666 ( .a(n_17906), .b(n_17997), .c(n_17866), .o(n_18070) );
no02f80 FE_RC_2045_0 ( .a(FE_RN_683_0), .b(FE_RN_686_0), .o(FE_RN_687_0) );
no02f80 g750357 ( .a(n_29659), .b(n_29640), .o(n_29701) );
na02f80 g773456 ( .a(n_7527), .b(n_6830), .o(n_7565) );
oa12f80 g743814 ( .a(n_36336), .b(n_36335), .c(n_36334), .o(n_36387) );
oa22f80 FE_RC_1501_0 ( .a(n_25702), .b(n_25426), .c(n_25703), .d(n_25396), .o(n_25826) );
na02f80 g781238 ( .a(n_117), .b(n_44), .o(n_136) );
na02f80 g755725 ( .a(FE_OCP_RBN2338_n_24325), .b(n_23972), .o(n_24348) );
no02f80 g760219 ( .a(n_20249), .b(FE_OCP_RBN1688_n_18986), .o(n_20309) );
in01f80 g746068 ( .a(n_33975), .o(n_34003) );
in01f80 g765414 ( .a(n_15294), .o(n_15295) );
in01f80 g758190 ( .a(n_22498), .o(n_22499) );
in01f80 g767576 ( .a(n_13288), .o(n_13289) );
in01f80 newInst_1654 ( .a(newNet_1537), .o(newNet_1654) );
no02f80 g766129 ( .a(n_14450), .b(n_14416), .o(n_14451) );
na02f80 g779782 ( .a(n_1452), .b(delay_sub_ln23_0_unr2_stage2_stallmux_q_10_), .o(n_1441) );
oa12f80 g748023 ( .a(n_31751), .b(n_31777), .c(n_31612), .o(n_31881) );
no02f80 g752286 ( .a(n_27970), .b(n_27937), .o(n_27966) );
na02f80 g769192 ( .a(n_12016), .b(n_12050), .o(n_12544) );
na02f80 g761445 ( .a(n_19787), .b(n_19927), .o(n_19981) );
na02f80 g759775 ( .a(n_21517), .b(n_21516), .o(n_21995) );
in01f80 g773627 ( .a(n_7726), .o(n_7725) );
in01f80 FE_OFC784_delay_sub_ln23_0_unr15_stage6_stallmux_q ( .a(FE_OFN782_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q) );
no02f80 g766264 ( .a(n_14249), .b(n_13418), .o(n_14466) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_3_ ( .ck(newNet_955), .d(n_22704), .o(delay_xor_ln21_unr15_stage6_stallmux_q_3_) );
na02f80 g779777 ( .a(n_1780), .b(n_1381), .o(n_1396) );
no02f80 g743436 ( .a(n_36567), .b(n_36750), .o(n_36568) );
in01f80 FE_RC_2302_0 ( .a(n_25253), .o(FE_RN_870_0) );
ao12f80 g744472 ( .a(n_35393), .b(n_35467), .c(n_35418), .o(n_35503) );
na02f80 g749935 ( .a(n_29984), .b(n_29868), .o(n_29962) );
in01f80 g762257 ( .a(n_18619), .o(n_18698) );
in01f80 newInst_2657 ( .a(newNet_2301), .o(newNet_2657) );
na02f80 g752823 ( .a(n_27355), .b(n_27273), .o(n_27470) );
in01f80 g761375 ( .a(n_19712), .o(n_20011) );
in01f80 g740160 ( .a(n_39980), .o(n_40043) );
in01f80 g771711 ( .a(n_9275), .o(n_9392) );
na02f80 FE_RC_2457_0 ( .a(n_13697), .b(FE_RN_984_0), .o(FE_RN_985_0) );
in01f80 g736387 ( .a(n_43842), .o(n_43843) );
oa12f80 g784642 ( .a(n_18170), .b(n_18113), .c(n_17973), .o(n_46972) );
na02f80 g770586 ( .a(n_10498), .b(n_10461), .o(n_10462) );
in01f80 g753984 ( .a(n_26316), .o(n_26317) );
na02f80 g771197 ( .a(n_9452), .b(n_9408), .o(n_9538) );
in01f80 g745830 ( .a(n_34241), .o(n_34239) );
oa22f80 g739777 ( .a(n_40448), .b(n_40311), .c(n_40449), .d(n_40312), .o(n_40489) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_18_ ( .ck(newNet_2480), .d(n_32262), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_18_) );
na02f80 FE_RC_3637_0 ( .a(FE_RN_1595_0), .b(n_31466), .o(n_31751) );
oa22f80 g753167 ( .a(n_27287), .b(FE_OCP_RBN1200_n_25763), .c(n_27377), .d(FE_OCP_RBN1201_n_25763), .o(n_27542) );
in01f80 newInst_3394 ( .a(newNet_3393), .o(newNet_3394) );
na02f80 g741606 ( .a(n_38587), .b(FE_OCP_RBN2452_n_38537), .o(n_38603) );
in01f80 newInst_3045 ( .a(newNet_1415), .o(newNet_3045) );
ms00f80 delay_sub_ln21_0_unr8_stage4_stallmux_q_reg_16_ ( .ck(newNet_2013), .d(n_11307), .o(delay_sub_ln21_0_unr8_stage4_stallmux_q_16_) );
in01f80 g765857 ( .a(n_14862), .o(n_14884) );
in01f80 g775108 ( .a(n_6077), .o(n_6092) );
in01f80 FE_OCP_RBC1359_FE_RN_677_0 ( .a(FE_RN_677_0), .o(FE_OCP_RBN1359_FE_RN_677_0) );
ao12f80 g751747 ( .a(n_29047), .b(n_28989), .c(n_28919), .o(n_29048) );
in01f80 newInst_954 ( .a(newNet_953), .o(newNet_954) );
na02f80 g768507 ( .a(n_45659), .b(delay_xor_ln22_unr9_stage4_stallmux_q_22_), .o(n_12406) );
ms00f80 delay_xor_ln21_unr12_stage5_stallmux_q_reg_9_ ( .ck(newNet_990), .d(n_17567), .o(delay_xor_ln21_unr12_stage5_stallmux_q_9_) );
no02f80 g767565 ( .a(n_12978), .b(n_12941), .o(n_13146) );
no02f80 g778769 ( .a(n_2272), .b(n_2313), .o(n_2328) );
in01f80 g761488 ( .a(n_19849), .o(n_19824) );
na02f80 FE_RC_3159_0 ( .a(FE_RN_1400_0), .b(n_17417), .o(n_17523) );
in01f80 FE_OCP_RBC3416_n_12739 ( .a(FE_OCP_RBN3413_n_12739), .o(FE_OCP_RBN3416_n_12739) );
na02f80 g750962 ( .a(n_30231), .b(n_30162), .o(n_30232) );
in01f80 g780062 ( .a(n_1231), .o(n_1235) );
ao12f80 g747169 ( .a(n_33891), .b(n_33890), .c(n_33889), .o(n_34523) );
in01f80 g746975 ( .a(n_32957), .o(n_32958) );
ao12f80 g774064 ( .a(n_6711), .b(n_6729), .c(n_6710), .o(n_6860) );
in01f80 g773440 ( .a(n_7678), .o(n_7737) );
oa12f80 g750154 ( .a(n_30128), .b(n_30835), .c(n_30091), .o(n_30921) );
in01f80 g763851 ( .a(n_16726), .o(n_16748) );
na02f80 g761263 ( .a(n_19910), .b(n_19909), .o(n_19911) );
oa12f80 g776858 ( .a(n_4208), .b(n_4209), .c(n_4037), .o(n_4204) );
ms00f80 delay_xor_ln21_unr9_stage4_stallmux_q_reg_14_ ( .ck(newNet_659), .d(n_46359), .o(delay_xor_ln21_unr9_stage4_stallmux_q_14_) );
in01f80 newInst_2624 ( .a(newNet_1296), .o(newNet_2624) );
in01f80 g774723 ( .a(n_6382), .o(n_6383) );
no02f80 FE_RC_1120_0 ( .a(FE_RN_336_0), .b(FE_RN_337_0), .o(FE_RN_338_0) );
oa22f80 FE_RC_3827_0 ( .a(n_24059), .b(n_27726), .c(n_27796), .d(n_27704), .o(n_27748) );
in01f80 g765322 ( .a(n_15302), .o(n_15771) );
no02f80 g755233 ( .a(n_25039), .b(n_25037), .o(n_25097) );
in01f80 g745146 ( .a(n_35749), .o(n_34660) );
no02f80 g743084 ( .a(delay_add_ln22_unr23_stage9_stallmux_q_6_), .b(delay_sub_ln22_unr24_stage9_stallmux_q_6_), .o(n_36989) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_15_ ( .ck(newNet_2404), .d(n_36396), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_15_) );
na02f80 g765159 ( .a(n_15930), .b(n_15835), .o(n_15931) );
na02f80 g767238 ( .a(n_13535), .b(n_13530), .o(n_13531) );
no03m80 FE_RC_2548_0 ( .a(n_37154), .b(n_37311), .c(n_37374), .o(n_37451) );
oa12f80 g778220 ( .a(n_2690), .b(n_2689), .c(n_2688), .o(n_4435) );
in01f80 g779029 ( .a(n_2141), .o(n_2142) );
in01f80 FE_OCPC1755_n_16923 ( .a(FE_OCP_RBN3727_FE_RN_1787_0), .o(FE_OCPN1755_n_16923) );
in01f80 newInst_178 ( .a(newNet_72), .o(newNet_178) );
in01f80 g741520 ( .a(n_38705), .o(n_38706) );
na02f80 g757748 ( .a(n_23155), .b(n_23154), .o(n_23156) );
no02f80 g756343 ( .a(n_23929), .b(n_23600), .o(n_24000) );
no02f80 g776979 ( .a(n_4049), .b(n_4121), .o(n_4122) );
in01f80 g754302 ( .a(n_25925), .o(n_25926) );
no02f80 g759059 ( .a(n_21466), .b(n_45080), .o(n_21495) );
in01f80 fopt782972 ( .a(FE_OCP_RBN1297_n_30451), .o(n_44437) );
na02f80 FE_RC_3751_0 ( .a(FE_RN_1645_0), .b(FE_RN_1646_0), .o(FE_RN_1647_0) );
na02f80 g764787 ( .a(n_15692), .b(n_14452), .o(n_15763) );
ao12f80 g770516 ( .a(n_9651), .b(n_10527), .c(n_9730), .o(n_10577) );
in01f80 FE_OCP_RBC3515_n_8498 ( .a(n_8498), .o(FE_OCP_RBN3515_n_8498) );
in01f80 newInst_1499 ( .a(newNet_1498), .o(newNet_1499) );
no02f80 g779632 ( .a(n_1752), .b(n_1801), .o(n_2134) );
na02f80 g747435 ( .a(n_32592), .b(n_32632), .o(n_32647) );
no02f80 g747378 ( .a(n_32661), .b(delay_add_ln22_unr20_stage8_stallmux_q_0_), .o(n_32662) );
oa12f80 g767299 ( .a(n_13676), .b(n_13675), .c(n_13674), .o(n_14170) );
na02f80 g749355 ( .a(n_30541), .b(n_27014), .o(n_30566) );
in01f80 g749859 ( .a(n_31279), .o(n_31339) );
in01f80 g765256 ( .a(n_15601), .o(n_15602) );
na02f80 g751035 ( .a(n_29805), .b(n_29804), .o(n_29806) );
na02f80 g762187 ( .a(n_18161), .b(delay_add_ln22_unr11_stage5_stallmux_q_17_), .o(n_18220) );
na02f80 g758907 ( .a(n_21292), .b(n_21329), .o(n_21476) );
in01f80 g745201 ( .a(n_34594), .o(n_34595) );
in01f80 g756832 ( .a(n_23956), .o(n_23957) );
na02f80 g745574 ( .a(n_34297), .b(FE_OCPN3749_n_34296), .o(n_34348) );
ao12f80 g757871 ( .a(FE_OFN735_n_22641), .b(n_23119), .c(n_23056), .o(n_23120) );
in01f80 g763840 ( .a(n_16669), .o(n_16670) );
in01f80 newInst_2791 ( .a(newNet_612), .o(newNet_2791) );
na02f80 g741240 ( .a(FE_OCP_RBN2635_n_38806), .b(n_38433), .o(n_38880) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_15_ ( .ck(newNet_1760), .d(n_22245), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_15_) );
na02f80 g745599 ( .a(n_34297), .b(n_33616), .o(n_34374) );
no02f80 g757253 ( .a(n_23137), .b(delay_add_ln22_unr14_stage6_stallmux_q_5_), .o(n_23170) );
na02f80 g766270 ( .a(FE_OCP_RBN2482_n_14326), .b(FE_OCP_RBN3535_n_13765), .o(n_14409) );
na02f80 g775000 ( .a(n_5924), .b(n_5965), .o(n_6102) );
ao12f80 FE_RC_2848_0 ( .a(FE_RN_1225_0), .b(FE_RN_1226_0), .c(n_38747), .o(n_38780) );
in01f80 g769274 ( .a(n_11459), .o(n_11514) );
in01f80 FE_RC_793_0 ( .a(n_41434), .o(FE_RN_241_0) );
in01f80 g739387 ( .a(n_40787), .o(n_40688) );
no02f80 g780513 ( .a(n_819), .b(n_818), .o(n_820) );
na02f80 g772684 ( .a(n_8238), .b(FE_OCP_RBN2337_n_8269), .o(n_8299) );
na03f80 FE_RC_757_0 ( .a(n_11603), .b(n_11599), .c(n_11569), .o(n_11777) );
in01f80 g751412 ( .a(n_28610), .o(n_28652) );
in01f80 g751138 ( .a(n_30587), .o(n_30612) );
oa22f80 g758870 ( .a(n_22119), .b(n_21564), .c(n_22056), .d(n_21565), .o(n_22144) );
na02f80 g777257 ( .a(n_3533), .b(n_2771), .o(n_3518) );
in01f80 newInst_2981 ( .a(newNet_1220), .o(newNet_2981) );
no02f80 g776669 ( .a(n_4278), .b(n_4304), .o(n_4572) );
in01f80 g749046 ( .a(n_31023), .o(n_31024) );
in01f80 g747190 ( .a(n_32774), .o(n_32734) );
na02f80 g745942 ( .a(n_34088), .b(n_34087), .o(n_34089) );
na02f80 g778438 ( .a(FE_OCP_RBN2286_n_2433), .b(n_2858), .o(n_2470) );
no02f80 g738404 ( .a(n_41642), .b(n_41587), .o(n_42095) );
no02f80 g753531 ( .a(n_26821), .b(n_26820), .o(n_26837) );
in01f80 newInst_1951 ( .a(newNet_1950), .o(newNet_1951) );
in01f80 g775224 ( .a(n_5996), .o(n_6017) );
oa12f80 g772769 ( .a(n_8126), .b(n_8125), .c(n_8124), .o(n_9784) );
in01f80 FE_RC_3853_0 ( .a(n_20123), .o(n_20159) );
no02f80 g759734 ( .a(n_21375), .b(n_21336), .o(n_21410) );
in01f80 FE_RC_2154_0 ( .a(n_15175), .o(FE_RN_761_0) );
ms00f80 delay_add_ln22_unr17_stage7_stallmux_q_reg_23_ ( .ck(newNet_3412), .d(n_27726), .o(delay_add_ln22_unr17_stage7_stallmux_q_23_) );
no02f80 g747246 ( .a(n_32667), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_3_), .o(n_32695) );
no02f80 g745985 ( .a(n_34034), .b(n_34011), .o(n_34086) );
in01f80 g739839 ( .a(n_40442), .o(n_40443) );
in01f80 g769653 ( .a(n_11323), .o(n_11324) );
in01f80 g740850 ( .a(n_39493), .o(n_39430) );
no02f80 g750982 ( .a(n_30127), .b(n_30088), .o(n_30128) );
in01f80 g762296 ( .a(n_18138), .o(n_18095) );
na02f80 g773028 ( .a(n_7703), .b(n_7702), .o(n_7704) );
na02f80 g738299 ( .a(n_41888), .b(n_41594), .o(n_41801) );
in01f80 FE_OCPC1034_n_28420 ( .a(FE_OCPN1033_n_28420), .o(FE_OCPN1034_n_28420) );
in01f80 FE_RC_1335_0 ( .a(n_5218), .o(FE_RN_397_0) );
in01f80 g749288 ( .a(n_30771), .o(n_30737) );
no02f80 g745125 ( .a(n_34767), .b(n_34514), .o(n_34897) );
na02f80 g736714 ( .a(n_43314), .b(n_43230), .o(n_43404) );
in01f80 g754508 ( .a(n_26829), .o(n_26830) );
no02f80 g744704 ( .a(n_35269), .b(n_33640), .o(n_35379) );
in01f80 fopt782841 ( .a(n_44267), .o(n_44268) );
in01f80 g754142 ( .a(n_26059), .o(n_26060) );
na02f80 g767749 ( .a(n_13069), .b(n_12254), .o(n_13777) );
in01f80 g758471 ( .a(n_23271), .o(n_26054) );
in01f80 g773590 ( .a(n_7447), .o(n_7448) );
in01f80 g738372 ( .a(n_41792), .o(n_41732) );
na02f80 g755030 ( .a(n_25800), .b(n_25799), .o(n_25801) );
no02f80 g775130 ( .a(n_5732), .b(n_4875), .o(n_5760) );
in01f80 g745569 ( .a(n_34743), .o(n_34744) );
ms00f80 delay_add_ln22_unr11_stage5_stallmux_q_reg_9_ ( .ck(newNet_3574), .d(n_16106), .o(delay_add_ln22_unr11_stage5_stallmux_q_9_) );
in01f80 FE_OCPC1047_n_24819 ( .a(n_24819), .o(FE_OCPN1047_n_24819) );
in01f80 g759459 ( .a(n_20995), .o(n_21030) );
no02f80 FE_RC_4000_0 ( .a(FE_RN_1735_0), .b(n_29967), .o(FE_RN_1734_0) );
in01f80 g748673 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_4_), .o(n_32670) );
no02f80 g754894 ( .a(FE_OCPN985_n_25210), .b(n_24116), .o(n_25331) );
oa12f80 g737282 ( .a(n_42299), .b(n_42842), .c(n_42297), .o(n_42888) );
ao12f80 g773600 ( .a(n_7375), .b(n_7381), .c(n_7374), .o(n_7439) );
in01f80 newInst_3308 ( .a(newNet_3307), .o(newNet_3308) );
in01f80 g747316 ( .a(n_32554), .o(n_32790) );
na02f80 FE_RC_3902_0 ( .a(FE_RN_1281_0), .b(FE_RN_1695_0), .o(n_29778) );
no02f80 g769187 ( .a(n_11686), .b(n_11630), .o(n_11648) );
ao12f80 g739093 ( .a(n_41059), .b(n_41058), .c(n_41057), .o(n_41433) );
ao12f80 g752163 ( .a(n_28587), .b(n_28586), .c(n_28585), .o(n_28837) );
no02f80 g743551 ( .a(n_36543), .b(n_36750), .o(n_36579) );
na02f80 g760924 ( .a(n_19378), .b(n_18010), .o(n_19425) );
no02f80 g771941 ( .a(FE_OCP_RBN2514_n_8739), .b(n_8679), .o(n_8800) );
in01f80 g736975 ( .a(n_43357), .o(n_43341) );
na02f80 g744044 ( .a(n_44223), .b(n_34712), .o(n_36303) );
in01f80 newInst_3663 ( .a(newNet_3662), .o(newNet_3663) );
oa12f80 g784796 ( .a(n_44875), .b(n_38269), .c(n_37935), .o(n_47336) );
in01f80 FE_OCPC1232_n_42201 ( .a(FE_OCPN1230_n_42201), .o(FE_OCPN1232_n_42201) );
no02f80 g777632 ( .a(n_3598), .b(FE_OCPN848_n_3597), .o(n_3648) );
na02f80 g743379 ( .a(n_36594), .b(n_36750), .o(n_36595) );
na02f80 g741463 ( .a(n_44166), .b(n_38729), .o(n_38793) );
in01f80 newInst_2382 ( .a(newNet_1392), .o(newNet_2382) );
in01f80 FE_OCP_RBC2370_n_38545 ( .a(FE_OCP_RBN2369_n_38545), .o(FE_OCP_RBN2370_n_38545) );
no02f80 g776777 ( .a(n_3967), .b(n_4061), .o(n_4110) );
in01f80 g768335 ( .a(n_12533), .o(n_12534) );
in01f80 g770020 ( .a(n_10878), .o(n_10910) );
in01f80 newInst_447 ( .a(newNet_446), .o(newNet_447) );
in01f80 g751835 ( .a(n_28265), .o(n_28266) );
na02f80 g759927 ( .a(FE_OCP_RBN3678_n_21051), .b(n_21405), .o(n_21516) );
in01f80 g753113 ( .a(n_27224), .o(n_27225) );
in01f80 newInst_2590 ( .a(newNet_774), .o(newNet_2590) );
no02f80 g758254 ( .a(FE_OCP_RBN2045_delay_sub_ln23_unr17_stage6_stallmux_q_1_), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_2_), .o(n_22649) );
na02f80 FE_RC_2765_0 ( .a(FE_OCPN1424_delay_sub_ln23_0_unr21_stage8_stallmux_q), .b(n_33872), .o(FE_RN_1178_0) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_19_ ( .ck(newNet_3537), .d(n_22715), .o(delay_add_ln22_unr14_stage6_stallmux_q_19_) );
na02f80 g766131 ( .a(n_14484), .b(n_14475), .o(n_14517) );
in01f80 FE_OCP_RBC3850_n_20290 ( .a(n_20290), .o(FE_OCP_RBN3850_n_20290) );
no02f80 g757962 ( .a(n_22950), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_27_), .o(n_23007) );
in01f80 FE_OCPC3790_n_36069 ( .a(n_36069), .o(FE_OCPN3790_n_36069) );
in01f80 newInst_2287 ( .a(newNet_2286), .o(newNet_2287) );
oa22f80 FE_RC_4270_0 ( .a(n_22490), .b(n_22661), .c(n_22624), .d(n_22491), .o(n_22818) );
no02f80 g776289 ( .a(n_4697), .b(n_4200), .o(n_4698) );
na02f80 g738186 ( .a(n_41974), .b(n_41862), .o(n_42003) );
no02f80 g765902 ( .a(n_14816), .b(n_14795), .o(n_14874) );
na02f80 g765508 ( .a(n_15719), .b(n_15718), .o(n_15837) );
no02f80 g771818 ( .a(n_9876), .b(n_9825), .o(n_9877) );
in01f80 g765997 ( .a(n_15086), .o(n_15087) );
na02f80 g765084 ( .a(n_15347), .b(n_14419), .o(n_15348) );
ao12f80 g764181 ( .a(n_16173), .b(n_16824), .c(n_16255), .o(n_16850) );
no02f80 g737753 ( .a(n_42368), .b(n_42274), .o(n_42329) );
na02f80 g767033 ( .a(FE_OCP_RBN3534_n_13765), .b(n_13501), .o(n_13966) );
na02f80 g739075 ( .a(n_41082), .b(n_40893), .o(n_41128) );
no02f80 g778725 ( .a(n_45903), .b(n_2218), .o(n_2219) );
na02f80 g738267 ( .a(n_41846), .b(n_41845), .o(n_41847) );
na02f80 FE_RC_2778_0 ( .a(FE_RN_1183_0), .b(FE_RN_1185_0), .o(n_38421) );
ms00f80 sin_out_reg_26_ ( .ck(newNet_41), .d(n_43915), .o(sin_out_26) );
no02f80 g740967 ( .a(n_39313), .b(n_39108), .o(n_39215) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_18_ ( .ck(newNet_3540), .d(n_22631), .o(delay_add_ln22_unr14_stage6_stallmux_q_18_) );
in01f80 g774792 ( .a(n_6295), .o(n_6291) );
na02f80 g777053 ( .a(n_3903), .b(delay_sub_ln23_0_unr1_stage2_stallmux_q_0_), .o(n_3904) );
na02f80 FE_RC_674_0 ( .a(FE_RN_215_0), .b(n_28292), .o(n_28348) );
na02f80 g772405 ( .a(n_8410), .b(FE_OCP_RBN3466_n_7886), .o(n_8477) );
na02f80 g777197 ( .a(n_3782), .b(n_3693), .o(n_3835) );
no02f80 g749180 ( .a(n_32114), .b(n_31512), .o(n_32205) );
in01f80 g768726 ( .a(n_12247), .o(n_12942) );
in01f80 newInst_1864 ( .a(newNet_1863), .o(newNet_1864) );
in01f80 newInst_1558 ( .a(newNet_692), .o(newNet_1558) );
ao22s80 g780343 ( .a(n_824), .b(n_1203), .c(n_823), .d(FE_OFN761_n_45813), .o(n_924) );
oa12f80 g749814 ( .a(n_31340), .b(FE_OCP_RBN3012_n_31117), .c(n_31288), .o(n_31619) );
in01f80 g767145 ( .a(n_14524), .o(n_14618) );
in01f80 FE_OCPC999_n_19311 ( .a(FE_OCP_RBN1347_n_19270), .o(FE_OCPN999_n_19311) );
na02f80 g763943 ( .a(n_16570), .b(n_16441), .o(n_16590) );
no02f80 g773615 ( .a(n_7376), .b(delay_sub_ln21_0_unr5_stage3_stallmux_q_19_), .o(n_7395) );
in01f80 g751968 ( .a(n_29049), .o(n_28921) );
in01f80 newInst_2628 ( .a(newNet_2627), .o(newNet_2628) );
in01f80 newInst_1521 ( .a(newNet_695), .o(newNet_1521) );
in01f80 newInst_1451 ( .a(newNet_1311), .o(newNet_1451) );
in01f80 g778348 ( .a(n_2535), .o(n_2536) );
no02f80 g765504 ( .a(n_15719), .b(n_15779), .o(n_15876) );
ao12f80 g742550 ( .a(n_37124), .b(n_37446), .c(n_37258), .o(n_37494) );
ao22s80 FE_RC_1597_0 ( .a(FE_OCP_RBN2728_n_4219), .b(n_5988), .c(FE_OCP_RBN2727_n_4219), .d(n_4751), .o(n_4922) );
na02f80 g756607 ( .a(n_23581), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_18_), .o(n_23683) );
no02f80 g771791 ( .a(n_9263), .b(n_9218), .o(n_9482) );
in01f80 g736966 ( .a(n_43303), .o(n_43304) );
na02f80 FE_RC_2859_0 ( .a(FE_RN_1231_0), .b(n_10503), .o(FE_RN_1232_0) );
in01f80 g767107 ( .a(n_14758), .o(n_14210) );
in01f80 g747812 ( .a(n_33413), .o(n_33414) );
in01f80 g762411 ( .a(n_19400), .o(n_18607) );
in01f80 FE_RC_1639_0 ( .a(n_23067), .o(FE_RN_457_0) );
na02f80 g761382 ( .a(n_18900), .b(n_18876), .o(n_18981) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_7_ ( .ck(newNet_3274), .d(n_31405), .o(delay_add_ln22_unr20_stage8_stallmux_q_7_) );
in01f80 newInst_2901 ( .a(newNet_2399), .o(newNet_2901) );
in01f80 g754749 ( .a(n_25404), .o(n_25405) );
in01f80 g745116 ( .a(n_35665), .o(n_34726) );
in01f80 g748171 ( .a(n_32208), .o(n_32209) );
na02f80 g744898 ( .a(FE_OCP_RBN2710_n_35075), .b(n_30546), .o(n_35115) );
in01f80 FE_RC_4235_0 ( .a(FE_OFN737_n_22641), .o(FE_RN_1860_0) );
in01f80 g746020 ( .a(n_35241), .o(n_35299) );
oa12f80 g738937 ( .a(n_41239), .b(n_41238), .c(n_41237), .o(n_41290) );
in01f80 FE_RC_214_0 ( .a(n_12492), .o(FE_RN_70_0) );
in01f80 g766948 ( .a(n_14345), .o(n_14298) );
in01f80 g777645 ( .a(n_3400), .o(n_3418) );
in01f80 g740776 ( .a(n_39561), .o(n_39978) );
na02f80 FE_RC_1781_0 ( .a(FE_RN_519_0), .b(n_1979), .o(n_2318) );
no02f80 g749416 ( .a(n_30579), .b(n_30244), .o(n_30623) );
oa22f80 FE_RC_1595_0 ( .a(n_4452), .b(n_4531), .c(n_4451), .d(n_4530), .o(n_4751) );
oa22f80 g763334 ( .a(n_17128), .b(FE_OFN767_n_15670), .c(n_17061), .d(n_16339), .o(n_17224) );
no02f80 g754536 ( .a(n_26235), .b(n_26234), .o(n_26236) );
ao12f80 g762115 ( .a(n_18499), .b(n_18703), .c(n_18701), .o(n_18780) );
no02f80 g776028 ( .a(FE_OCPN960_n_3951), .b(n_4692), .o(n_4749) );
na02f80 g744102 ( .a(n_35819), .b(FE_OCP_RBN2902_n_44174), .o(n_36034) );
no02f80 g741974 ( .a(n_38056), .b(FE_OCPN1239_n_37945), .o(n_38110) );
in01f80 g766864 ( .a(n_13629), .o(n_13630) );
in01f80 g748763 ( .a(n_31356), .o(n_31377) );
in01f80 FE_OCP_RBC1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_ ( .a(delay_sub_ln23_0_unr5_stage3_stallmux_q_31_), .o(FE_OCP_RBN1984_delay_sub_ln23_0_unr5_stage3_stallmux_q_31_) );
in01f80 g769372 ( .a(n_12077), .o(n_12046) );
in01f80 newInst_813 ( .a(newNet_812), .o(newNet_813) );
na02f80 g762649 ( .a(n_18020), .b(n_18018), .o(n_18019) );
oa12f80 g778049 ( .a(n_2961), .b(n_2960), .c(n_2959), .o(n_4333) );
na02f80 g744608 ( .a(n_35316), .b(n_35315), .o(n_35330) );
in01f80 g751627 ( .a(FE_OCPN1030_n_28423), .o(n_28424) );
no02f80 g747482 ( .a(n_32591), .b(n_44962), .o(n_32620) );
ao22s80 g756383 ( .a(n_23826), .b(n_23596), .c(n_23777), .d(n_23595), .o(n_23887) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_2_ ( .ck(newNet_3119), .d(n_39855), .o(delay_add_ln22_unr27_stage10_stallmux_q_2_) );
oa12f80 g744564 ( .a(n_35381), .b(n_35380), .c(n_35379), .o(n_35409) );
in01f80 g773707 ( .a(n_7268), .o(n_7269) );
na02f80 g742144 ( .a(FE_OCP_RBN2255_n_37844), .b(n_37394), .o(n_37956) );
in01f80 g774505 ( .a(n_6756), .o(n_6721) );
in01f80 g769270 ( .a(n_11458), .o(n_11657) );
no02f80 g752783 ( .a(n_28109), .b(n_28108), .o(n_28110) );
in01f80 g754979 ( .a(n_25504), .o(n_25505) );
in01f80 g744376 ( .a(n_46213), .o(n_36810) );
na02f80 g740363 ( .a(n_39803), .b(n_40202), .o(n_39835) );
no02f80 g766595 ( .a(n_13988), .b(n_13785), .o(n_13989) );
na02f80 g744097 ( .a(n_35614), .b(n_44174), .o(n_35691) );
in01f80 g742475 ( .a(n_37755), .o(n_37689) );
in01f80 FE_OCP_RBC3212_n_44365 ( .a(FE_OCP_RBN3213_n_44365), .o(FE_OCP_RBN3212_n_44365) );
in01f80 g744942 ( .a(n_36405), .o(n_36406) );
in01f80 FE_OFC830_n_2540 ( .a(n_2540), .o(FE_OFN830_n_2540) );
in01f80 FE_RC_3700_0 ( .a(n_2764), .o(FE_RN_1628_0) );
in01f80 g737868 ( .a(n_42194), .o(n_42195) );
na02f80 g752505 ( .a(n_27712), .b(n_27710), .o(n_27711) );
oa12f80 g760436 ( .a(n_20085), .b(n_20624), .c(n_20112), .o(n_20701) );
ao12f80 g756789 ( .a(n_24355), .b(n_24076), .c(n_24059), .o(n_24815) );
in01f80 g764506 ( .a(n_16266), .o(n_16314) );
in01f80 g751229 ( .a(n_30156), .o(n_30303) );
na02f80 g756464 ( .a(n_23883), .b(n_23819), .o(n_23925) );
in01f80 g780680 ( .a(n_663), .o(n_666) );
na02f80 g778958 ( .a(n_2232), .b(n_2231), .o(n_2247) );
ao22s80 FE_RC_1416_0 ( .a(n_5918), .b(n_5939), .c(n_5917), .d(n_5938), .o(n_6034) );
na02f80 FE_RC_3014_0 ( .a(FE_RN_1321_0), .b(FE_RN_1319_0), .o(n_15908) );
na02f80 g764896 ( .a(n_15438), .b(n_15390), .o(n_15561) );
in01f80 g767901 ( .a(n_12768), .o(n_12796) );
in01f80 g762209 ( .a(n_18811), .o(n_18812) );
na02f80 g765632 ( .a(n_14943), .b(n_14963), .o(n_15047) );
in01f80 newInst_2052 ( .a(newNet_2051), .o(newNet_2052) );
in01f80 newInst_111 ( .a(newNet_110), .o(newNet_111) );
na02f80 g743425 ( .a(n_36668), .b(n_36750), .o(n_36702) );
in01f80 newInst_2743 ( .a(newNet_2742), .o(newNet_2743) );
in01f80 newInst_49 ( .a(newNet_39), .o(newNet_49) );
no02f80 FE_RC_2350_0 ( .a(FE_RN_901_0), .b(FE_RN_902_0), .o(FE_RN_903_0) );
no02f80 FE_RC_2481_0 ( .a(n_40130), .b(n_40128), .o(FE_RN_1001_0) );
in01f80 g774068 ( .a(delay_xor_ln21_unr6_stage3_stallmux_q_22_), .o(n_6746) );
na02f80 g762136 ( .a(n_18165), .b(n_16779), .o(n_18246) );
in01f80 g764715 ( .a(FE_OCPN973_n_15900), .o(n_15939) );
na02f80 g753271 ( .a(n_27287), .b(FE_OCP_RBN2892_n_26152), .o(n_27414) );
in01f80 g779095 ( .a(n_2067), .o(n_2087) );
in01f80 FE_OCPC891_n_7802 ( .a(FE_OCPN889_n_7802), .o(FE_OCPN891_n_7802) );
ao22s80 g777205 ( .a(n_3639), .b(n_4642), .c(n_3638), .d(n_3025), .o(n_3677) );
ms00f80 delay_xor_ln21_unr15_stage6_stallmux_q_reg_2_ ( .ck(newNet_960), .d(n_22629), .o(delay_xor_ln21_unr15_stage6_stallmux_q_2_) );
in01f80 g741387 ( .a(FE_OCP_RBN2638_n_38806), .o(n_38870) );
ao12f80 g752492 ( .a(n_27373), .b(n_27620), .c(n_27462), .o(n_27690) );
na02f80 g754562 ( .a(n_26640), .b(n_26606), .o(n_26683) );
oa12f80 g759369 ( .a(n_21296), .b(n_21699), .c(n_21205), .o(n_21757) );
na02f80 g740426 ( .a(FE_OCP_RBN3026_n_39942), .b(n_39559), .o(n_40204) );
na02f80 g747207 ( .a(n_46413), .b(n_32712), .o(n_32672) );
in01f80 g773011 ( .a(n_8143), .o(n_8144) );
na02f80 g737044 ( .a(n_43230), .b(n_43172), .o(n_43485) );
in01f80 g780418 ( .a(n_823), .o(n_824) );
oa22f80 g784547 ( .a(FE_OFN801_n_46285), .b(n_46986), .c(FE_OCP_RBN3044_n_46337), .d(n_11412), .o(n_46368) );
in01f80 g771043 ( .a(delay_sub_ln23_0_unr8_stage4_stallmux_q_6_), .o(n_10035) );
ao12f80 g761037 ( .a(n_19609), .b(n_20115), .c(n_19913), .o(n_19914) );
in01f80 g748151 ( .a(n_31988), .o(n_31989) );
in01f80 g770235 ( .a(n_10669), .o(n_10670) );
in01f80 newInst_2642 ( .a(newNet_2515), .o(newNet_2642) );
in01f80 FE_OCP_RBC2401_n_13954 ( .a(n_13954), .o(FE_OCP_RBN2401_n_13954) );
oa22f80 g781155 ( .a(n_194), .b(n_149), .c(n_199), .d(n_150), .o(n_384) );
no02f80 g749130 ( .a(n_30847), .b(n_27130), .o(n_30963) );
in01f80 g745142 ( .a(n_34894), .o(n_35569) );
na02f80 g756869 ( .a(n_23867), .b(n_23832), .o(n_23868) );
na02f80 g741304 ( .a(FE_OCP_RBN2549_n_44944), .b(n_38872), .o(n_38959) );
in01f80 g779471 ( .a(n_1931), .o(n_1932) );
no02f80 g760182 ( .a(n_20605), .b(n_20567), .o(n_20658) );
in01f80 g737625 ( .a(n_42461), .o(n_42462) );
na02f80 g762303 ( .a(n_18059), .b(n_18061), .o(n_18153) );
ms00f80 delay_xor_ln22_unr9_stage4_stallmux_q_reg_6_ ( .ck(newNet_147), .d(n_46376), .o(delay_xor_ln22_unr9_stage4_stallmux_q_6_) );
in01f80 newInst_984 ( .a(newNet_181), .o(newNet_984) );
in01f80 newInst_841 ( .a(newNet_840), .o(newNet_841) );
na03f80 g763484 ( .a(n_17536), .b(n_17537), .c(n_17610), .o(n_17734) );
in01f80 g748578 ( .a(n_31426), .o(n_31385) );
in01f80 newInst_686 ( .a(newNet_685), .o(newNet_686) );
na02f80 g780408 ( .a(n_787), .b(n_1002), .o(n_817) );
na02f80 g777736 ( .a(n_3440), .b(n_3457), .o(n_3460) );
na02f80 g774464 ( .a(n_6789), .b(delay_sub_ln23_0_unr5_stage3_stallmux_q_23_), .o(n_6844) );
in01f80 g736871 ( .a(n_43607), .o(n_43608) );
in01f80 FE_OCP_RBC2443_n_42051 ( .a(n_42051), .o(FE_OCP_RBN2443_n_42051) );
na02f80 g757096 ( .a(n_23235), .b(n_23196), .o(n_23270) );
in01f80 newInst_1208 ( .a(newNet_1207), .o(newNet_1208) );
ao22s80 FE_RC_3959_0 ( .a(n_33287), .b(FE_OCP_RBN2254_n_33729), .c(n_33729), .d(n_33288), .o(n_33825) );
in01f80 fopt782909 ( .a(n_11726), .o(n_44356) );
na02f80 g759011 ( .a(n_21603), .b(n_21530), .o(n_21632) );
na02f80 g761787 ( .a(n_18894), .b(FE_OCPN1454_n_18559), .o(n_18561) );
no02f80 g752030 ( .a(n_28067), .b(n_28120), .o(n_28073) );
no02f80 g775550 ( .a(n_5632), .b(FE_OCP_RBN2746_n_47011), .o(n_5681) );
oa12f80 g742624 ( .a(n_37502), .b(n_37501), .c(n_37500), .o(n_37974) );
na02f80 g737920 ( .a(n_42202), .b(n_41960), .o(n_42327) );
oa22f80 FE_RC_3880_0 ( .a(n_22393), .b(n_24932), .c(n_22484), .d(n_24933), .o(n_25036) );
na02f80 g759301 ( .a(n_21118), .b(n_45091), .o(n_21152) );
na02f80 g766496 ( .a(n_14118), .b(FE_OCP_RBN2208_n_12907), .o(n_14230) );
oa12f80 g743983 ( .a(n_35683), .b(n_35689), .c(n_44180), .o(n_35916) );
no03m80 g743818 ( .a(n_37190), .b(n_37166), .c(n_37136), .o(n_37201) );
in01f80 fopt782792 ( .a(n_35487), .o(n_44211) );
no02f80 g744209 ( .a(n_36130), .b(n_35740), .o(n_36254) );
na02f80 g761030 ( .a(FE_OCP_RBN3830_n_19204), .b(n_19345), .o(n_19347) );
no02f80 g779619 ( .a(FE_OCP_RBN3362_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .b(delay_xor_ln21_unr3_stage2_stallmux_q_4_), .o(n_1390) );
in01f80 g738172 ( .a(n_41996), .o(n_41997) );
in01f80 FE_OCP_RBC2906_n_16230 ( .a(n_16230), .o(FE_OCP_RBN2906_n_16230) );
oa22f80 g739692 ( .a(n_40540), .b(n_40354), .c(n_40541), .d(n_40353), .o(n_40567) );
in01f80 g736799 ( .a(n_43347), .o(n_43348) );
na02f80 g762786 ( .a(n_17887), .b(n_17886), .o(n_17966) );
in01f80 newInst_2424 ( .a(newNet_2423), .o(newNet_2424) );
na02f80 g774884 ( .a(n_6281), .b(n_6204), .o(n_6302) );
in01f80 FE_OCP_DRV_C1580_n_35482 ( .a(FE_OCP_DRV_N1579_n_35482), .o(FE_OCP_DRV_N1580_n_35482) );
in01f80 g748863 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_1_), .o(n_31260) );
na02f80 g736768 ( .a(n_43320), .b(n_43181), .o(n_43182) );
no02f80 g762820 ( .a(n_17700), .b(n_17772), .o(n_17773) );
no02f80 g754941 ( .a(n_25185), .b(n_25184), .o(n_25186) );
na02f80 g763372 ( .a(FE_OCP_RBN3724_n_16975), .b(n_15479), .o(n_17331) );
no02f80 g766337 ( .a(n_14161), .b(n_14135), .o(n_14251) );
in01f80 FE_OCP_RBC3855_n_21224 ( .a(n_21224), .o(FE_OCP_RBN3855_n_21224) );
oa22f80 g747761 ( .a(n_32216), .b(n_32137), .c(n_32217), .d(n_32136), .o(n_32262) );
in01f80 FE_OCPC870_n_2737 ( .a(FE_OCP_RBN2292_n_2438), .o(FE_OCPN870_n_2737) );
in01f80 g743413 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_31_), .o(n_36590) );
in01f80 g761611 ( .a(n_19787), .o(n_19845) );
ao12f80 g777712 ( .a(n_3125), .b(n_3345), .c(n_3329), .o(n_3357) );
na02f80 g759232 ( .a(n_21344), .b(FE_OCP_DRV_N1590_n_21343), .o(n_21381) );
no02f80 g752027 ( .a(n_28071), .b(n_27968), .o(n_28102) );
na02f80 g768303 ( .a(n_12531), .b(n_12387), .o(n_12532) );
na02f80 g776977 ( .a(n_3941), .b(n_4036), .o(n_4037) );
oa22f80 g775111 ( .a(n_5941), .b(n_5599), .c(n_5927), .d(n_5598), .o(n_6063) );
no02f80 g739329 ( .a(n_45144), .b(n_40695), .o(n_40781) );
ao22s80 g757461 ( .a(FE_OCP_RBN3823_n_44061), .b(delay_xor_ln22_unr15_stage6_stallmux_q_5_), .c(n_22865), .d(FE_OCP_RBN3822_n_44061), .o(n_22937) );
oa12f80 g777918 ( .a(n_2358), .b(n_3096), .c(n_2314), .o(n_3133) );
na02f80 g751199 ( .a(n_29818), .b(n_29817), .o(n_29884) );
oa12f80 g761501 ( .a(n_18434), .b(FE_OCP_RBN1836_FE_RN_1542_0), .c(n_18346), .o(n_18873) );
na02f80 g756172 ( .a(n_25251), .b(n_25250), .o(n_24793) );
ao12f80 g745178 ( .a(n_34631), .b(n_34656), .c(n_34630), .o(n_34706) );
na02f80 FE_RC_2722_0 ( .a(n_8355), .b(FE_RN_1149_0), .o(FE_RN_1150_0) );
in01f80 g760761 ( .a(FE_OCP_RBN2419_n_19601), .o(n_19654) );
na02f80 g751463 ( .a(n_28720), .b(n_28719), .o(n_28737) );
na02f80 g742136 ( .a(n_38120), .b(n_38291), .o(n_38327) );
oa12f80 g741489 ( .a(n_38711), .b(n_38710), .c(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38746) );
in01f80 g764814 ( .a(n_15761), .o(n_15847) );
in01f80 g745595 ( .a(n_34339), .o(n_34846) );
no02f80 g743933 ( .a(n_36146), .b(n_44223), .o(n_36245) );
oa12f80 g742015 ( .a(n_38009), .b(FE_OCP_RBN3445_n_37945), .c(n_37566), .o(n_38461) );
na02f80 g773770 ( .a(n_7205), .b(n_7233), .o(n_7578) );
na02f80 g767293 ( .a(n_13538), .b(n_13625), .o(n_13551) );
ao12f80 g784433 ( .a(n_46224), .b(n_46197), .c(delay_sub_ln23_0_unr28_stage9_stallmux_q_10_), .o(n_46245) );
na02f80 g739586 ( .a(n_40602), .b(n_44610), .o(n_40612) );
in01f80 g736506 ( .a(n_43675), .o(n_43676) );
na02f80 FE_RC_2634_0 ( .a(FE_RN_1096_0), .b(FE_RN_1097_0), .o(FE_RN_68_0) );
na02f80 g769062 ( .a(FE_OCP_RBN2009_n_45622), .b(n_45224), .o(n_11774) );
in01f80 g759383 ( .a(n_20862), .o(n_20859) );
na02f80 g774241 ( .a(n_6526), .b(n_6619), .o(n_6637) );
na02f80 g738744 ( .a(n_41537), .b(n_41372), .o(n_41684) );
in01f80 g764009 ( .a(n_18140), .o(n_18230) );
in01f80 g757411 ( .a(n_23014), .o(n_23222) );
in01f80 FE_OCP_RBC1198_n_30619 ( .a(n_30619), .o(FE_OCP_RBN1198_n_30619) );
ms00f80 delay_sub_ln21_0_unr2_stage2_stallmux_q_reg_9_ ( .ck(newNet_2132), .d(n_934), .o(delay_sub_ln21_0_unr2_stage2_stallmux_q_9_) );
in01f80 g755553 ( .a(n_24745), .o(n_24774) );
in01f80 FE_OCP_RBC2157_n_1614 ( .a(n_1614), .o(FE_OCP_RBN2157_n_1614) );
in01f80 FE_OCP_RBC2844_n_10326 ( .a(FE_OCP_RBN2843_n_10326), .o(FE_OCP_RBN2844_n_10326) );
oa22f80 g748565 ( .a(n_31545), .b(n_31487), .c(n_31544), .d(n_31486), .o(n_31673) );
in01f80 g752669 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .o(n_27475) );
no02f80 g771984 ( .a(FE_OCP_RBN3546_n_44575), .b(n_8781), .o(n_8959) );
no02f80 g770687 ( .a(n_9941), .b(FE_OCP_RBN2474_n_8664), .o(n_10020) );
oa22f80 FE_RC_357_0 ( .a(n_17349), .b(n_17333), .c(n_17350), .d(n_17392), .o(n_17594) );
oa12f80 g771554 ( .a(n_9393), .b(n_9392), .c(FE_OFN361_n_9391), .o(n_9474) );
no02f80 g779154 ( .a(FE_OCP_RBN2182_n_1916), .b(n_1685), .o(n_1967) );
no02f80 g753814 ( .a(n_26433), .b(FE_RN_1667_0), .o(n_26436) );
in01f80 g737999 ( .a(n_42201), .o(n_42270) );
na02f80 g774959 ( .a(n_6220), .b(n_6148), .o(n_6225) );
in01f80 g743603 ( .a(n_36444), .o(n_36472) );
in01f80 g740881 ( .a(n_39218), .o(n_39219) );
na02f80 g771065 ( .a(n_9629), .b(FE_OCPN903_n_44581), .o(n_9644) );
in01f80 newInst_1389 ( .a(newNet_1388), .o(newNet_1389) );
oa22f80 FE_RC_988_0 ( .a(n_24350), .b(n_27800), .c(n_27796), .d(n_27767), .o(n_27858) );
na02f80 g777283 ( .a(FE_OCPN959_n_3951), .b(FE_OFN819_n_4298), .o(n_4361) );
no02f80 g744582 ( .a(n_35296), .b(n_35152), .o(n_35332) );
na02f80 g765346 ( .a(n_15258), .b(FE_OCP_RBN2760_n_15180), .o(n_15259) );
no02f80 g765660 ( .a(n_14962), .b(FE_OCP_RBN3485_n_13667), .o(n_14987) );
in01f80 g766562 ( .a(n_13955), .o(n_13956) );
in01f80 g778283 ( .a(n_2911), .o(n_2912) );
in01f80 g756326 ( .a(n_23949), .o(n_24005) );
no02f80 g764283 ( .a(n_16321), .b(n_16273), .o(n_16379) );
in01f80 g736647 ( .a(n_43441), .o(n_43479) );
oa12f80 g736273 ( .a(n_310), .b(n_43862), .c(FE_OFN4_n_43918), .o(n_43898) );
na02f80 g752550 ( .a(n_27602), .b(n_27397), .o(n_27621) );
na02f80 g749539 ( .a(n_31709), .b(n_31212), .o(n_31782) );
in01f80 g772753 ( .a(n_8106), .o(n_8138) );
na02f80 g766313 ( .a(n_14286), .b(n_14240), .o(n_14241) );
ms00f80 delay_sub_ln23_0_unr12_stage5_stallmux_q_reg_26_ ( .ck(newNet_1830), .d(n_17017), .o(delay_sub_ln23_0_unr12_stage5_stallmux_q_26_) );
no02f80 g760845 ( .a(n_19439), .b(FE_OFN780_n_17093), .o(n_19530) );
no02f80 g760960 ( .a(n_19214), .b(FE_OFN779_n_17093), .o(n_19254) );
no02f80 g740181 ( .a(n_39812), .b(n_39945), .o(n_39977) );
in01f80 FE_RC_4189_0 ( .a(n_24158), .o(FE_RN_1835_0) );
in01f80 g777586 ( .a(n_3562), .o(n_3638) );
oa12f80 g777687 ( .a(n_3355), .b(n_3354), .c(n_3353), .o(n_5197) );
in01f80 g777545 ( .a(n_4556), .o(n_4606) );
na02f80 g742520 ( .a(n_37581), .b(delay_sub_ln23_0_unr24_stage9_stallmux_q), .o(n_37601) );
in01f80 fopt783797 ( .a(n_45479), .o(n_45474) );
in01f80 g761081 ( .a(n_19213), .o(n_19207) );
in01f80 g776610 ( .a(FE_OCP_RBN2669_n_4158), .o(n_5009) );
no02f80 g753963 ( .a(n_26188), .b(n_23466), .o(n_26217) );
ao12f80 g749579 ( .a(n_30017), .b(n_30285), .c(n_30021), .o(n_30494) );
in01f80 FE_OCP_RBC2262_n_33691 ( .a(n_33691), .o(FE_OCP_RBN2262_n_33691) );
na02f80 g751772 ( .a(n_29203), .b(n_29149), .o(n_29204) );
no02f80 g753558 ( .a(n_27406), .b(n_26860), .o(n_27449) );
in01f80 g778626 ( .a(n_2617), .o(n_2618) );
no02f80 g780444 ( .a(n_764), .b(n_7), .o(n_796) );
no02f80 FE_RC_1137_0 ( .a(FE_RN_344_0), .b(n_2821), .o(n_2840) );
in01f80 newInst_3741 ( .a(newNet_3740), .o(newNet_3741) );
no02f80 g778110 ( .a(n_2761), .b(n_2891), .o(n_2892) );
na02f80 g746375 ( .a(n_33471), .b(n_33470), .o(n_33472) );
no02f80 FE_RC_3108_0 ( .a(n_26846), .b(FE_RN_1374_0), .o(FE_RN_1375_0) );
na02f80 g765002 ( .a(FE_OCP_RBN3661_n_15429), .b(n_14452), .o(n_15467) );
in01f80 g763030 ( .a(n_17717), .o(n_17645) );
na02f80 FE_RC_4098_0 ( .a(FE_OCP_RBN1198_n_30619), .b(n_30729), .o(FE_RN_1792_0) );
in01f80 g775645 ( .a(n_5308), .o(n_5309) );
oa12f80 g755936 ( .a(n_24250), .b(n_24270), .c(n_24249), .o(n_24342) );
ao12f80 g742936 ( .a(n_37000), .b(n_46256), .c(delay_add_ln22_unr23_stage9_stallmux_q_21_), .o(n_37431) );
in01f80 fopt783582 ( .a(n_45213), .o(n_45212) );
in01f80 g754706 ( .a(n_26308), .o(n_26346) );
in01f80 FE_OCPC985_n_25210 ( .a(FE_OCPN984_n_25210), .o(FE_OCPN985_n_25210) );
in01f80 newInst_2822 ( .a(newNet_2821), .o(newNet_2822) );
na02f80 g753645 ( .a(n_26627), .b(n_26626), .o(n_26723) );
na02f80 g758037 ( .a(n_22812), .b(n_22699), .o(n_22700) );
in01f80 g747999 ( .a(n_31908), .o(n_31938) );
no02f80 g736971 ( .a(FE_OCPN913_n_43022), .b(n_43208), .o(n_43359) );
no02f80 g778424 ( .a(n_2616), .b(delay_sub_ln21_0_unr2_stage2_stallmux_q_26_), .o(n_2731) );
no02f80 g755272 ( .a(n_26310), .b(n_25683), .o(n_25684) );
oa12f80 g738272 ( .a(n_41734), .b(n_41824), .c(n_41619), .o(n_41940) );
na02f80 g766103 ( .a(n_14553), .b(FE_OCP_RBN2450_n_14114), .o(n_14609) );
no02f80 g769073 ( .a(n_11537), .b(n_11640), .o(n_11775) );
ao12f80 g773113 ( .a(n_7816), .b(n_8309), .c(n_7105), .o(n_8479) );
in01f80 g773135 ( .a(n_7857), .o(n_7914) );
in01f80 g752363 ( .a(n_27785), .o(n_27758) );
in01f80 g752959 ( .a(n_28176), .o(n_28075) );
in01f80 FE_OCP_RBC2736_n_14985 ( .a(n_14985), .o(FE_OCP_RBN2736_n_14985) );
in01f80 newInst_2676 ( .a(newNet_2675), .o(newNet_2676) );
in01f80 newInst_155 ( .a(newNet_154), .o(newNet_155) );
in01f80 g744467 ( .a(n_35490), .o(n_35491) );
in01f80 newInst_1050 ( .a(newNet_1049), .o(newNet_1050) );
no02f80 g742027 ( .a(n_38082), .b(n_44033), .o(n_38083) );
ms00f80 cos_out_reg_9_ ( .ck(newNet_3663), .d(n_43767), .o(cos_out_9) );
na02f80 g736785 ( .a(n_43341), .b(n_43393), .o(n_43427) );
in01f80 g769981 ( .a(n_11069), .o(n_11070) );
oa22f80 g758369 ( .a(n_21904), .b(n_21956), .c(n_21903), .d(n_21955), .o(n_21973) );
in01f80 g740843 ( .a(n_39349), .o(n_39350) );
no02f80 FE_RC_1844_0 ( .a(n_35872), .b(FE_RN_559_0), .o(FE_RN_560_0) );
in01f80 FE_OCP_RBC3534_n_13765 ( .a(FE_OCP_RBN3530_n_13765), .o(FE_OCP_RBN3534_n_13765) );
no02f80 g776194 ( .a(n_4887), .b(n_4886), .o(n_4956) );
in01f80 newInst_3217 ( .a(newNet_1619), .o(newNet_3217) );
ms00f80 delay_add_ln22_unr14_stage6_stallmux_q_reg_10_ ( .ck(newNet_3568), .d(n_21915), .o(delay_add_ln22_unr14_stage6_stallmux_q_10_) );
na02f80 g740821 ( .a(n_39265), .b(n_39292), .o(n_39878) );
in01f80 g759096 ( .a(n_21130), .o(n_21131) );
no02f80 g755267 ( .a(n_24944), .b(n_24943), .o(n_24972) );
in01f80 g756368 ( .a(n_25085), .o(n_24382) );
in01f80 newInst_3064 ( .a(newNet_3063), .o(newNet_3064) );
in01f80 g738368 ( .a(n_41771), .o(n_41772) );
in01f80 FE_OCP_RBC3088_FE_OCPN1052_n_31674 ( .a(FE_OCPN1052_n_31674), .o(FE_OCP_RBN3088_FE_OCPN1052_n_31674) );
in01f80 g753897 ( .a(n_26376), .o(n_26324) );
na02f80 g771524 ( .a(n_9595), .b(n_9558), .o(n_9559) );
no02f80 g751170 ( .a(n_29932), .b(n_29710), .o(n_30094) );
ms00f80 sin_out_reg_31_ ( .ck(newNet_27), .d(n_43916), .o(sin_out_31) );
na02f80 g777767 ( .a(n_3375), .b(n_3226), .o(n_3376) );
no02f80 g740829 ( .a(n_39436), .b(n_38998), .o(n_39437) );
in01f80 g756199 ( .a(n_24084), .o(n_24085) );
no02f80 g778738 ( .a(FE_OCPN1234_n_2414), .b(n_2562), .o(n_2609) );
no02f80 g744242 ( .a(n_46216), .b(n_36854), .o(n_37839) );
in01f80 g747528 ( .a(n_32518), .o(n_32470) );
in01f80 FE_RC_1978_0 ( .a(n_19722), .o(FE_RN_642_0) );
in01f80 g778585 ( .a(n_2712), .o(n_2706) );
no02f80 g747226 ( .a(n_33795), .b(n_33794), .o(n_33796) );
in01f80 g775720 ( .a(n_5212), .o(n_5213) );
na02f80 g775440 ( .a(n_5568), .b(n_5581), .o(n_5654) );
in01f80 g743237 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_3_), .o(n_36872) );
no02f80 g738619 ( .a(n_41376), .b(n_41374), .o(n_41405) );
ms00f80 delay_sub_ln21_0_unr5_stage3_stallmux_q_reg_30_ ( .ck(newNet_2068), .d(n_6739), .o(delay_sub_ln21_0_unr5_stage3_stallmux_q_30_) );
no02f80 FE_RC_3978_0 ( .a(FE_OFN788_n_25834), .b(FE_RN_1723_0), .o(FE_RN_1724_0) );
in01f80 g757867 ( .a(n_22421), .o(n_22422) );
no02f80 g766557 ( .a(FE_OCP_RBN2413_n_13960), .b(FE_OCP_RBN3507_n_13860), .o(n_14055) );
in01f80 FE_RC_3408_0 ( .a(FE_RN_740_0), .o(FE_RN_1475_0) );
in01f80 g736663 ( .a(n_43374), .o(n_43333) );
na02f80 g760930 ( .a(n_19284), .b(n_18463), .o(n_19333) );
in01f80 FE_OCP_RBC3598_FE_OCPN1243_n_44460 ( .a(FE_OCP_RBN3597_FE_OCPN1243_n_44460), .o(FE_OCP_RBN3598_FE_OCPN1243_n_44460) );
ms00f80 delay_add_ln22_unr8_stage4_stallmux_q_reg_7_ ( .ck(newNet_2802), .d(n_10496), .o(delay_add_ln22_unr8_stage4_stallmux_q_7_) );
in01f80 g768909 ( .a(n_11941), .o(n_11942) );
no02f80 g739238 ( .a(n_40972), .b(n_40988), .o(n_41032) );
no02f80 g781323 ( .a(n_7), .b(beta_19), .o(n_135) );
in01f80 FE_RC_3098_0 ( .a(n_16333), .o(FE_RN_1369_0) );
in01f80 g755522 ( .a(n_25261), .o(n_25262) );
oa12f80 g768778 ( .a(n_11715), .b(n_11874), .c(n_11514), .o(n_11985) );
no02f80 g747668 ( .a(n_33990), .b(n_33700), .o(n_33760) );
oa12f80 g767370 ( .a(n_13586), .b(n_13585), .c(n_13584), .o(n_14107) );
no02f80 g772644 ( .a(n_8205), .b(n_8184), .o(n_8296) );
oa22f80 g737302 ( .a(n_42889), .b(n_42788), .c(n_42855), .d(n_42789), .o(n_43208) );
in01f80 newInst_942 ( .a(newNet_209), .o(newNet_942) );
no02f80 g756234 ( .a(n_24670), .b(n_24355), .o(n_24742) );
in01f80 FE_OFC4_n_43918 ( .a(FE_OFN0_n_43918), .o(FE_OFN4_n_43918) );
na02f80 g761353 ( .a(n_19128), .b(n_19127), .o(n_19129) );
na02f80 g764496 ( .a(n_16041), .b(n_14524), .o(n_16090) );
na02f80 g778612 ( .a(FE_OCPN871_n_2737), .b(n_2719), .o(n_2817) );
na02f80 g770464 ( .a(n_10557), .b(n_10603), .o(n_10725) );
in01f80 g755764 ( .a(n_24486), .o(n_24633) );
in01f80 g760073 ( .a(n_21626), .o(n_21719) );
no02f80 g764790 ( .a(n_45134), .b(n_15271), .o(n_15596) );
in01f80 g737229 ( .a(n_43251), .o(n_42969) );
no02f80 g757091 ( .a(n_23263), .b(n_23322), .o(n_23345) );
in01f80 g759029 ( .a(n_21236), .o(n_21281) );
oa22f80 FE_RC_435_0 ( .a(n_17330), .b(n_17599), .c(n_17494), .d(n_17327), .o(n_17728) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_19_ ( .ck(newNet_1412), .d(n_36666), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_19_) );
no02f80 FE_RC_3396_0 ( .a(FE_RN_1469_0), .b(FE_RN_1470_0), .o(FE_RN_1471_0) );
in01f80 g770434 ( .a(n_10582), .o(n_10564) );
na02f80 g766510 ( .a(n_14092), .b(n_12877), .o(n_14117) );
in01f80 FE_OCP_RBC2154_n_32772 ( .a(n_32772), .o(FE_OCP_RBN2154_n_32772) );
oa22f80 g746427 ( .a(n_33308), .b(n_33262), .c(n_33307), .d(n_33263), .o(n_34294) );
in01f80 newInst_2451 ( .a(newNet_2450), .o(newNet_2451) );
oa22f80 g779139 ( .a(n_1916), .b(n_1720), .c(FE_OCP_RBN2181_n_1916), .d(n_1719), .o(n_2004) );
in01f80 g769338 ( .a(n_11607), .o(n_11547) );
in01f80 FE_OCP_RBC1852_n_22556 ( .a(n_22556), .o(FE_OCP_RBN1852_n_22556) );
in01f80 FE_OCP_RBC3723_n_16975 ( .a(n_16975), .o(FE_OCP_RBN3723_n_16975) );
na02f80 FE_RC_911_0 ( .a(FE_RN_267_0), .b(FE_RN_268_0), .o(FE_RN_269_0) );
in01f80 FE_OCP_RBC2931_n_5307 ( .a(n_5307), .o(FE_OCP_RBN2931_n_5307) );
na02f80 g744699 ( .a(n_35269), .b(n_35268), .o(n_35270) );
no02f80 g748257 ( .a(FE_OCP_RBN3734_n_31819), .b(n_30541), .o(n_32054) );
in01f80 g771469 ( .a(n_9116), .o(n_9166) );
in01f80 newInst_3024 ( .a(newNet_380), .o(newNet_3024) );
na02f80 g778296 ( .a(n_2559), .b(n_2464), .o(n_2688) );
no02f80 g746206 ( .a(n_33664), .b(n_34037), .o(n_33782) );
in01f80 g781291 ( .a(n_52), .o(n_158) );
no02f80 g755455 ( .a(n_24603), .b(FE_OFN784_delay_sub_ln23_0_unr15_stage6_stallmux_q), .o(n_24788) );
no02f80 g741689 ( .a(n_38529), .b(delay_sub_ln23_0_unr25_stage9_stallmux_q), .o(n_38566) );
na02f80 g756726 ( .a(n_23431), .b(n_23315), .o(n_23445) );
na02f80 g741324 ( .a(FE_OCP_RBN2546_n_44944), .b(FE_OCP_RBN2485_n_38601), .o(n_39175) );
na02f80 g751992 ( .a(n_28781), .b(n_28834), .o(n_28858) );
no02f80 g768279 ( .a(n_12573), .b(n_12567), .o(n_12568) );
na02f80 g736436 ( .a(FE_OCP_RBN3131_n_43762), .b(n_43642), .o(n_43792) );
ao12f80 g751318 ( .a(n_29243), .b(n_29601), .c(n_29285), .o(n_29638) );
in01f80 newInst_3674 ( .a(newNet_2830), .o(newNet_3674) );
no02f80 g756166 ( .a(n_24791), .b(n_24354), .o(n_24818) );
na02f80 FE_RC_2599_0 ( .a(FE_RN_1077_0), .b(n_3456), .o(FE_RN_1078_0) );
in01f80 FE_OCP_RBC2918_n_16084 ( .a(n_16084), .o(FE_OCP_RBN2918_n_16084) );
in01f80 g771071 ( .a(n_9800), .o(n_9801) );
no02f80 g750698 ( .a(n_29232), .b(n_28739), .o(n_29323) );
no02f80 FE_RC_2814_0 ( .a(n_34365), .b(n_45185), .o(FE_RN_1205_0) );
ao12f80 g738613 ( .a(n_41828), .b(n_41716), .c(n_41484), .o(n_42008) );
in01f80 g764644 ( .a(n_15816), .o(n_15912) );
in01f80 g753361 ( .a(n_26993), .o(n_26922) );
oa12f80 g739014 ( .a(n_41053), .b(n_41119), .c(n_41038), .o(n_41147) );
in01f80 FE_OCP_RBC1136_n_17040 ( .a(n_17040), .o(FE_OCP_RBN1136_n_17040) );
no02f80 FE_RC_983_0 ( .a(n_27254), .b(n_27639), .o(FE_RN_283_0) );
na02f80 g763698 ( .a(n_17367), .b(n_17265), .o(n_17368) );
no02f80 FE_RC_3195_0 ( .a(FE_RN_1418_0), .b(FE_RN_1419_0), .o(FE_RN_1420_0) );
na02f80 g763201 ( .a(n_17249), .b(n_17233), .o(n_17402) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_26_ ( .ck(newNet_3131), .d(n_40559), .o(delay_add_ln22_unr27_stage10_stallmux_q_26_) );
na02f80 g759418 ( .a(n_20886), .b(n_20885), .o(n_20917) );
in01f80 g767948 ( .a(n_12788), .o(n_12843) );
in01f80 g753425 ( .a(n_26883), .o(n_26828) );
no02f80 g753676 ( .a(n_26588), .b(FE_OCPN1526_n_26587), .o(n_26659) );
in01f80 g766222 ( .a(n_14511), .o(n_14467) );
in01f80 g747504 ( .a(delay_xor_ln22_unr21_stage8_stallmux_q_0_), .o(n_32543) );
na02f80 g748654 ( .a(n_31209), .b(n_31030), .o(n_31273) );
no02f80 g762834 ( .a(n_18104), .b(n_17469), .o(n_18158) );
na02f80 g766161 ( .a(n_14444), .b(n_13514), .o(n_14477) );
in01f80 FE_OCP_RBC2161_n_40687 ( .a(n_40687), .o(FE_OCP_RBN2161_n_40687) );
in01f80 g779757 ( .a(n_1663), .o(n_1739) );
in01f80 FE_OCP_DRV_C1565_n_28654 ( .a(n_28654), .o(FE_OCP_DRV_N1565_n_28654) );
in01f80 g773450 ( .a(n_7881), .o(n_7851) );
oa12f80 g755079 ( .a(n_25075), .b(n_25074), .c(n_25073), .o(n_26752) );
ms00f80 delay_xor_ln22_unr15_stage6_stallmux_q_reg_9_ ( .ck(newNet_477), .d(n_22802), .o(delay_xor_ln22_unr15_stage6_stallmux_q_9_) );
ao12f80 g779515 ( .a(n_1685), .b(FE_OCP_RBN3243_delay_sub_ln23_0_unr2_stage2_stallmux_q_29_), .c(delay_xor_ln22_unr3_stage2_stallmux_q_13_), .o(n_1719) );
oa12f80 g779216 ( .a(n_1724), .b(n_1838), .c(n_1678), .o(n_1874) );
na02f80 g750506 ( .a(n_29450), .b(FE_OFN788_n_25834), .o(n_29484) );
no02f80 g738677 ( .a(n_41525), .b(n_41656), .o(n_41725) );
no02f80 g763444 ( .a(FE_OCP_RBN3724_n_16975), .b(n_16192), .o(n_17120) );
oa12f80 g742156 ( .a(n_37810), .b(n_37863), .c(n_37832), .o(n_37917) );
na02f80 g767688 ( .a(n_13101), .b(n_12969), .o(n_13132) );
oa22f80 g769883 ( .a(n_11069), .b(n_10206), .c(n_11070), .d(n_10207), .o(n_11153) );
oa12f80 g742694 ( .a(n_37356), .b(n_37355), .c(n_37354), .o(n_37889) );
no02f80 g754540 ( .a(n_26385), .b(n_26345), .o(n_26452) );
no02f80 g776446 ( .a(n_4588), .b(n_4587), .o(n_4735) );
in01f80 newInst_341 ( .a(newNet_61), .o(newNet_341) );
na02f80 g747107 ( .a(n_32969), .b(n_33007), .o(n_33110) );
oa22f80 g756355 ( .a(n_23948), .b(n_23652), .c(n_23889), .d(n_23651), .o(n_25126) );
na02f80 g767524 ( .a(n_13222), .b(n_13221), .o(n_13223) );
in01f80 FE_OCP_RBC3567_n_29857 ( .a(FE_OCP_RBN3565_n_29857), .o(FE_OCP_RBN3567_n_29857) );
na02f80 g745956 ( .a(n_33944), .b(n_33965), .o(n_34052) );
in01f80 g762870 ( .a(n_17720), .o(n_17721) );
na02f80 FE_RC_3153_0 ( .a(n_21353), .b(n_21159), .o(FE_RN_1399_0) );
ms00f80 delay_xor_ln22_unr12_stage5_stallmux_q_reg_15_ ( .ck(newNet_582), .d(n_17776), .o(delay_xor_ln22_unr12_stage5_stallmux_q_15_) );
in01f80 g755541 ( .a(n_24578), .o(n_24579) );
in01f80 g768891 ( .a(n_11945), .o(n_11946) );
na02f80 g776653 ( .a(n_4340), .b(n_4339), .o(n_4501) );
in01f80 g773174 ( .a(n_7919), .o(n_7920) );
in01f80 g745802 ( .a(n_34479), .o(n_34480) );
in01f80 g741038 ( .a(n_39331), .o(n_39332) );
ms00f80 delay_sub_ln23_0_unr16_stage6_stallmux_q_reg_16_ ( .ck(newNet_1759), .d(n_22244), .o(delay_sub_ln23_0_unr16_stage6_stallmux_q_16_) );
ao22s80 g736547 ( .a(n_43572), .b(n_43615), .c(n_43571), .d(n_43616), .o(n_43663) );
na02f80 g748222 ( .a(n_31718), .b(n_31740), .o(n_31741) );
in01f80 g754306 ( .a(n_26016), .o(n_25956) );
in01f80 FE_RC_2198_0 ( .a(n_26196), .o(FE_RN_789_0) );
no02f80 FE_RC_1839_0 ( .a(FE_OCPN1017_n_23307), .b(FE_OCPN1022_n_23195), .o(FE_RN_556_0) );
in01f80 g749296 ( .a(n_30841), .o(n_30867) );
na02f80 g761313 ( .a(n_18978), .b(n_18973), .o(n_19004) );
no02f80 g746061 ( .a(n_33809), .b(n_33784), .o(n_33908) );
in01f80 g743369 ( .a(n_37828), .o(n_37829) );
oa22f80 FE_RC_735_0 ( .a(FE_OCP_RBN3465_n_7886), .b(n_8402), .c(FE_OCP_RBN3463_n_7886), .d(FE_OCP_RBN2437_n_8402), .o(n_8525) );
no02f80 g766546 ( .a(FE_OCP_RBN2429_n_14018), .b(FE_OCP_RBN2250_n_13017), .o(n_14090) );
in01f80 g743900 ( .a(n_37020), .o(n_37021) );
in01f80 g766844 ( .a(n_13703), .o(n_13745) );
in01f80 g772947 ( .a(n_7929), .o(n_7930) );
in01f80 g762726 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_28_), .o(n_17805) );
in01f80 g768085 ( .a(n_13196), .o(n_13312) );
ao12f80 g750383 ( .a(n_30090), .b(n_30634), .c(n_29976), .o(n_30690) );
in01f80 newInst_452 ( .a(newNet_451), .o(newNet_452) );
no02f80 FE_RC_3650_0 ( .a(n_21923), .b(FE_RN_1601_0), .o(FE_RN_1602_0) );
no02f80 g759295 ( .a(n_21064), .b(n_45024), .o(n_21220) );
na02f80 g770862 ( .a(n_9866), .b(n_9932), .o(n_10100) );
oa12f80 g743853 ( .a(n_37027), .b(n_46250), .c(n_46236), .o(n_37190) );
in01f80 newInst_2089 ( .a(newNet_1462), .o(newNet_2089) );
in01f80 g756557 ( .a(n_23876), .o(n_23945) );
in01f80 g781349 ( .a(beta_0), .o(n_50) );
in01f80 g774605 ( .a(n_46993), .o(n_6479) );
na02f80 g739911 ( .a(n_40231), .b(n_39914), .o(n_40298) );
na02f80 g773426 ( .a(n_7558), .b(delay_add_ln22_unr5_stage3_stallmux_q_28_), .o(n_7554) );
na02f80 g773839 ( .a(n_7089), .b(n_6993), .o(n_7144) );
in01f80 g744481 ( .a(delay_sub_ln21_0_unr23_stage9_stallmux_q_2_), .o(n_35466) );
no02f80 g764652 ( .a(n_15773), .b(n_15336), .o(n_15858) );
in01f80 g754259 ( .a(n_26795), .o(n_26947) );
in01f80 newInst_3143 ( .a(newNet_3142), .o(newNet_3143) );
no02f80 g742203 ( .a(n_37853), .b(n_37808), .o(n_37891) );
in01f80 g736863 ( .a(n_43541), .o(n_43542) );
oa22f80 g759701 ( .a(n_21750), .b(n_21714), .c(n_21721), .d(n_21691), .o(n_21865) );
in01f80 newInst_732 ( .a(newNet_314), .o(newNet_732) );
na02f80 g784396 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_), .o(n_46208) );
in01f80 newInst_2233 ( .a(newNet_1863), .o(newNet_2233) );
in01f80 FE_OCP_RBC2821_n_10023 ( .a(n_10023), .o(FE_OCP_RBN2821_n_10023) );
in01f80 g763427 ( .a(n_16920), .o(n_17488) );
in01f80 newInst_853 ( .a(newNet_676), .o(newNet_853) );
na02f80 g779252 ( .a(n_1795), .b(n_1667), .o(n_1796) );
in01f80 g748329 ( .a(n_31836), .o(n_31837) );
in01f80 g761710 ( .a(n_18716), .o(n_18793) );
ao12f80 g745196 ( .a(n_34598), .b(n_34597), .c(n_34596), .o(n_34707) );
na02f80 g760779 ( .a(n_19615), .b(n_19616), .o(n_19687) );
in01f80 newInst_3319 ( .a(newNet_3318), .o(newNet_3319) );
in01f80 newInst_1438 ( .a(newNet_998), .o(newNet_1438) );
na02f80 g758138 ( .a(FE_OCPN3184_n_22294), .b(n_22417), .o(n_22419) );
na02f80 g763147 ( .a(n_17348), .b(n_17347), .o(n_17482) );
na02f80 g739907 ( .a(n_40092), .b(n_39925), .o(n_40200) );
na02f80 g770696 ( .a(n_10309), .b(FE_OCP_RBN3538_n_8597), .o(n_10423) );
na02f80 g748412 ( .a(n_31730), .b(FE_OCP_RBN2829_n_30731), .o(n_31729) );
ms00f80 delay_sub_ln23_0_unr28_stage9_stallmux_q_reg_5_ ( .ck(newNet_1366), .d(n_36330), .o(delay_sub_ln23_0_unr28_stage9_stallmux_q_5_) );
ao22s80 g736638 ( .a(n_43117), .b(n_43089), .c(n_43116), .d(n_43090), .o(n_43236) );
oa12f80 g738070 ( .a(n_42097), .b(n_42096), .c(n_42095), .o(n_42130) );
no02f80 g772321 ( .a(n_8707), .b(n_8706), .o(n_8708) );
na02f80 g770940 ( .a(n_9895), .b(FE_OCP_RBN3596_FE_OCPN1243_n_44460), .o(n_9968) );
in01f80 newInst_2840 ( .a(newNet_2839), .o(newNet_2840) );
in01f80 fopt783484 ( .a(FE_RN_1585_0), .o(n_45091) );
ao12f80 g767382 ( .a(n_12558), .b(n_13139), .c(n_12576), .o(n_13270) );
in01f80 newInst_11 ( .a(newNet_10), .o(newNet_11) );
no02f80 g756409 ( .a(n_23998), .b(n_24040), .o(n_24041) );
in01f80 g752980 ( .a(n_27088), .o(n_27089) );
na02f80 FE_RC_1731_0 ( .a(n_17865), .b(n_17843), .o(FE_RN_481_0) );
in01f80 g774111 ( .a(n_6723), .o(n_6724) );
in01f80 FE_OCP_RBC2957_n_26231 ( .a(FE_OCP_RBN2955_n_26231), .o(FE_OCP_RBN2957_n_26231) );
ao22s80 g768625 ( .a(n_12185), .b(n_11877), .c(n_47211), .d(n_11878), .o(n_12316) );
ms00f80 delay_sub_ln21_0_unr27_stage10_stallmux_q_reg_17_ ( .ck(newNet_2301), .d(n_40465), .o(delay_sub_ln21_0_unr27_stage10_stallmux_q_17_) );
no02f80 g746576 ( .a(n_33254), .b(n_33236), .o(n_33237) );
na02f80 g743692 ( .a(n_36375), .b(n_35955), .o(n_36424) );
na03f80 g780473 ( .a(n_951), .b(n_977), .c(n_865), .o(n_943) );
no02f80 g749920 ( .a(n_30577), .b(n_30244), .o(n_30263) );
in01f80 g748071 ( .a(n_33314), .o(n_32902) );
na02f80 g770509 ( .a(n_10529), .b(FE_OCP_RBN2539_n_8781), .o(n_10603) );
oa12f80 g745886 ( .a(n_34089), .b(n_34088), .c(n_34087), .o(n_35292) );
oa22f80 FE_RC_236_0 ( .a(n_13016), .b(n_13633), .c(n_13044), .d(n_13594), .o(n_13667) );
na02f80 g769794 ( .a(n_11191), .b(n_11190), .o(n_11293) );
in01f80 g772483 ( .a(n_8513), .o(n_8537) );
in01f80 newInst_3680 ( .a(newNet_3679), .o(newNet_3680) );
in01f80 g777006 ( .a(n_4032), .o(n_4033) );
in01f80 fopt783660 ( .a(n_40306), .o(n_45306) );
ms00f80 delay_add_ln22_unr20_stage8_stallmux_q_reg_27_ ( .ck(newNet_3296), .d(n_32340), .o(delay_add_ln22_unr20_stage8_stallmux_q_27_) );
na02f80 g754554 ( .a(n_26863), .b(n_26862), .o(n_26901) );
no02f80 g753931 ( .a(n_26228), .b(n_25673), .o(n_26265) );
in01f80 g753125 ( .a(n_27423), .o(n_27424) );
in01f80 g736490 ( .a(n_43717), .o(n_43718) );
ms00f80 delay_sub_ln21_0_unr23_stage9_stallmux_q_reg_25_ ( .ck(newNet_2379), .d(n_36520), .o(delay_sub_ln21_0_unr23_stage9_stallmux_q_25_) );
in01f80 FE_OCP_RBC3334_n_44962 ( .a(FE_OCP_RBN3335_n_44962), .o(FE_OCP_RBN3334_n_44962) );
in01f80 fopt783065 ( .a(FE_OFN753_n_44461), .o(n_44463) );
oa12f80 g752012 ( .a(n_28793), .b(n_28396), .c(n_28810), .o(n_28946) );
na02f80 g753834 ( .a(n_26461), .b(n_26393), .o(n_26526) );
na02f80 g755066 ( .a(n_25320), .b(n_25205), .o(n_25380) );
in01f80 g779448 ( .a(n_2070), .o(n_2071) );
na02f80 g742587 ( .a(n_37489), .b(n_37101), .o(n_37532) );
na02f80 g739724 ( .a(n_40505), .b(n_40257), .o(n_40503) );
in01f80 g747215 ( .a(n_32846), .o(n_32847) );
na02f80 g757001 ( .a(n_23345), .b(n_23094), .o(n_23384) );
no02f80 g756858 ( .a(n_23363), .b(delay_add_ln22_unr14_stage6_stallmux_q_10_), .o(n_23407) );
in01f80 g751155 ( .a(n_29821), .o(n_29822) );
in01f80 newInst_3201 ( .a(newNet_3200), .o(newNet_3201) );
ao12f80 g750671 ( .a(n_29340), .b(n_29389), .c(n_29436), .o(n_29513) );
in01f80 newInst_2993 ( .a(newNet_2992), .o(newNet_2993) );
in01f80 g741804 ( .a(n_38344), .o(n_38455) );
in01f80 g740328 ( .a(n_40357), .o(n_40358) );
na02f80 g738150 ( .a(n_42004), .b(n_41793), .o(n_42071) );
na02f80 g772654 ( .a(n_8318), .b(n_7886), .o(n_8319) );
in01f80 g776988 ( .a(n_4147), .o(n_4148) );
in01f80 g771754 ( .a(n_10248), .o(n_10249) );
oa12f80 g745332 ( .a(n_35891), .b(FE_OCP_RBN2995_n_35539), .c(n_35800), .o(n_36164) );
na02f80 g781120 ( .a(n_224), .b(n_143), .o(n_229) );
no02f80 g774710 ( .a(n_6213), .b(n_6485), .o(n_6486) );
na02f80 g737946 ( .a(n_42201), .b(n_42161), .o(n_42341) );
in01f80 FE_OCP_RBC3080_n_16977 ( .a(n_16977), .o(FE_OCP_RBN3080_n_16977) );
in01f80 g752674 ( .a(n_28158), .o(n_28159) );
in01f80 g744048 ( .a(n_35747), .o(n_35698) );
in01f80 FE_RC_489_0 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_16_), .o(FE_RN_144_0) );
in01f80 g780249 ( .a(n_1106), .o(n_1132) );
na02f80 g772889 ( .a(n_7984), .b(n_7937), .o(n_8067) );
in01f80 FE_OCP_RBC1207_n_16814 ( .a(n_16814), .o(FE_OCP_RBN1207_n_16814) );
no02f80 g760650 ( .a(n_20277), .b(n_20256), .o(n_20257) );
ao12f80 g747964 ( .a(n_32724), .b(n_33029), .c(n_32490), .o(n_33128) );
no02f80 g773064 ( .a(n_45887), .b(n_7228), .o(n_7706) );
ao12f80 g745139 ( .a(n_34785), .b(n_34784), .c(n_34783), .o(n_35613) );
no02f80 g744267 ( .a(n_44180), .b(n_34947), .o(n_36133) );
na02f80 g744030 ( .a(n_35550), .b(n_34262), .o(n_35596) );
in01f80 g763257 ( .a(n_17237), .o(n_17238) );
in01f80 g758217 ( .a(n_22850), .o(n_22810) );
in01f80 g762385 ( .a(n_18724), .o(n_18809) );
na02f80 g744834 ( .a(n_35027), .b(n_30612), .o(n_35065) );
na02f80 g748381 ( .a(FE_OCPN1052_n_31674), .b(n_30526), .o(n_31862) );
no02f80 g760741 ( .a(n_19692), .b(n_19624), .o(n_19742) );
in01f80 FE_OCP_RBC3383_n_12365 ( .a(n_12365), .o(FE_OCP_RBN3383_n_12365) );
na02f80 g754201 ( .a(n_26013), .b(n_25989), .o(n_26146) );
na02f80 g740516 ( .a(n_39766), .b(n_39765), .o(n_39767) );
in01f80 g744124 ( .a(n_36262), .o(n_36263) );
in01f80 g766616 ( .a(n_16138), .o(n_16244) );
no02f80 g755117 ( .a(n_25374), .b(n_25316), .o(n_25377) );
na02f80 g742248 ( .a(n_37834), .b(n_37866), .o(n_37918) );
in01f80 g739745 ( .a(delay_add_ln22_unr27_stage10_stallmux_q_17_), .o(n_40756) );
na02f80 g740433 ( .a(n_39728), .b(n_39720), .o(n_39764) );
in01f80 g737484 ( .a(n_42639), .o(n_42599) );
in01f80 g766234 ( .a(n_14464), .o(n_14465) );
no02f80 g769709 ( .a(n_11225), .b(n_11262), .o(n_11358) );
ao12f80 g737292 ( .a(n_42724), .b(n_42889), .c(n_42766), .o(n_42894) );
no02f80 g765043 ( .a(FE_OCP_RBN2742_n_15206), .b(n_14340), .o(n_15285) );
in01f80 FE_OCP_RBC2827_FE_RN_1573_0 ( .a(FE_RN_1573_0), .o(FE_OCP_RBN2827_FE_RN_1573_0) );
na02f80 FE_RC_2507_0 ( .a(FE_RN_1017_0), .b(FE_RN_1018_0), .o(FE_RN_1019_0) );
in01f80 g776201 ( .a(n_4855), .o(n_4856) );
in01f80 FE_RC_2063_0 ( .a(n_45221), .o(FE_RN_700_0) );
in01f80 g768005 ( .a(n_12664), .o(n_12658) );
na02f80 g769266 ( .a(n_11454), .b(n_11407), .o(n_11500) );
na02f80 g741841 ( .a(n_38413), .b(n_38412), .o(n_38414) );
oa22f80 FE_RC_1487_0 ( .a(n_27306), .b(n_27614), .c(n_27305), .d(n_27615), .o(n_27714) );
na02f80 g769878 ( .a(n_11097), .b(n_10920), .o(n_11161) );
in01f80 newInst_3755 ( .a(newNet_2870), .o(newNet_3755) );
no02f80 g745747 ( .a(n_34618), .b(n_34201), .o(n_34682) );
oa12f80 g758823 ( .a(n_21547), .b(n_21546), .c(n_21545), .o(n_21613) );
oa22f80 FE_RC_729_0 ( .a(n_36005), .b(n_36492), .c(FE_OCP_RBN1674_n_36492), .d(n_36004), .o(n_36569) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_16_ ( .ck(newNet_2483), .d(n_32235), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_16_) );
na02f80 g768577 ( .a(n_12146), .b(n_11901), .o(n_12161) );
oa22f80 g739778 ( .a(n_40446), .b(n_40392), .c(n_40447), .d(n_40393), .o(n_40488) );
na02f80 g771690 ( .a(n_8965), .b(FE_OCP_RBN2386_n_8342), .o(n_9201) );
in01f80 FE_OCP_RBC1925_cordic_combinational_sub_ln23_0_unr12_z_0__ ( .a(FE_OCP_RBN1922_cordic_combinational_sub_ln23_0_unr12_z_0__), .o(FE_OCP_RBN1925_cordic_combinational_sub_ln23_0_unr12_z_0__) );
na02f80 g764955 ( .a(n_15504), .b(n_15467), .o(n_15584) );
in01f80 g753198 ( .a(n_27119), .o(n_27230) );
na02f80 g741584 ( .a(n_38665), .b(n_38664), .o(n_38714) );
in01f80 g757857 ( .a(n_22425), .o(n_22390) );
in01f80 g770037 ( .a(n_10955), .o(n_10956) );
oa12f80 g751932 ( .a(n_28758), .b(n_28757), .c(n_28756), .o(n_29172) );
no02f80 g771863 ( .a(n_10122), .b(n_44511), .o(n_10246) );
na02f80 g767469 ( .a(n_13426), .b(n_13425), .o(n_13427) );
in01f80 g767754 ( .a(n_13203), .o(n_13281) );
in01f80 newInst_3298 ( .a(newNet_3297), .o(newNet_3298) );
in01f80 newInst_1066 ( .a(newNet_1065), .o(newNet_1066) );
in01f80 g746162 ( .a(n_33677), .o(n_33695) );
na02f80 g750545 ( .a(FE_OCP_RBN2326_n_29378), .b(FE_RN_1513_0), .o(n_29427) );
in01f80 g745490 ( .a(FE_OCP_RBN2988_n_35539), .o(n_35956) );
na02f80 g754548 ( .a(n_26813), .b(n_26866), .o(n_26946) );
in01f80 g778890 ( .a(n_2277), .o(n_2289) );
in01f80 g775701 ( .a(n_5556), .o(n_5557) );
na02f80 g774986 ( .a(n_6152), .b(n_6133), .o(n_6233) );
ms00f80 delay_xor_ln22_unr3_stage2_stallmux_q_reg_11_ ( .ck(newNet_369), .d(n_44624), .o(delay_xor_ln22_unr3_stage2_stallmux_q_11_) );
in01f80 g749805 ( .a(n_31532), .o(n_31533) );
in01f80 FE_OCPC1528_n_26296 ( .a(FE_OCPN1527_n_26296), .o(FE_OCPN1528_n_26296) );
ao12f80 g779441 ( .a(n_1947), .b(n_1852), .c(delay_xor_ln22_unr3_stage2_stallmux_q_20_), .o(n_1960) );
in01f80 g737879 ( .a(n_42310), .o(n_42280) );
in01f80 g737469 ( .a(n_43070), .o(n_42748) );
in01f80 FE_OFC749_n_45003 ( .a(n_45003), .o(FE_OFN749_n_45003) );
oa12f80 g752455 ( .a(n_27461), .b(n_27672), .c(n_27336), .o(n_27674) );
in01f80 g737907 ( .a(n_42213), .o(n_42214) );
in01f80 g757026 ( .a(n_23833), .o(n_24256) );
na02f80 g743126 ( .a(n_36636), .b(delay_sub_ln21_unr24_stage9_stallmux_q_8_), .o(n_37101) );
na02f80 g773746 ( .a(n_7259), .b(n_7037), .o(n_7335) );
in01f80 g745731 ( .a(n_34396), .o(n_34397) );
na02f80 FE_RC_3583_0 ( .a(FE_RN_1560_0), .b(FE_RN_1561_0), .o(FE_RN_1562_0) );
na02f80 g748424 ( .a(FE_OCPN1052_n_31674), .b(n_30906), .o(n_31759) );
na02f80 g760708 ( .a(FE_OCP_RBN2419_n_19601), .b(FE_OCP_RBN1702_n_19560), .o(n_19664) );
no02f80 g741980 ( .a(n_38008), .b(n_38038), .o(n_38039) );
in01f80 g736903 ( .a(n_43533), .o(n_43534) );
in01f80 g750083 ( .a(n_30969), .o(n_31065) );
ao12f80 g768823 ( .a(n_11996), .b(n_12036), .c(delay_sub_ln21_0_unr8_stage4_stallmux_q_1_), .o(n_12122) );
in01f80 g759819 ( .a(n_21853), .o(n_21854) );
no02f80 g761971 ( .a(n_18964), .b(n_18844), .o(n_18965) );
ao12f80 g769283 ( .a(n_12078), .b(n_45659), .c(delay_sub_ln23_0_unr8_stage4_stallmux_q_28_), .o(n_12710) );
no02f80 g764608 ( .a(n_15917), .b(n_15950), .o(n_16122) );
oa22f80 FE_RC_3342_0 ( .a(n_18551), .b(n_18433), .c(n_18468), .d(n_19893), .o(n_18789) );
na02f80 g768315 ( .a(n_12580), .b(n_11298), .o(n_12640) );
in01f80 newInst_2915 ( .a(newNet_683), .o(newNet_2915) );
na02f80 g755484 ( .a(n_24694), .b(n_22484), .o(n_24690) );
in01f80 newInst_3440 ( .a(newNet_3439), .o(newNet_3440) );
ao22s80 FE_RC_4055_0 ( .a(n_30997), .b(n_31161), .c(n_30998), .d(n_31160), .o(n_31304) );
oa22f80 g752731 ( .a(n_27159), .b(n_27021), .c(n_27158), .d(n_27022), .o(n_27278) );
in01f80 newInst_797 ( .a(newNet_796), .o(newNet_797) );
in01f80 g773165 ( .a(n_7880), .o(n_7954) );
na02f80 g738390 ( .a(n_41680), .b(n_41830), .o(n_41708) );
ao22s80 g780308 ( .a(n_855), .b(n_936), .c(n_922), .d(n_935), .o(n_969) );
no02f80 g779338 ( .a(n_1644), .b(n_1617), .o(n_1691) );
in01f80 newInst_3445 ( .a(newNet_515), .o(newNet_3445) );
na02f80 g759353 ( .a(n_21121), .b(n_45032), .o(n_21147) );
in01f80 g775173 ( .a(n_5769), .o(n_5801) );
in01f80 g737596 ( .a(n_42631), .o(n_42632) );
na02f80 g752578 ( .a(n_28298), .b(n_28278), .o(n_28279) );
oa12f80 g760251 ( .a(n_20222), .b(FE_OCP_RBN3848_FE_RN_1548_0), .c(FE_OCP_RBN3844_FE_RN_1242_0), .o(n_20267) );
no02f80 g763299 ( .a(n_17081), .b(n_16978), .o(n_17134) );
oa12f80 g745468 ( .a(n_34067), .b(n_34167), .c(n_34095), .o(n_34226) );
na02f80 g764383 ( .a(n_16417), .b(n_16361), .o(n_16482) );
in01f80 FE_OCP_RBC3273_n_45224 ( .a(n_45224), .o(FE_OCP_RBN3273_n_45224) );
ms00f80 delay_sub_ln21_0_unr14_stage6_stallmux_q_reg_10_ ( .ck(newNet_2689), .d(n_21920), .o(delay_sub_ln21_0_unr14_stage6_stallmux_q_10_) );
na02f80 g776481 ( .a(n_4252), .b(n_3106), .o(n_4366) );
in01f80 newInst_714 ( .a(newNet_713), .o(newNet_714) );
na02f80 g748066 ( .a(n_31810), .b(n_31666), .o(n_32086) );
no02f80 g761928 ( .a(n_18268), .b(n_17722), .o(n_18595) );
na02f80 g753456 ( .a(n_26957), .b(n_26956), .o(n_27020) );
no02f80 g750554 ( .a(n_29498), .b(FE_OCP_RBN1365_n_29444), .o(n_29543) );
no02f80 g749249 ( .a(n_30630), .b(n_30659), .o(n_30714) );
na02f80 FE_RC_1910_0 ( .a(FE_RN_600_0), .b(n_27888), .o(n_27910) );
no02f80 g744846 ( .a(n_35053), .b(n_30612), .o(n_35080) );
in01f80 FE_RC_1719_0 ( .a(n_28058), .o(FE_RN_474_0) );
no02f80 g767582 ( .a(FE_OCP_RBN2206_n_12907), .b(n_12739), .o(n_12978) );
oa22f80 g739800 ( .a(n_40301), .b(n_40287), .c(n_40302), .d(n_40288), .o(n_40405) );
ao22s80 g780258 ( .a(n_991), .b(FE_OFN794_n_45813), .c(n_992), .d(n_1203), .o(n_1087) );
na02f80 g755293 ( .a(n_25065), .b(n_25064), .o(n_25144) );
in01f80 g746032 ( .a(n_33978), .o(n_33979) );
na02f80 g750738 ( .a(n_29216), .b(FE_OCP_RBN2282_n_29111), .o(n_29269) );
no02f80 g773868 ( .a(n_6997), .b(n_6988), .o(n_6989) );
in01f80 FE_OCP_RBC3718_n_39913 ( .a(FE_OCP_RBN3716_n_39913), .o(FE_OCP_RBN3718_n_39913) );
na02f80 g760514 ( .a(n_19946), .b(n_19965), .o(n_20022) );
in01f80 FE_OCP_RBC3487_n_2438 ( .a(FE_OCP_RBN2293_n_2438), .o(FE_OCP_RBN3487_n_2438) );
na02f80 g756338 ( .a(n_24002), .b(n_24001), .o(n_24003) );
in01f80 FE_RC_1986_0 ( .a(n_13204), .o(FE_RN_647_0) );
in01f80 g761872 ( .a(n_18370), .o(n_18371) );
na02f80 g759065 ( .a(n_21230), .b(n_21229), .o(n_21391) );
in01f80 newInst_268 ( .a(newNet_240), .o(newNet_268) );
in01f80 FE_OCP_RBC2620_n_44561 ( .a(FE_OCP_RBN3594_n_44561), .o(FE_OCP_RBN2620_n_44561) );
no02f80 g765880 ( .a(n_14818), .b(n_14801), .o(n_14858) );
in01f80 g753615 ( .a(delay_sub_ln21_0_unr17_stage7_stallmux_q_3_), .o(n_28115) );
no02f80 g769369 ( .a(n_45685), .b(delay_sub_ln23_0_unr8_stage4_stallmux_q_26_), .o(n_12080) );
no02f80 g767786 ( .a(n_46933), .b(delay_add_ln22_unr8_stage4_stallmux_q_25_), .o(n_12932) );
in01f80 newInst_1490 ( .a(newNet_26), .o(newNet_1490) );
oa12f80 g780749 ( .a(n_426), .b(n_584), .c(n_404), .o(n_590) );
no02f80 g755500 ( .a(n_24778), .b(n_24564), .o(n_24800) );
no02f80 g744795 ( .a(n_35194), .b(n_30587), .o(n_35197) );
in01f80 g775779 ( .a(n_5626), .o(n_5582) );
na02f80 g773072 ( .a(n_7891), .b(n_7857), .o(n_7892) );
no02f80 g768060 ( .a(n_12881), .b(n_12135), .o(n_12958) );
ao12f80 g779020 ( .a(n_2064), .b(n_2063), .c(n_2062), .o(n_2858) );
in01f80 g766396 ( .a(n_14397), .o(n_15518) );
in01f80 newInst_2461 ( .a(newNet_1587), .o(newNet_2461) );
in01f80 g771478 ( .a(n_8941), .o(n_8942) );
in01f80 FE_OCP_RBC3828_n_19204 ( .a(n_19204), .o(FE_OCP_RBN3828_n_19204) );
no02f80 g784415 ( .a(n_46197), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_27_), .o(n_46227) );
no02f80 g747238 ( .a(n_32617), .b(n_32548), .o(n_32627) );
ao12f80 g754471 ( .a(n_25630), .b(n_25629), .c(n_25628), .o(n_25789) );
no02f80 g762194 ( .a(n_18113), .b(n_18137), .o(n_18174) );
in01f80 g771114 ( .a(delay_add_ln22_unr8_stage4_stallmux_q_1_), .o(n_11871) );
in01f80 g742400 ( .a(n_37791), .o(n_37792) );
ao12f80 g738975 ( .a(n_40768), .b(n_41204), .c(n_40858), .o(n_41267) );
in01f80 g737884 ( .a(n_42608), .o(n_42609) );
na02f80 g739303 ( .a(n_45155), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .o(n_40971) );
no02f80 g779301 ( .a(n_1705), .b(n_1712), .o(n_1733) );
in01f80 FE_OCP_RBC2968_n_26398 ( .a(n_26398), .o(FE_OCP_RBN2968_n_26398) );
no02f80 g738583 ( .a(n_41807), .b(n_41457), .o(n_41864) );
oa12f80 g778300 ( .a(n_2519), .b(n_2528), .c(n_2518), .o(n_3361) );
na02f80 g770033 ( .a(n_10922), .b(FE_OCP_RBN3643_n_44490), .o(n_10995) );
no02f80 g775832 ( .a(n_5493), .b(n_47015), .o(n_5516) );
no02f80 g771596 ( .a(n_10284), .b(n_10283), .o(n_10285) );
in01f80 g743130 ( .a(n_37038), .o(n_37039) );
na03f80 FE_RC_1665_0 ( .a(n_29487), .b(n_29023), .c(n_29488), .o(n_29489) );
no02f80 FE_RC_939_0 ( .a(n_22383), .b(n_22569), .o(FE_RN_277_0) );
in01f80 g755695 ( .a(n_24553), .o(n_24554) );
in01f80 FE_OCP_RBC3017_n_31117 ( .a(FE_OCP_RBN3014_n_31117), .o(FE_OCP_RBN3017_n_31117) );
na02f80 g758751 ( .a(n_21684), .b(n_21654), .o(n_21685) );
na02f80 g753999 ( .a(n_26180), .b(n_26210), .o(n_26361) );
na02f80 g753234 ( .a(n_27167), .b(FE_OCP_RBN2939_n_26276), .o(n_27296) );
in01f80 g746731 ( .a(n_34738), .o(n_34229) );
in01f80 FE_RC_3527_0 ( .a(FE_RN_1525_0), .o(n_23330) );
no02f80 g741315 ( .a(FE_OCP_RBN2548_n_44944), .b(n_38872), .o(n_38901) );
in01f80 FE_OCP_RBC1926_cordic_combinational_sub_ln23_0_unr12_z_0__ ( .a(cordic_combinational_sub_ln23_0_unr12_z_0_), .o(FE_OCP_RBN1926_cordic_combinational_sub_ln23_0_unr12_z_0__) );
no02f80 FE_RC_1037_0 ( .a(FE_RN_297_0), .b(FE_RN_298_0), .o(FE_RN_299_0) );
na02f80 g762319 ( .a(n_18077), .b(delay_sub_ln21_0_unr11_stage5_stallmux_q_12_), .o(n_18136) );
na02f80 g770323 ( .a(n_10663), .b(FE_OCPN955_n_44460), .o(n_10690) );
na02f80 g766539 ( .a(n_13954), .b(n_13375), .o(n_13999) );
no02f80 g739445 ( .a(n_44804), .b(delay_sub_ln21_0_unr27_stage10_stallmux_q_26_), .o(n_40850) );
no02f80 g743108 ( .a(FE_OCP_RBN3354_delay_sub_ln21_unr24_stage9_stallmux_q_8_), .b(delay_sub_ln21_0_unr23_stage9_stallmux_q_20_), .o(n_37098) );
in01f80 FE_RC_3318_0 ( .a(FE_RN_1460_0), .o(FE_RN_1459_0) );
in01f80 FE_RC_2394_0 ( .a(n_42112), .o(FE_RN_940_0) );
na02f80 g773882 ( .a(n_7083), .b(n_6695), .o(n_7084) );
na02f80 g775458 ( .a(n_5641), .b(n_5720), .o(n_5771) );
in01f80 FE_OCP_RBC3830_n_19204 ( .a(FE_OCP_RBN3829_n_19204), .o(FE_OCP_RBN3830_n_19204) );
in01f80 FE_OCPC972_n_15900 ( .a(n_15900), .o(FE_OCPN972_n_15900) );
no02f80 g764263 ( .a(n_16438), .b(n_16461), .o(n_16486) );
no02f80 g777103 ( .a(n_3604), .b(n_3650), .o(n_3760) );
no02f80 g748602 ( .a(n_31305), .b(n_31157), .o(n_31337) );
in01f80 g770439 ( .a(n_10712), .o(n_10630) );
in01f80 g740167 ( .a(n_40001), .o(n_40002) );
na02f80 g757357 ( .a(n_23100), .b(delay_add_ln22_unr14_stage6_stallmux_q_3_), .o(n_23187) );
na02f80 g741695 ( .a(n_38564), .b(n_38562), .o(n_38563) );
in01f80 FE_OCP_RBC2246_n_13017 ( .a(FE_OCP_RBN2243_n_13017), .o(FE_OCP_RBN2246_n_13017) );
in01f80 newInst_1464 ( .a(newNet_773), .o(newNet_1464) );
na02f80 g740917 ( .a(n_39256), .b(n_39300), .o(n_39370) );
na02f80 g753163 ( .a(n_27342), .b(n_27387), .o(n_27482) );
in01f80 g758934 ( .a(n_21429), .o(n_21542) );
no02f80 g744141 ( .a(n_35736), .b(n_35659), .o(n_35688) );
in01f80 newInst_605 ( .a(newNet_604), .o(newNet_605) );
na02f80 g741527 ( .a(n_38742), .b(n_38725), .o(n_38756) );
in01f80 newInst_3179 ( .a(newNet_503), .o(newNet_3179) );
in01f80 newInst_1843 ( .a(newNet_1842), .o(newNet_1843) );
in01f80 newInst_1049 ( .a(newNet_1048), .o(newNet_1049) );
na03f80 g761537 ( .a(n_18759), .b(n_18718), .c(n_18366), .o(n_18799) );
in01f80 FE_OCP_RBC2249_n_13017 ( .a(FE_OCP_RBN2247_n_13017), .o(FE_OCP_RBN2249_n_13017) );
in01f80 FE_OCP_RBC1158_n_18517 ( .a(n_18517), .o(FE_OCP_RBN1158_n_18517) );
in01f80 FE_RC_2326_0 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_15_), .o(FE_RN_886_0) );
in01f80 g759914 ( .a(n_21297), .o(n_21377) );
oa12f80 g776083 ( .a(n_4666), .b(n_4656), .c(n_4804), .o(n_4878) );
in01f80 g753915 ( .a(n_26291), .o(n_26290) );
na02f80 g748817 ( .a(n_32457), .b(n_32484), .o(n_32837) );
in01f80 g777890 ( .a(n_4761), .o(n_3195) );
in01f80 g753001 ( .a(n_27469), .o(n_27507) );
no02f80 g754222 ( .a(n_25932), .b(FE_OCP_DRV_N3745_FE_OFN737_n_22641), .o(n_25993) );
oa12f80 g762123 ( .a(n_18175), .b(n_18174), .c(n_18173), .o(n_18205) );
na02f80 g744547 ( .a(n_35368), .b(n_35367), .o(n_35410) );
no02f80 g741879 ( .a(n_38244), .b(n_44034), .o(n_38287) );
in01f80 fopt782831 ( .a(n_35550), .o(n_44256) );
in01f80 g772411 ( .a(n_8670), .o(n_8671) );
in01f80 g774735 ( .a(delay_sub_ln21_0_unr5_stage3_stallmux_q_24_), .o(n_7521) );
na03f80 FE_RC_75_0 ( .a(n_17848), .b(n_17894), .c(n_17827), .o(n_17895) );
no02f80 g776786 ( .a(n_4114), .b(n_4046), .o(n_4310) );
na02f80 g741627 ( .a(n_38592), .b(n_38778), .o(n_38613) );
no02f80 g770609 ( .a(n_10270), .b(n_44464), .o(n_10286) );
ms00f80 delay_sub_ln21_0_unr20_stage8_stallmux_q_reg_2_ ( .ck(newNet_2449), .d(n_31193), .o(delay_sub_ln21_0_unr20_stage8_stallmux_q_2_) );
no02f80 g747242 ( .a(n_32655), .b(n_32654), .o(n_32718) );
no02f80 g776369 ( .a(n_4735), .b(n_4650), .o(n_4890) );
no02f80 g767820 ( .a(n_12768), .b(n_12247), .o(n_12769) );
in01f80 g742910 ( .a(n_37120), .o(n_37121) );
na02f80 g753307 ( .a(n_27110), .b(n_25827), .o(n_27139) );
no02f80 g757059 ( .a(n_23643), .b(n_23642), .o(n_23644) );
ao12f80 g739151 ( .a(n_40693), .b(n_40897), .c(n_40742), .o(n_40915) );
na03f80 g743878 ( .a(n_37022), .b(n_37020), .c(n_36916), .o(n_37136) );
na02f80 g779344 ( .a(n_1625), .b(delay_add_ln22_unr2_stage2_stallmux_q_2_), .o(n_1652) );
oa22f80 g771559 ( .a(n_9234), .b(n_9128), .c(n_9235), .d(n_9127), .o(n_9441) );
no02f80 g765561 ( .a(n_15142), .b(n_14224), .o(n_15216) );
na02f80 g742739 ( .a(n_37439), .b(n_37438), .o(n_37440) );
no02f80 g750054 ( .a(n_29869), .b(n_29082), .o(n_29960) );
ao12f80 g757716 ( .a(n_22171), .b(n_22450), .c(n_22139), .o(n_22542) );
no02f80 g737272 ( .a(n_42918), .b(n_42440), .o(n_42905) );
na02f80 g763962 ( .a(n_16569), .b(n_16537), .o(n_16645) );
no02f80 g744549 ( .a(n_35368), .b(FE_OCPN1516_n_35367), .o(n_35385) );
in01f80 g771276 ( .a(n_9657), .o(n_9658) );
ao12f80 g772288 ( .a(n_8708), .b(n_8707), .c(n_8706), .o(n_9939) );
ao22s80 g752355 ( .a(FE_OCP_RBN3364_n_44722), .b(n_44422), .c(n_44420), .d(FE_OCP_RBN3306_n_44722), .o(n_27859) );
na02f80 g776553 ( .a(n_4112), .b(n_4167), .o(n_4317) );
in01f80 g746920 ( .a(n_33231), .o(n_33232) );
na02f80 g741840 ( .a(n_38416), .b(n_38415), .o(n_38417) );
oa12f80 g739082 ( .a(n_41095), .b(n_41108), .c(n_41094), .o(n_41126) );
na02f80 g778402 ( .a(n_2412), .b(n_2538), .o(n_2604) );
no02f80 g736739 ( .a(n_43357), .b(n_43356), .o(n_43358) );
ao12f80 g737638 ( .a(n_42467), .b(n_42392), .c(n_42421), .o(n_42760) );
no02f80 g744870 ( .a(n_35030), .b(n_35055), .o(n_35143) );
in01f80 FE_RC_2886_0 ( .a(n_13515), .o(FE_RN_1249_0) );
oa12f80 g758729 ( .a(n_21542), .b(n_21558), .c(n_21661), .o(n_21686) );
in01f80 g757646 ( .a(delay_xor_ln21_unr15_stage6_stallmux_q_2_), .o(n_22795) );
no02f80 g768587 ( .a(n_12242), .b(n_12241), .o(n_12243) );
na02f80 g775291 ( .a(n_5644), .b(n_4556), .o(n_5667) );
in01f80 newInst_1940 ( .a(newNet_1939), .o(newNet_1940) );
ao12f80 g774380 ( .a(n_6815), .b(n_6624), .c(delay_sub_ln23_0_unr5_stage3_stallmux_q_30_), .o(n_7623) );
no02f80 g755043 ( .a(n_25293), .b(n_25295), .o(n_25296) );
in01f80 g756038 ( .a(n_24997), .o(n_25055) );
oa12f80 g741871 ( .a(n_38381), .b(n_38380), .c(n_38379), .o(n_38862) );
in01f80 g746663 ( .a(n_34666), .o(n_34810) );
na02f80 g781058 ( .a(cos_out_8), .b(FE_OFN2_n_43918), .o(n_313) );
oa12f80 g767365 ( .a(n_13603), .b(n_13620), .c(n_13602), .o(n_13649) );
na02f80 g746790 ( .a(n_33200), .b(n_33150), .o(n_33201) );
in01f80 g743287 ( .a(n_36757), .o(n_36758) );
oa22f80 FE_RC_3720_0 ( .a(n_5782), .b(n_5975), .c(n_5779), .d(n_5974), .o(n_6074) );
in01f80 newInst_381 ( .a(newNet_209), .o(newNet_381) );
na02f80 g744135 ( .a(n_35615), .b(FE_OCPN1422_n_35611), .o(n_35612) );
in01f80 g745426 ( .a(n_35715), .o(n_35716) );
in01f80 g741773 ( .a(n_38471), .o(n_38472) );
no02f80 g769644 ( .a(n_11358), .b(n_11357), .o(n_11383) );
oa12f80 g739396 ( .a(n_45145), .b(delay_add_ln22_unr27_stage10_stallmux_q_8_), .c(delay_add_ln22_unr27_stage10_stallmux_q_9_), .o(n_40687) );
in01f80 FE_OCP_RBC2786_n_15079 ( .a(n_15079), .o(FE_OCP_RBN2786_n_15079) );
oa22f80 g784555 ( .a(FE_OFN801_n_46285), .b(n_11278), .c(FE_OCP_RBN3044_n_46337), .d(n_11232), .o(n_46376) );
na02f80 g745839 ( .a(n_44102), .b(FE_OCP_RBN2269_n_33803), .o(n_34238) );
in01f80 g738699 ( .a(n_41534), .o(n_41535) );
in01f80 g759696 ( .a(n_20640), .o(n_20723) );
in01f80 newInst_2546 ( .a(newNet_2545), .o(newNet_2546) );
no02f80 g762609 ( .a(n_18040), .b(n_17951), .o(n_18086) );
no02f80 g770287 ( .a(n_10718), .b(n_9956), .o(n_10869) );
na02f80 g771147 ( .a(n_9788), .b(n_8239), .o(n_9843) );
no02f80 g762265 ( .a(n_18766), .b(n_18585), .o(n_19541) );
in01f80 newInst_2524 ( .a(newNet_2523), .o(newNet_2524) );
na02f80 g756906 ( .a(n_23347), .b(delay_sub_ln21_0_unr14_stage6_stallmux_q_9_), .o(n_23374) );
no02f80 g746179 ( .a(n_33647), .b(n_34037), .o(n_33693) );
oa12f80 g755906 ( .a(n_25030), .b(n_25160), .c(n_25090), .o(n_25579) );
no02f80 g770409 ( .a(n_10483), .b(n_44463), .o(n_10547) );
na02f80 g772366 ( .a(n_8572), .b(n_7941), .o(n_8682) );
na02f80 g742029 ( .a(n_38050), .b(FE_OCP_RBN3426_n_44881), .o(n_38138) );
no02f80 g750074 ( .a(n_29896), .b(n_30192), .o(n_30262) );
ao12f80 g773656 ( .a(n_7324), .b(n_7323), .c(n_7322), .o(n_7376) );
no02f80 g776043 ( .a(n_47005), .b(FE_OCP_RBN2534_n_47018), .o(n_5032) );
ao12f80 g768518 ( .a(n_12332), .b(n_12331), .c(n_12341), .o(n_13330) );
no02f80 g742560 ( .a(n_37619), .b(n_37618), .o(n_37617) );
ao12f80 g761840 ( .a(n_18127), .b(n_18318), .c(n_18126), .o(n_18475) );
na02f80 g748793 ( .a(n_32586), .b(n_32457), .o(n_32458) );
in01f80 g778138 ( .a(n_2967), .o(n_2968) );
in01f80 g740064 ( .a(n_40114), .o(n_40115) );
na02f80 g756431 ( .a(n_23770), .b(n_23757), .o(n_23824) );
in01f80 g771577 ( .a(FE_OCP_RBN2529_n_9044), .o(n_9121) );
na02f80 g759638 ( .a(n_20720), .b(n_45066), .o(n_20911) );
in01f80 g772979 ( .a(n_7834), .o(n_7863) );
in01f80 g770527 ( .a(n_10401), .o(n_10437) );
na02f80 g754114 ( .a(n_26021), .b(FE_OCPN1530_n_26090), .o(n_26369) );
na02f80 g749494 ( .a(n_30452), .b(n_30199), .o(n_30467) );
no02f80 FE_RC_3592_0 ( .a(FE_RN_1567_0), .b(n_14478), .o(n_14515) );
na02f80 g767017 ( .a(n_14210), .b(n_13650), .o(n_14295) );
oa12f80 g767596 ( .a(n_12943), .b(n_12949), .c(n_12942), .o(n_13052) );
oa12f80 g774975 ( .a(FE_OCP_RBN3047_n_6013), .b(n_6090), .c(n_6089), .o(n_6115) );
na02f80 g744616 ( .a(n_35324), .b(FE_OCP_DRV_N1578_n_33904), .o(n_35360) );
in01f80 g740708 ( .a(n_39597), .o(n_39598) );
in01f80 FE_OCP_RBC3736_n_27535 ( .a(n_27535), .o(FE_OCP_RBN3736_n_27535) );
no02f80 g745412 ( .a(n_35543), .b(n_35542), .o(n_35605) );
oa22f80 g752850 ( .a(n_27285), .b(n_27923), .c(n_27948), .d(delay_sub_ln23_0_unr20_stage7_stallmux_q_17_), .o(n_28558) );
na02f80 g766931 ( .a(n_13901), .b(n_13898), .o(n_14307) );
na02f80 g768022 ( .a(n_12910), .b(n_12887), .o(n_13248) );
ao12f80 g773725 ( .a(n_7191), .b(n_7194), .c(n_7190), .o(n_7237) );
oa12f80 g772759 ( .a(n_8094), .b(n_8155), .c(n_7802), .o(n_8258) );
in01f80 FE_OCP_RBC2843_n_10326 ( .a(n_10326), .o(FE_OCP_RBN2843_n_10326) );
no03m80 g748774 ( .a(n_32499), .b(n_32498), .c(n_32391), .o(n_32500) );
na02f80 g739252 ( .a(n_40856), .b(n_40772), .o(n_40857) );
no02f80 g765281 ( .a(n_15873), .b(n_15876), .o(n_15877) );
ao12f80 g761523 ( .a(n_18920), .b(n_18948), .c(n_18919), .o(n_19028) );
in01f80 newInst_2761 ( .a(newNet_2760), .o(newNet_2761) );
na02f80 g778482 ( .a(n_2878), .b(n_2759), .o(n_2882) );
in01f80 newInst_439 ( .a(newNet_438), .o(newNet_439) );
no02f80 g744903 ( .a(n_36420), .b(n_36419), .o(n_36463) );
ao12f80 g751024 ( .a(n_29837), .b(n_29945), .c(n_29938), .o(n_29946) );
no02f80 g775670 ( .a(n_5709), .b(n_5577), .o(n_5598) );
no02f80 g745825 ( .a(n_44133), .b(n_33673), .o(n_34201) );
no02f80 g740854 ( .a(n_39347), .b(n_39278), .o(n_39348) );
in01f80 g759472 ( .a(n_20973), .o(n_20937) );
na02f80 g736557 ( .a(n_43532), .b(n_43111), .o(n_43629) );
na02f80 g755147 ( .a(n_25105), .b(n_25047), .o(n_25157) );
oa22f80 g764134 ( .a(n_16821), .b(n_15962), .c(n_16820), .d(n_15963), .o(n_16927) );
in01f80 g748723 ( .a(n_31160), .o(n_31161) );
in01f80 newInst_209 ( .a(newNet_208), .o(newNet_209) );
in01f80 g742858 ( .a(n_37188), .o(n_37165) );
ao12f80 g779466 ( .a(n_1832), .b(n_1800), .c(delay_xor_ln21_unr3_stage2_stallmux_q_16_), .o(n_1854) );
ao12f80 g751621 ( .a(n_28371), .b(n_28391), .c(n_28293), .o(n_28426) );
na02f80 g750433 ( .a(n_29577), .b(n_29576), .o(n_29592) );
no02f80 g742966 ( .a(n_37082), .b(n_36610), .o(n_37126) );
na02f80 g770789 ( .a(n_10136), .b(n_10091), .o(n_10309) );
in01f80 FE_OCPC3747_n_29439 ( .a(FE_OCPN3746_n_29439), .o(FE_OCPN3747_n_29439) );
in01f80 FE_OCP_DRV_C1612_n_21706 ( .a(FE_OCP_DRV_N1611_n_21706), .o(FE_OCP_DRV_N1612_n_21706) );
no03m80 FE_RC_3684_0 ( .a(n_23308), .b(FE_RN_1618_0), .c(FE_OCPN1022_n_23195), .o(n_23312) );
na02f80 g748523 ( .a(n_31467), .b(n_31425), .o(n_31497) );
in01f80 g759577 ( .a(n_20621), .o(n_20622) );
no02f80 g759713 ( .a(n_20504), .b(n_45101), .o(n_20546) );
no02f80 g760471 ( .a(n_20624), .b(n_19982), .o(n_20655) );
oa12f80 g748016 ( .a(n_32485), .b(n_44347), .c(n_32414), .o(n_33046) );
oa12f80 g780696 ( .a(n_488), .b(n_646), .c(n_480), .o(n_653) );
na02f80 g761912 ( .a(n_18268), .b(n_17696), .o(n_18742) );
na02f80 g737684 ( .a(n_42367), .b(n_42459), .o(n_42460) );
no02f80 g749368 ( .a(n_30692), .b(n_29228), .o(n_30758) );
oa12f80 g780740 ( .a(n_595), .b(n_594), .c(n_593), .o(n_734) );
in01f80 FE_RC_2628_0 ( .a(n_12056), .o(FE_RN_1094_0) );
oa12f80 g754750 ( .a(n_25209), .b(n_25366), .c(n_25154), .o(n_25404) );
in01f80 g759778 ( .a(n_21715), .o(n_21716) );
in01f80 newInst_2208 ( .a(newNet_2207), .o(newNet_2208) );
na02f80 g754900 ( .a(FE_OCP_RBN2597_n_25181), .b(n_24332), .o(n_25301) );
no02f80 g761695 ( .a(n_19405), .b(n_18737), .o(n_19496) );
oa22f80 FE_RC_369_0 ( .a(n_12755), .b(n_13267), .c(n_12756), .d(n_13266), .o(n_13453) );
in01f80 newInst_3182 ( .a(newNet_3181), .o(newNet_3182) );
no02f80 g767766 ( .a(n_13084), .b(delay_sub_ln21_0_unr8_stage4_stallmux_q_29_), .o(n_13371) );
na02f80 g742673 ( .a(n_37372), .b(n_37135), .o(n_37465) );
na02f80 g767899 ( .a(n_12990), .b(FE_OCPN860_n_12880), .o(n_13065) );
na02f80 g743044 ( .a(n_37044), .b(n_37161), .o(n_37438) );
no02f80 g757565 ( .a(n_22817), .b(n_22796), .o(n_22927) );
in01f80 newInst_655 ( .a(newNet_654), .o(newNet_655) );
ao22s80 FE_RC_810_0 ( .a(n_44352), .b(n_7520), .c(n_7519), .d(n_44351), .o(n_8380) );
in01f80 FE_OCP_RBC1344_n_32520 ( .a(n_32520), .o(FE_OCP_RBN1344_n_32520) );
na02f80 FE_RC_3972_0 ( .a(n_24553), .b(n_24556), .o(FE_RN_1720_0) );
no02f80 g764168 ( .a(n_16474), .b(FE_OCP_RBN2679_n_14768), .o(n_16498) );
in01f80 g744496 ( .a(n_35475), .o(n_35443) );
na02f80 g766994 ( .a(n_13531), .b(n_47253), .o(n_13582) );
na02f80 g769114 ( .a(n_11626), .b(n_11671), .o(n_11803) );
in01f80 newInst_2747 ( .a(newNet_2746), .o(newNet_2747) );
in01f80 g750148 ( .a(n_30071), .o(n_30072) );
na02f80 g763194 ( .a(n_17340), .b(delay_add_ln22_unr11_stage5_stallmux_q_3_), .o(n_17477) );
na02f80 g747256 ( .a(n_32693), .b(n_32692), .o(n_32694) );
oa12f80 g737257 ( .a(n_42486), .b(n_42857), .c(n_42549), .o(n_42907) );
in01f80 g773447 ( .a(n_7542), .o(n_7579) );
in01f80 g780422 ( .a(n_1079), .o(n_853) );
in01f80 g779557 ( .a(n_2113), .o(n_2114) );
in01f80 g757112 ( .a(n_24059), .o(n_27845) );
oa22f80 FE_RC_3914_0 ( .a(n_22299), .b(n_22556), .c(n_22335), .d(FE_OCP_RBN1852_n_22556), .o(n_22709) );
ao12f80 g755149 ( .a(n_24695), .b(n_24989), .c(n_24690), .o(n_25071) );
in01f80 FE_RC_1837_0 ( .a(n_23074), .o(FE_RN_554_0) );
ms00f80 delay_sub_ln23_0_unr2_stage2_stallmux_q_reg_25_ ( .ck(newNet_1309), .d(n_1273), .o(delay_sub_ln23_0_unr2_stage2_stallmux_q_25_) );
in01f80 g756622 ( .a(n_23666), .o(n_23602) );
no02f80 g764587 ( .a(n_16000), .b(n_15984), .o(n_16076) );
na02f80 g749728 ( .a(n_31428), .b(n_31511), .o(n_31537) );
oa22f80 FE_RC_1471_0 ( .a(n_24350), .b(n_27739), .c(n_27796), .d(n_27730), .o(n_27779) );
oa22f80 g752519 ( .a(n_27628), .b(n_27495), .c(n_27629), .d(n_27494), .o(n_27726) );
in01f80 FE_OCPC1420_n_14003 ( .a(FE_OCPN1419_n_14003), .o(FE_OCPN1420_n_14003) );
in01f80 g741211 ( .a(n_38831), .o(n_38832) );
in01f80 g750745 ( .a(n_29279), .o(n_29234) );
na02f80 g758287 ( .a(FE_OCPN992_n_22249), .b(n_20862), .o(n_22374) );
in01f80 g739515 ( .a(n_40709), .o(n_40710) );
in01f80 newInst_1966 ( .a(newNet_1965), .o(newNet_1966) );
in01f80 g777222 ( .a(n_3832), .o(n_3833) );
no02f80 FE_RC_3497_0 ( .a(FE_RN_1508_0), .b(n_31908), .o(n_31959) );
in01f80 g742908 ( .a(n_37122), .o(n_37123) );
na02f80 FE_RC_400_0 ( .a(FE_RN_119_0), .b(n_15475), .o(n_46982) );
no02f80 g775632 ( .a(n_47001), .b(n_5603), .o(n_5638) );
no02f80 g758142 ( .a(n_22461), .b(n_22370), .o(n_22462) );
no02f80 g742794 ( .a(n_37277), .b(n_37099), .o(n_37316) );
in01f80 FE_RC_3169_0 ( .a(n_22482), .o(FE_RN_1403_0) );
na02f80 g760285 ( .a(FE_OCP_RBN3613_n_20249), .b(n_19347), .o(n_20608) );
oa12f80 g743657 ( .a(n_35917), .b(n_36329), .c(n_35739), .o(n_36378) );
na02f80 g740109 ( .a(n_40071), .b(n_40179), .o(n_40279) );
no02f80 g757037 ( .a(n_23743), .b(n_23903), .o(n_23981) );
in01f80 FE_OCP_RBC3452_n_37945 ( .a(FE_OCP_RBN3450_n_37945), .o(FE_OCP_RBN3452_n_37945) );
in01f80 FE_OCP_RBC2527_n_3421 ( .a(FE_OCP_RBN2526_n_3421), .o(FE_OCP_RBN2527_n_3421) );
in01f80 g739292 ( .a(n_40846), .o(n_40847) );
ao12f80 g757526 ( .a(n_22313), .b(n_22720), .c(n_22214), .o(n_22719) );
no02f80 g771697 ( .a(n_8848), .b(n_8794), .o(n_8911) );
no02f80 g763696 ( .a(n_17266), .b(n_17210), .o(n_17430) );
in01f80 g771320 ( .a(n_9091), .o(n_9092) );
in01f80 g764725 ( .a(n_15951), .o(n_15898) );
oa12f80 g742945 ( .a(n_36897), .b(n_36995), .c(n_36878), .o(n_37058) );
oa12f80 g782662 ( .a(FE_OCP_RBN3552_n_44575), .b(n_9035), .c(n_9034), .o(n_44055) );
no02f80 g772779 ( .a(n_7944), .b(n_7414), .o(n_7990) );
ao12f80 g752834 ( .a(n_28175), .b(n_27948), .c(delay_sub_ln23_0_unr20_stage7_stallmux_q_23_), .o(n_28692) );
no02f80 FE_RC_4231_0 ( .a(FE_RN_1857_0), .b(FE_OCP_RBN1222_n_45522), .o(n_15415) );
oa12f80 g775860 ( .a(n_4577), .b(n_5193), .c(n_4460), .o(n_5339) );
no02f80 g780793 ( .a(n_422), .b(n_419), .o(n_423) );
na02f80 g737919 ( .a(n_42547), .b(n_42271), .o(n_42581) );
ao22s80 g737365 ( .a(n_42779), .b(n_42729), .c(n_42778), .d(n_42728), .o(n_42829) );
in01f80 g768095 ( .a(n_12615), .o(n_12627) );
no02f80 g760311 ( .a(n_20151), .b(n_20043), .o(n_20173) );
in01f80 g753969 ( .a(n_26354), .o(n_26387) );
oa12f80 g756945 ( .a(n_24025), .b(n_24188), .c(n_23985), .o(n_24513) );
na02f80 g749128 ( .a(n_30849), .b(FE_OCPN1410_n_27014), .o(n_30879) );
in01f80 g761620 ( .a(n_19609), .o(n_19569) );
in01f80 g749847 ( .a(n_31088), .o(n_31089) );
na02f80 g750772 ( .a(n_29259), .b(n_29293), .o(n_29392) );
in01f80 g764773 ( .a(delay_add_ln22_unr11_stage5_stallmux_q_7_), .o(n_15892) );
na02f80 g765271 ( .a(n_14991), .b(FE_OCP_RBN2507_n_13896), .o(n_15025) );
in01f80 newInst_1954 ( .a(newNet_1953), .o(newNet_1954) );
na02f80 g767009 ( .a(n_14210), .b(n_13715), .o(n_14386) );
na02f80 g750313 ( .a(n_29718), .b(n_29696), .o(n_29788) );
ao22s80 g743566 ( .a(n_37586), .b(n_36869), .c(n_37517), .d(n_36868), .o(n_37613) );
in01f80 g773890 ( .a(n_7022), .o(n_7023) );
no02f80 g766669 ( .a(n_13690), .b(n_13782), .o(n_13840) );
no02f80 g761765 ( .a(n_19293), .b(n_19292), .o(n_19294) );
no02f80 g740380 ( .a(n_39803), .b(n_39881), .o(n_39882) );
na02f80 g750412 ( .a(n_29579), .b(n_29554), .o(n_29628) );
no02f80 g776177 ( .a(n_4654), .b(FE_OCP_RBN2691_FE_OCPN843_n_3912), .o(n_4842) );
in01f80 newInst_246 ( .a(newNet_245), .o(newNet_246) );
no02f80 g751910 ( .a(n_28863), .b(n_28901), .o(n_28882) );
oa12f80 g772549 ( .a(n_8373), .b(n_8372), .c(n_8371), .o(n_9381) );
no02f80 g754723 ( .a(FE_OCP_RBN2965_n_26231), .b(n_26604), .o(n_26637) );
na02f80 g773759 ( .a(n_7156), .b(delay_add_ln22_unr5_stage3_stallmux_q_14_), .o(n_7225) );
ao12f80 g775934 ( .a(n_4949), .b(n_5020), .c(n_4935), .o(n_5283) );
in01f80 newInst_3195 ( .a(newNet_3194), .o(newNet_3195) );
na02f80 g774588 ( .a(n_6331), .b(n_6386), .o(n_6387) );
no02f80 g768548 ( .a(n_12312), .b(n_11946), .o(n_12339) );
in01f80 g756884 ( .a(n_23988), .o(n_24029) );
in01f80 g739638 ( .a(delay_sub_ln21_0_unr27_stage10_stallmux_q_27_), .o(n_40573) );
no02f80 g750121 ( .a(FE_OCP_RBN3562_n_29857), .b(n_29231), .o(n_30212) );
in01f80 newInst_3630 ( .a(newNet_3629), .o(newNet_3630) );
in01f80 g770712 ( .a(n_10379), .o(n_10428) );
in01f80 g751562 ( .a(n_28722), .o(n_28672) );
in01f80 g778095 ( .a(n_3055), .o(n_3054) );
oa22f80 g747547 ( .a(n_32255), .b(n_32287), .c(n_32240), .d(n_28336), .o(n_32289) );
in01f80 FE_OCPC948_n_41382 ( .a(FE_OCPN947_n_41382), .o(FE_OCPN948_n_41382) );
na02f80 g755621 ( .a(n_24465), .b(n_24367), .o(n_24507) );
oa12f80 g784632 ( .a(n_27920), .b(n_27919), .c(n_27839), .o(n_46961) );
in01f80 g773213 ( .a(n_8038), .o(n_7993) );
in01f80 FE_OCP_RBC2621_n_44561 ( .a(FE_OCP_RBN2620_n_44561), .o(FE_OCP_RBN2621_n_44561) );
na02f80 g749303 ( .a(n_30681), .b(n_27131), .o(n_30744) );
in01f80 g769197 ( .a(n_11632), .o(n_11633) );
in01f80 FE_OCP_RBC2878_n_15553 ( .a(n_15553), .o(FE_OCP_RBN2878_n_15553) );
no02f80 g747381 ( .a(FE_OCP_RBN2103_n_44962), .b(delay_xor_ln22_unr21_stage8_stallmux_q_4_), .o(n_32635) );
no02f80 g741935 ( .a(n_44881), .b(n_38203), .o(n_38241) );
no02f80 g766680 ( .a(n_13807), .b(n_13280), .o(n_13856) );
no02f80 g758810 ( .a(n_21789), .b(n_21788), .o(n_21807) );
ao12f80 g751071 ( .a(n_30157), .b(n_30303), .c(n_30086), .o(n_30837) );
in01f80 g736735 ( .a(n_43360), .o(n_43401) );
in01f80 g749690 ( .a(n_31482), .o(n_31483) );
no02f80 g758051 ( .a(n_22782), .b(delay_sub_ln23_0_unr16_stage6_stallmux_q_23_), .o(n_22849) );
in01f80 g749572 ( .a(n_30354), .o(n_30355) );
in01f80 FE_OCPC1469_n_23818 ( .a(n_23818), .o(FE_OCPN1469_n_23818) );
in01f80 g762024 ( .a(n_18391), .o(n_18392) );
no02f80 g764279 ( .a(n_16204), .b(n_16228), .o(n_16297) );
in01f80 g744854 ( .a(n_35167), .o(n_35168) );
in01f80 g777064 ( .a(n_4034), .o(n_3970) );
in01f80 FE_OCP_RBC2756_FE_RN_722_0 ( .a(FE_RN_722_0), .o(FE_OCP_RBN2756_FE_RN_722_0) );
ao22s80 FE_RC_4033_0 ( .a(FE_OCP_RBN3667_n_20812), .b(n_21197), .c(FE_OCP_RBN3668_n_20812), .d(n_21198), .o(n_21360) );
no02f80 g750107 ( .a(FE_OCP_RBN2572_n_29922), .b(n_29260), .o(n_30198) );
na02f80 g755232 ( .a(n_24992), .b(n_24805), .o(n_24993) );
na02f80 g751730 ( .a(n_28334), .b(n_28332), .o(n_28333) );
na02f80 g776846 ( .a(n_4005), .b(n_3885), .o(n_4126) );
ao12f80 g777745 ( .a(n_3282), .b(n_3281), .c(n_3280), .o(n_4693) );
na02f80 g740339 ( .a(n_40100), .b(n_40267), .o(n_40390) );
oa12f80 g747858 ( .a(n_33372), .b(n_32777), .c(n_33370), .o(n_33579) );
na02f80 g773582 ( .a(n_7396), .b(n_7432), .o(n_7437) );
no02f80 g744681 ( .a(n_35253), .b(n_35221), .o(n_35254) );
no02f80 g743461 ( .a(n_37680), .b(n_46244), .o(n_37681) );
na02f80 g746966 ( .a(FE_OCP_RBN2168_n_32892), .b(delay_sub_ln21_0_unr20_stage8_stallmux_q_29_), .o(n_33136) );
in01f80 g751501 ( .a(n_28912), .o(n_28913) );
in01f80 FE_RC_2430_0 ( .a(n_6887), .o(FE_RN_966_0) );
in01f80 g743769 ( .a(n_36338), .o(n_36339) );
in01f80 g737778 ( .a(n_42625), .o(n_42626) );
na02f80 g779000 ( .a(n_2161), .b(delay_add_ln22_unr2_stage2_stallmux_q_17_), .o(n_2202) );
in01f80 g746527 ( .a(n_34642), .o(n_34700) );
na02f80 g758006 ( .a(n_22200), .b(FE_OCP_RBN3221_n_22068), .o(n_22269) );
na02f80 g766484 ( .a(n_13959), .b(n_14005), .o(n_14096) );
na02f80 g780589 ( .a(n_666), .b(n_665), .o(n_677) );
no02f80 g742829 ( .a(n_37223), .b(n_36990), .o(n_37243) );
in01f80 g754733 ( .a(n_25432), .o(n_25464) );
no02f80 g746139 ( .a(n_33849), .b(n_33806), .o(n_33873) );
in01f80 FE_RC_2877_0 ( .a(n_13515), .o(FE_RN_1243_0) );
in01f80 newInst_413 ( .a(newNet_171), .o(newNet_413) );
in01f80 newInst_2108 ( .a(newNet_1989), .o(newNet_2108) );
na02f80 g762210 ( .a(n_18773), .b(n_45002), .o(n_18811) );
in01f80 FE_OCP_RBC3607_n_8981 ( .a(FE_OCP_RBN3605_n_8981), .o(FE_OCP_RBN3607_n_8981) );
na02f80 g764538 ( .a(n_16049), .b(n_16047), .o(n_16194) );
no02f80 g775139 ( .a(n_5927), .b(n_5577), .o(n_5987) );
na02f80 g744079 ( .a(n_44223), .b(n_35027), .o(n_36198) );
na02f80 g766322 ( .a(n_14533), .b(FE_OCP_RBN2510_n_13896), .o(n_14681) );
in01f80 g771187 ( .a(n_9359), .o(n_9417) );
na02f80 g738141 ( .a(n_42011), .b(n_41854), .o(n_42028) );
no02f80 g753491 ( .a(n_26874), .b(n_26873), .o(n_26913) );
no02f80 g766015 ( .a(n_14710), .b(n_14575), .o(n_14761) );
in01f80 newInst_1767 ( .a(newNet_1025), .o(newNet_1767) );
in01f80 g740005 ( .a(n_40150), .o(n_40151) );
ao12f80 g759083 ( .a(n_21452), .b(n_21909), .c(n_21410), .o(n_21959) );
na02f80 g764793 ( .a(n_15626), .b(n_15172), .o(n_15804) );
no02f80 g778233 ( .a(n_2718), .b(n_2717), .o(n_2749) );
no02f80 g758118 ( .a(n_44277), .b(n_22076), .o(n_22098) );
in01f80 FE_OCP_RBC2448_n_14114 ( .a(FE_OCP_RBN2447_n_14114), .o(FE_OCP_RBN2448_n_14114) );
in01f80 g766256 ( .a(n_14412), .o(n_14413) );
no02f80 g776868 ( .a(n_3887), .b(n_3847), .o(n_3917) );
oa12f80 g775610 ( .a(n_5518), .b(n_5552), .c(n_5517), .o(n_5578) );
in01f80 newInst_3383 ( .a(newNet_2234), .o(newNet_3383) );
in01f80 g742366 ( .a(n_37815), .o(n_37816) );
na02f80 g774813 ( .a(n_6324), .b(n_6234), .o(n_6368) );
in01f80 newInst_1297 ( .a(newNet_1062), .o(newNet_1297) );
no02f80 g737454 ( .a(n_42652), .b(n_42376), .o(n_42705) );
oa22f80 g739940 ( .a(n_40122), .b(n_40363), .c(n_40159), .d(n_40364), .o(n_40427) );
na02f80 g739572 ( .a(n_40610), .b(n_40612), .o(n_40627) );
in01f80 g764344 ( .a(n_16575), .o(n_16551) );
na02f80 g760873 ( .a(n_19467), .b(FE_OFN780_n_17093), .o(n_19468) );
in01f80 g767316 ( .a(n_13409), .o(n_13430) );
in01f80 g736611 ( .a(n_43636), .o(n_43642) );
na02f80 g767690 ( .a(n_12867), .b(n_47250), .o(n_12961) );
in01f80 g742118 ( .a(n_38233), .o(n_38234) );
na02f80 g738859 ( .a(n_41263), .b(n_41217), .o(n_41264) );
in01f80 g751360 ( .a(n_28612), .o(n_28552) );
in01f80 g771100 ( .a(n_9713), .o(n_9714) );
ao22s80 FE_RC_569_0 ( .a(n_42887), .b(n_42481), .c(n_42480), .d(n_42886), .o(n_42947) );
no02f80 g780563 ( .a(n_713), .b(n_712), .o(n_751) );
in01f80 g752194 ( .a(n_28059), .o(n_28060) );
oa22f80 FE_RC_373_0 ( .a(n_17387), .b(n_17657), .c(n_17386), .d(n_17629), .o(n_17811) );
in01f80 g757803 ( .a(n_22591), .o(n_22592) );
in01f80 g762931 ( .a(n_17792), .o(n_17793) );
in01f80 g748909 ( .a(n_32495), .o(n_32410) );
in01f80 newInst_1398 ( .a(newNet_1397), .o(newNet_1398) );
no02f80 g773056 ( .a(n_7706), .b(n_7742), .o(n_7832) );
na02f80 g777934 ( .a(n_3142), .b(n_2759), .o(n_3169) );
no02f80 g747728 ( .a(n_33668), .b(n_33701), .o(n_34106) );
in01f80 FE_OCP_RBC2961_n_26231 ( .a(FE_OCP_RBN2956_n_26231), .o(FE_OCP_RBN2961_n_26231) );
oa22f80 g775019 ( .a(n_6097), .b(n_5342), .c(n_6096), .d(n_5343), .o(n_6183) );
na02f80 g759981 ( .a(n_20675), .b(n_20657), .o(n_20676) );
na02f80 g770366 ( .a(n_10582), .b(n_44464), .o(n_10665) );
in01f80 g746194 ( .a(n_33825), .o(n_33846) );
na02f80 g766274 ( .a(n_14197), .b(n_13048), .o(n_14247) );
in01f80 FE_OCPC1503_n_47257 ( .a(n_47257), .o(FE_OCPN1503_n_47257) );
na02f80 g774279 ( .a(n_6895), .b(n_6857), .o(n_6858) );
in01f80 g750264 ( .a(n_30920), .o(n_31277) );
no02f80 g746462 ( .a(n_33344), .b(n_33343), .o(n_33345) );
in01f80 g744989 ( .a(n_34906), .o(n_34907) );
ms00f80 delay_xor_ln22_unr18_stage7_stallmux_q_reg_8_ ( .ck(newNet_429), .d(n_27779), .o(delay_xor_ln22_unr18_stage7_stallmux_q_8_) );
no02f80 FE_RC_3611_0 ( .a(n_26781), .b(FE_OCP_RBN2967_n_26580), .o(FE_RN_1579_0) );
in01f80 g740563 ( .a(n_39730), .o(n_39731) );
na02f80 g736674 ( .a(n_43232), .b(n_43199), .o(n_43369) );
in01f80 g775471 ( .a(n_5444), .o(n_5469) );
no02f80 g764436 ( .a(n_16050), .b(n_14805), .o(n_16093) );
in01f80 g772542 ( .a(FE_OCP_RBN2394_n_8288), .o(n_8334) );
in01f80 g752681 ( .a(FE_RN_1274_0), .o(n_27532) );
in01f80 g753865 ( .a(n_26304), .o(n_26305) );
na02f80 FE_RC_2324_0 ( .a(FE_RN_884_0), .b(n_28812), .o(n_28911) );
ao12f80 g737505 ( .a(n_42536), .b(n_42535), .c(n_42534), .o(n_43083) );
no02f80 g756412 ( .a(n_24040), .b(n_23970), .o(n_23971) );
na02f80 g745246 ( .a(n_36223), .b(n_36222), .o(n_36224) );
in01f80 g743574 ( .a(n_36559), .o(n_36608) );
in01f80 g747824 ( .a(n_33495), .o(n_33496) );
no02f80 g741540 ( .a(n_38715), .b(n_38716), .o(n_38726) );
in01f80 FE_OFC763_n_15670 ( .a(n_15670), .o(FE_OFN763_n_15670) );
oa12f80 g769009 ( .a(n_11993), .b(n_11689), .c(FE_OCP_RBN3268_n_45224), .o(n_11997) );
in01f80 FE_OCP_RBC2841_n_4784 ( .a(n_4784), .o(FE_OCP_RBN2841_n_4784) );
na02f80 g752935 ( .a(n_27899), .b(delay_sub_ln23_0_unr20_stage7_stallmux_q_14_), .o(n_27949) );
in01f80 g760945 ( .a(n_19453), .o(n_19497) );
in01f80 FE_OCP_RBC2810_n_15433 ( .a(n_15433), .o(FE_OCP_RBN2810_n_15433) );
no02f80 FE_RC_3961_0 ( .a(FE_RN_1715_0), .b(n_24200), .o(n_24248) );
no03m80 FE_RC_3401_0 ( .a(FE_RN_164_0), .b(n_23823), .c(n_24127), .o(n_24186) );
in01f80 g774822 ( .a(n_6414), .o(n_6391) );
na02f80 g756877 ( .a(n_23334), .b(n_23332), .o(n_23333) );
na02f80 g750818 ( .a(n_29118), .b(n_28770), .o(n_29144) );
in01f80 g758176 ( .a(n_22785), .o(n_22660) );
in01f80 FE_OCP_RBC2959_n_26231 ( .a(FE_OCP_RBN2955_n_26231), .o(FE_OCP_RBN2959_n_26231) );
no02f80 g770040 ( .a(n_10827), .b(n_9114), .o(n_10857) );
no02f80 g744055 ( .a(n_44223), .b(n_34772), .o(n_36294) );
ms00f80 delay_add_ln22_unr5_stage3_stallmux_q_reg_5_ ( .ck(newNet_2905), .d(n_4997), .o(delay_add_ln22_unr5_stage3_stallmux_q_5_) );
no02f80 g771702 ( .a(n_8791), .b(n_8784), .o(n_8880) );
oa12f80 g764761 ( .a(n_15273), .b(n_45139), .c(n_15269), .o(n_15629) );
ao12f80 g747585 ( .a(n_31947), .b(n_32324), .c(n_31898), .o(n_32382) );
in01f80 g750167 ( .a(n_29842), .o(n_29843) );
no02f80 g767376 ( .a(n_13417), .b(n_13384), .o(n_13492) );
oa12f80 g775841 ( .a(n_5263), .b(n_5262), .c(n_5261), .o(n_5371) );
in01f80 g763063 ( .a(n_17637), .o(n_17638) );
in01f80 FE_RC_2584_0 ( .a(n_17758), .o(FE_RN_1067_0) );
in01f80 g758253 ( .a(n_22649), .o(n_22728) );
in01f80 g769766 ( .a(n_11221), .o(n_11222) );
no02f80 g774082 ( .a(n_7172), .b(delay_xor_ln21_unr6_stage3_stallmux_q_21_), .o(n_7173) );
in01f80 newInst_1693 ( .a(newNet_823), .o(newNet_1693) );
in01f80 newInst_1183 ( .a(newNet_1182), .o(newNet_1183) );
na02f80 FE_RC_2905_0 ( .a(FE_RN_1257_0), .b(FE_RN_1261_0), .o(n_20167) );
na02f80 g748033 ( .a(n_44346), .b(n_32535), .o(n_33003) );
in01f80 g765728 ( .a(FE_OFN765_n_15670), .o(n_15874) );
in01f80 g752918 ( .a(n_27790), .o(n_27853) );
oa12f80 g776884 ( .a(n_3977), .b(n_3945), .c(n_3944), .o(n_4157) );
oa22f80 FE_RC_3222_0 ( .a(n_11750), .b(n_11947), .c(n_11913), .d(n_11749), .o(n_12144) );
in01f80 g764204 ( .a(n_16822), .o(n_16823) );
no02f80 g765488 ( .a(n_15874), .b(n_15957), .o(n_16173) );
ms00f80 delay_sub_ln23_0_unr24_stage9_stallmux_q_reg ( .ck(newNet_1458), .d(delay_sub_ln23_unr25_stage8_stallmux_q_3_), .o(delay_sub_ln23_0_unr24_stage9_stallmux_q) );
in01f80 g759932 ( .a(n_21482), .o(n_21402) );
in01f80 FE_OCP_RBC3377_n_1675 ( .a(n_1675), .o(FE_OCP_RBN3377_n_1675) );
in01f80 g745653 ( .a(n_34450), .o(n_34451) );
ao12f80 g742651 ( .a(n_37255), .b(n_37455), .c(n_37095), .o(n_37572) );
in01f80 FE_RC_1057_0 ( .a(FE_RN_311_0), .o(n_24269) );
na02f80 g749777 ( .a(n_31571), .b(n_31526), .o(n_31629) );
oa12f80 g761365 ( .a(n_19850), .b(n_19980), .c(n_19796), .o(n_20384) );
na02f80 g776257 ( .a(n_4536), .b(n_4665), .o(n_4804) );
no02f80 g776376 ( .a(n_4799), .b(n_4674), .o(n_4929) );
in01f80 FE_OCP_RBC3539_n_3335 ( .a(n_3335), .o(FE_OCP_RBN3539_n_3335) );
in01f80 g746598 ( .a(n_34800), .o(n_34801) );
no02f80 g755162 ( .a(n_25374), .b(n_24531), .o(n_25553) );
na02f80 g760565 ( .a(n_19858), .b(n_19696), .o(n_19920) );
in01f80 g758268 ( .a(n_22879), .o(n_22759) );
in01f80 g769921 ( .a(n_11026), .o(n_11085) );
na02f80 g741961 ( .a(n_38053), .b(n_38118), .o(n_38119) );
no02f80 g768329 ( .a(n_12514), .b(n_12513), .o(n_12515) );
in01f80 newInst_1989 ( .a(newNet_1988), .o(newNet_1989) );
ao12f80 g773542 ( .a(n_7483), .b(n_45864), .c(n_7481), .o(n_7877) );
na02f80 g765848 ( .a(n_14804), .b(n_14442), .o(n_14886) );
na02f80 g739115 ( .a(n_41014), .b(n_40887), .o(n_41015) );
in01f80 FE_OCP_RBC3359_delay_sub_ln23_unr13_stage5_stallmux_q_1_ ( .a(FE_OCP_RBN3296_delay_sub_ln23_unr13_stage5_stallmux_q_1_), .o(FE_OCP_RBN3359_delay_sub_ln23_unr13_stage5_stallmux_q_1_) );
ao12f80 g771025 ( .a(n_9556), .b(n_9761), .c(n_9635), .o(n_9926) );
no02f80 g740957 ( .a(n_39252), .b(n_38928), .o(n_39213) );
in01f80 FE_OCP_RBC3111_n_43871 ( .a(n_43871), .o(FE_OCP_RBN3111_n_43871) );
na02f80 g751876 ( .a(n_28946), .b(n_28907), .o(n_28908) );
in01f80 FE_OCP_RBC3835_n_19241 ( .a(FE_OCP_RBN3834_n_19241), .o(FE_OCP_RBN3835_n_19241) );
ao12f80 g754592 ( .a(n_26637), .b(n_26856), .c(n_26604), .o(n_26888) );
na02f80 g769610 ( .a(n_11375), .b(n_11419), .o(n_11426) );
in01f80 newInst_1603 ( .a(newNet_1602), .o(newNet_1603) );
no02f80 g778028 ( .a(n_3018), .b(n_2741), .o(n_3049) );
no02f80 g780844 ( .a(n_478), .b(n_445), .o(n_630) );
na03f80 FE_RC_1491_0 ( .a(n_22816), .b(n_22820), .c(n_22708), .o(n_22990) );
na02f80 g746701 ( .a(n_34276), .b(n_33813), .o(n_34277) );
no02f80 g755879 ( .a(n_25191), .b(n_25285), .o(n_25192) );
in01f80 newInst_2693 ( .a(newNet_2692), .o(newNet_2693) );
no02f80 g750048 ( .a(n_29869), .b(n_29898), .o(n_29928) );
in01f80 g753731 ( .a(n_26502), .o(n_26503) );
na02f80 g758071 ( .a(n_22507), .b(FE_OCP_RBN1709_n_22150), .o(n_22508) );
in01f80 g751683 ( .a(n_28458), .o(n_28597) );
na02f80 g760677 ( .a(n_19690), .b(FE_OCP_RBN1700_n_19353), .o(n_19746) );
in01f80 g764026 ( .a(n_18032), .o(n_18099) );
no02f80 g761813 ( .a(n_18322), .b(n_18193), .o(n_18348) );
in01f80 g760540 ( .a(n_19946), .o(n_19967) );
in01f80 g752699 ( .a(n_27313), .o(n_27314) );
in01f80 g771038 ( .a(n_9625), .o(n_9668) );
ao12f80 g743524 ( .a(n_36841), .b(n_37584), .c(n_36852), .o(n_37680) );
in01f80 g761569 ( .a(n_20231), .o(n_22580) );
no02f80 g763480 ( .a(n_15656), .b(n_16814), .o(n_16839) );
na02f80 g762109 ( .a(n_18884), .b(n_18810), .o(n_18885) );
in01f80 g736883 ( .a(n_43597), .o(n_43598) );
na02f80 g754825 ( .a(n_25303), .b(FE_OCPN985_n_25210), .o(n_25361) );
no02f80 FE_RC_3673_0 ( .a(FE_RN_1613_0), .b(n_31379), .o(n_31439) );
ao12f80 g738259 ( .a(n_41874), .b(n_41873), .c(n_41872), .o(n_41921) );
no02f80 g765934 ( .a(n_14812), .b(n_14788), .o(n_14871) );
in01f80 g737295 ( .a(n_42941), .o(n_42926) );
no02f80 g778944 ( .a(n_2257), .b(n_1971), .o(n_2268) );
no02f80 FE_RC_858_0 ( .a(FE_RN_257_0), .b(n_43152), .o(n_43153) );
na02f80 g765218 ( .a(n_16023), .b(n_15968), .o(n_16062) );
in01f80 g747312 ( .a(n_34474), .o(n_33929) );
in01f80 g761919 ( .a(n_18319), .o(n_18320) );
in01f80 g748112 ( .a(n_31746), .o(n_31688) );
in01f80 g754426 ( .a(n_25731), .o(n_25730) );
na02f80 g757219 ( .a(n_23527), .b(n_23526), .o(n_23528) );
na02f80 g759314 ( .a(n_46968), .b(n_21212), .o(n_21342) );
in01f80 g776810 ( .a(n_4015), .o(n_4016) );
no02f80 g784408 ( .a(n_46204), .b(delay_sub_ln23_0_unr28_stage9_stallmux_q_13_), .o(n_46220) );
in01f80 g773576 ( .a(n_7384), .o(n_7385) );
ao12f80 g746388 ( .a(n_33220), .b(n_33501), .c(n_33152), .o(n_33561) );
no02f80 g750512 ( .a(n_29505), .b(FE_OCPN1432_n_29504), .o(n_29525) );
na02f80 g756016 ( .a(n_25160), .b(n_25250), .o(n_25741) );
no02f80 g740198 ( .a(n_40210), .b(n_40247), .o(n_40248) );
in01f80 g751268 ( .a(n_29767), .o(n_29768) );
no02f80 g740658 ( .a(n_39525), .b(n_39528), .o(n_39557) );
no02f80 g766333 ( .a(n_14164), .b(n_13323), .o(n_14279) );
no02f80 g739323 ( .a(n_45149), .b(delay_add_ln22_unr27_stage10_stallmux_q_27_), .o(n_40859) );
in01f80 g756633 ( .a(n_24275), .o(n_24257) );
in01f80 g761283 ( .a(n_19037), .o(n_19038) );
no02f80 g737006 ( .a(n_43230), .b(n_42993), .o(n_43387) );
in01f80 FE_OCP_DRV_C1590_n_21343 ( .a(FE_OCP_DRV_N1589_n_21343), .o(FE_OCP_DRV_N1590_n_21343) );
in01f80 g740419 ( .a(n_40097), .o(n_40051) );
na02f80 FE_RC_599_0 ( .a(FE_RN_186_0), .b(FE_RN_187_0), .o(FE_RN_188_0) );
ms00f80 delay_add_ln22_unr27_stage10_stallmux_q_reg_0_ ( .ck(newNet_3178), .d(n_39708), .o(delay_add_ln22_unr27_stage10_stallmux_q_0_) );
na02f80 g742088 ( .a(FE_OCP_RBN3451_n_37945), .b(n_37597), .o(n_38216) );
na02f80 g741811 ( .a(n_38484), .b(n_39232), .o(n_38485) );
in01f80 g746044 ( .a(n_35259), .o(n_35804) );
in01f80 FE_OCP_RBC3708_n_31396 ( .a(n_31396), .o(FE_OCP_RBN3708_n_31396) );
ao12f80 g782652 ( .a(n_27923), .b(n_27931), .c(n_27854), .o(n_44046) );
oa12f80 g749467 ( .a(n_30170), .b(n_30471), .c(n_30470), .o(n_30501) );
no02f80 g738946 ( .a(n_41159), .b(n_40962), .o(n_41249) );
na02f80 g739552 ( .a(n_44027), .b(n_40660), .o(n_40685) );
no02f80 g780921 ( .a(n_357), .b(n_362), .o(n_369) );
ao12f80 g772268 ( .a(n_8113), .b(n_8684), .c(n_8048), .o(n_8824) );
no02f80 g773560 ( .a(n_7402), .b(n_7401), .o(n_7411) );
na02f80 g745960 ( .a(n_35299), .b(n_35279), .o(n_35280) );
no02f80 g764292 ( .a(n_16330), .b(n_14588), .o(n_16332) );
in01f80 FE_OCPC916_n_46991 ( .a(n_46991), .o(FE_OCPN916_n_46991) );
ao22s80 g736549 ( .a(n_43569), .b(n_43178), .c(n_43570), .d(n_43177), .o(n_43652) );
no02f80 g769811 ( .a(n_11192), .b(n_44498), .o(n_11193) );
in01f80 g742065 ( .a(n_38033), .o(n_38084) );
in01f80 g736877 ( .a(n_43603), .o(n_43604) );
no02f80 g758068 ( .a(n_22729), .b(n_22644), .o(n_22761) );
in01f80 newInst_2141 ( .a(newNet_2140), .o(newNet_2141) );
na02f80 g753282 ( .a(n_27377), .b(n_26276), .o(n_27461) );
na02f80 g766798 ( .a(n_13748), .b(n_13747), .o(n_13749) );
in01f80 newInst_1027 ( .a(newNet_1026), .o(newNet_1027) );
in01f80 g752943 ( .a(n_27763), .o(n_27764) );
na02f80 g737760 ( .a(n_42307), .b(n_42417), .o(n_42353) );
oa12f80 g780111 ( .a(n_1013), .b(n_1029), .c(n_1012), .o(n_1082) );
ao12f80 g768846 ( .a(n_11821), .b(n_11699), .c(n_11440), .o(n_11822) );
no02f80 g765221 ( .a(n_15785), .b(n_15750), .o(n_15838) );
in01f80 FE_OCPUNCOC1805_n_19801 ( .a(n_19801), .o(FE_OCPUNCON1805_n_19801) );
in01f80 FE_OCP_RBC2001_delay_sub_ln23_unr9_stage4_stallmux_q_3_ ( .a(delay_sub_ln23_unr9_stage4_stallmux_q_3_), .o(FE_OCP_RBN2001_delay_sub_ln23_unr9_stage4_stallmux_q_3_) );
in01f80 newInst_2573 ( .a(newNet_2572), .o(newNet_2573) );
na02f80 g779292 ( .a(n_1659), .b(delay_add_ln22_unr2_stage2_stallmux_q_5_), .o(n_1745) );
na02f80 g765638 ( .a(n_15006), .b(n_14919), .o(n_15074) );
no02f80 g737230 ( .a(n_42919), .b(n_42931), .o(n_43251) );
na02f80 g766559 ( .a(n_13921), .b(n_13471), .o(n_14023) );
no02f80 g776655 ( .a(n_47009), .b(FE_OCP_RBN2465_n_4336), .o(n_4394) );
oa22f80 g763213 ( .a(n_46973), .b(n_17336), .c(n_17187), .d(n_17753), .o(n_17337) );
in01f80 FE_OCP_RBC2485_n_38601 ( .a(n_38601), .o(FE_OCP_RBN2485_n_38601) );
na02f80 g751572 ( .a(n_28437), .b(delay_sub_ln21_0_unr17_stage7_stallmux_q_14_), .o(n_28547) );
in01f80 g777386 ( .a(n_3643), .o(n_3711) );
oa12f80 g744022 ( .a(n_46203), .b(n_36860), .c(delay_sub_ln23_unr29_stage9_stallmux_q_2_), .o(n_37631) );
ao22s80 g754195 ( .a(n_26016), .b(n_25662), .c(n_25956), .d(n_25661), .o(n_26081) );
in01f80 g760046 ( .a(n_20439), .o(n_20440) );
in01f80 g777981 ( .a(n_47022), .o(n_3144) );
ao12f80 g742758 ( .a(n_37221), .b(n_37291), .c(n_36969), .o(n_37326) );
no02f80 g738500 ( .a(FE_OCPN952_n_41540), .b(n_41415), .o(n_41786) );
na02f80 g780521 ( .a(n_698), .b(n_685), .o(n_765) );
in01f80 g747566 ( .a(delay_add_ln22_unr20_stage8_stallmux_q_22_), .o(n_32303) );
in01f80 g748181 ( .a(n_32124), .o(n_32125) );
na02f80 g748716 ( .a(n_31165), .b(n_31164), .o(n_31271) );
no02f80 g755037 ( .a(n_25233), .b(n_25208), .o(n_25514) );
no02f80 g778539 ( .a(n_2278), .b(n_2031), .o(n_2323) );
in01f80 g760269 ( .a(n_20428), .o(n_20456) );
na02f80 FE_RC_2856_0 ( .a(FE_RN_1230_0), .b(n_13857), .o(n_13884) );
na02f80 g745308 ( .a(n_36119), .b(n_36118), .o(n_36120) );
na02f80 g776112 ( .a(n_5024), .b(n_4442), .o(n_5078) );
ao12f80 g746115 ( .a(n_35128), .b(n_35127), .c(n_35126), .o(n_35765) );
in01f80 newInst_2965 ( .a(newNet_2367), .o(newNet_2965) );
in01f80 g771745 ( .a(n_8919), .o(n_8920) );
in01f80 g745455 ( .a(n_34459), .o(n_34487) );
na02f80 g770444 ( .a(n_10577), .b(n_10576), .o(n_10578) );
na02f80 g773975 ( .a(n_7217), .b(delay_xor_ln21_unr6_stage3_stallmux_q_24_), .o(n_7239) );
in01f80 g744820 ( .a(n_36494), .o(n_36495) );
na02f80 g745216 ( .a(n_36226), .b(n_36225), .o(n_36227) );
in01f80 FE_RC_1635_0 ( .a(n_11908), .o(FE_RN_454_0) );
na02f80 g754572 ( .a(FE_OCP_RBN2959_n_26231), .b(n_26734), .o(n_26832) );
no02f80 g736950 ( .a(FE_OCPN912_n_43022), .b(n_42941), .o(n_43280) );
no02f80 FE_RC_3661_0 ( .a(n_21552), .b(FE_RN_1607_0), .o(n_21769) );
no02f80 g741294 ( .a(n_44944), .b(n_38472), .o(n_38939) );
in01f80 FE_OFC776_n_17093 ( .a(n_17093), .o(FE_OFN776_n_17093) );
na02f80 g751270 ( .a(n_28790), .b(n_28777), .o(n_28778) );
in01f80 g745856 ( .a(n_35406), .o(n_35407) );
in01f80 g751479 ( .a(n_28703), .o(n_28704) );
oa12f80 g775464 ( .a(n_5382), .b(n_5486), .c(n_5440), .o(n_5487) );
in01f80 newInst_3380 ( .a(newNet_3379), .o(newNet_3380) );
in01f80 g772731 ( .a(n_8263), .o(n_8264) );
oa22f80 g748619 ( .a(n_31485), .b(n_31490), .c(n_31484), .d(n_29966), .o(n_31646) );
no02f80 g744802 ( .a(n_35130), .b(n_30633), .o(n_35170) );
na02f80 g736795 ( .a(n_43518), .b(n_43385), .o(n_43554) );
no02f80 FE_RC_3933_0 ( .a(n_11918), .b(FE_RN_1701_0), .o(n_11770) );
no02f80 g743723 ( .a(n_37342), .b(n_37434), .o(n_37382) );
no02f80 g751338 ( .a(n_28806), .b(n_28744), .o(n_28851) );
na02f80 g762335 ( .a(n_18383), .b(n_18382), .o(n_18384) );
na02f80 g751443 ( .a(n_28742), .b(n_28741), .o(n_28743) );
in01f80 g778250 ( .a(n_2792), .o(n_2756) );
na02f80 g737895 ( .a(n_42201), .b(n_42139), .o(n_42383) );
ao12f80 g775846 ( .a(n_4578), .b(n_4776), .c(n_4659), .o(n_4907) );
na02f80 g776860 ( .a(n_4175), .b(n_4066), .o(n_4226) );
in01f80 newInst_2946 ( .a(newNet_2781), .o(newNet_2946) );
ao12f80 g761214 ( .a(n_18945), .b(n_19025), .c(FE_OFN779_n_17093), .o(n_19104) );
in01f80 g738827 ( .a(n_41372), .o(n_41366) );
oa22f80 FE_RC_1607_0 ( .a(FE_OCP_RBN1349_n_19270), .b(n_20429), .c(FE_OCPN999_n_19311), .d(n_20428), .o(n_20578) );
na02f80 g776597 ( .a(n_4484), .b(n_4395), .o(n_4563) );
in01f80 g743275 ( .a(delay_sub_ln21_unr24_stage9_stallmux_q_1_), .o(n_36844) );
no02f80 g775818 ( .a(n_5359), .b(n_5143), .o(n_5435) );
in01f80 FE_OCPC3166_n_44267 ( .a(FE_OCPN3165_n_44267), .o(FE_OCPN3166_n_44267) );
na02f80 g744081 ( .a(n_44223), .b(n_34996), .o(n_36143) );
in01f80 g766369 ( .a(n_14160), .o(n_14161) );
in01f80 g780054 ( .a(n_1238), .o(n_1239) );
in01f80 g747658 ( .a(delay_sub_ln21_0_unr20_stage8_stallmux_q_17_), .o(n_32362) );
in01f80 g757341 ( .a(n_23131), .o(n_23104) );
na02f80 g741718 ( .a(n_38506), .b(n_38156), .o(n_38523) );
ao12f80 g757614 ( .a(n_22676), .b(n_22675), .c(delay_add_ln22_unr14_stage6_stallmux_q_0_), .o(n_24119) );

endmodule
