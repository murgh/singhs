module top;

// Start PIs
input pmem_d_14;
input io_di_7;
input dmem_di_0;
input dmem_di_2;
input pmem_d_0;
input tau_clk;
input pmem_d_10;
input io_di_2;
input io_di_3;
input pmem_d_2;
input pmem_d_11;
input dmem_di_7;
input dmem_di_6;
input pmem_d_15;
input io_di_5;
input io_di_1;
input rst;
input pmem_d_13;
input pmem_d_9;
input io_di_4;
input pmem_d_8;
input io_di_0;
input dmem_di_5;
input pmem_d_3;
input dmem_di_4;
input pmem_d_4;
input pmem_d_5;
input pmem_d_6;
input dmem_di_3;
input dmem_di_1;
input io_di_6;
input pmem_d_12;
input pmem_d_1;
input pmem_d_7;

// Start POs
output dmem_do_3;
output dmem_a_4;
output io_do_1;
output dmem_a_9;
output pmem_a_9;
output dmem_a_10;
output io_we;
output dmem_a_6;
output pmem_ce;
output io_do_3;
output dmem_do_0;
output io_do_6;
output pmem_a_0;
output pmem_a_10;
output dmem_a_11;
output dmem_do_6;
output dmem_a_5;
output pmem_a_7;
output pmem_a_8;
output io_do_5;
output dmem_a_3;
output dmem_a_0;
output io_do_4;
output dmem_do_4;
output pmem_a_4;
output pmem_a_3;
output io_a_0;
output dmem_do_1;
output io_re;
output dmem_a_7;
output dmem_a_12;
output dmem_ce;
output dmem_do_2;
output pmem_a_1;
output dmem_do_5;
output io_do_2;
output io_do_7;
output io_a_1;
output io_do_0;
output io_a_4;
output pmem_a_2;
output pmem_a_5;
output dmem_we;
output io_a_3;
output dmem_a_8;
output dmem_do_7;
output dmem_a_2;
output io_a_5;
output io_a_2;
output pmem_a_6;
output dmem_a_1;

// Start wires
wire n_1514;
wire n_356;
wire newNet_1460;
wire n_707;
wire n_2478;
wire newNet_1761;
wire n_4132;
wire newNet_166;
wire n_997;
wire io_sel_0_;
wire n_685;
wire n_192;
wire n_1822;
wire n_2907;
wire newNet_451;
wire newNet_73;
wire n_1266;
wire n_3389;
wire n_1363;
wire GPR_10__2_;
wire newNet_828;
wire newNet_342;
wire n_1759;
wire n_61;
wire n_4316;
wire n_4185;
wire n_502;
wire n_3332;
wire n_4608;
wire newNet_1849;
wire n_2048;
wire n_98;
wire n_4115;
wire n_3775;
wire state_0_;
wire n_4165;
wire newNet_1302;
wire GPR_22__7_;
wire newNet_1689;
wire n_2794;
wire n_89;
wire n_2030;
wire newNet_862;
wire n_868;
wire n_4095;
wire n_3171;
wire n_2992;
wire final_adder_mux_R16_278_6_n_37;
wire n_3935;
wire n_1313;
wire n_1452;
wire n_2839;
wire n_861;
wire GPR_10__3_;
wire n_114;
wire newNet_857;
wire newNet_562;
wire n_1047;
wire n_1519;
wire n_3289;
wire n_3450;
wire n_1062;
wire newNet_1685;
wire newNet_1213;
wire newNet_1178;
wire n_682;
wire newNet_546;
wire n_2226;
wire n_2719;
wire n_2889;
wire n_4660;
wire n_3959;
wire newNet_1303;
wire n_68;
wire n_3044;
wire n_4147;
wire GPR_14__2_;
wire newNet_662;
wire newNet_1162;
wire n_2979;
wire n_4652;
wire n_2234;
wire n_2155;
wire pZ_0_;
wire newNet_674;
wire R16_6_;
wire n_811;
wire n_4262;
wire n_629;
wire newNet_1641;
wire n_3181;
wire n_4427;
wire n_1347;
wire n_3167;
wire newNet_183;
wire n_1731;
wire n_2116;
wire newNet_1648;
wire newNet_1339;
wire n_4648;
wire n_3534;
wire n_2217;
wire n_2821;
wire n_4570;
wire n_1279;
wire n_3257;
wire n_1948;
wire n_4042;
wire n_2158;
wire newNet_1202;
wire newNet_346;
wire n_1856;
wire n_937;
wire n_2138;
wire newNet_1237;
wire n_2287;
wire newNet_627;
wire newNet_319;
wire newNet_1855;
wire n_2582;
wire n_2810;
wire newNet_689;
wire n_1271;
wire n_4407;
wire final_adder_mux_R16_278_6_n_81;
wire n_3845;
wire n_2148;
wire n_2980;
wire n_3340;
wire n_4394;
wire n_2547;
wire n_2999;
wire newNet_1773;
wire n_958;
wire n_3015;
wire n_4312;
wire n_2423;
wire n_3398;
wire n_1233;
wire newNet_927;
wire n_324;
wire n_1674;
wire newNet_1446;
wire n_1585;
wire final_adder_mux_R16_278_6_n_44;
wire n_486;
wire n_2628;
wire Rd_2_;
wire newNet_1615;
wire newNet_1350;
wire n_800;
wire n_1355;
wire n_1650;
wire PC_0_;
wire newNet_1467;
wire n_1175;
wire n_1160;
wire n_1944;
wire n_1039;
wire n_3806;
wire pY_7_;
wire n_4267;
wire n_3472;
wire n_2970;
wire newNet_1023;
wire newNet_5;
wire newNet_1430;
wire n_4180;
wire newNet_521;
wire n_1045;
wire newNet_1711;
wire n_2925;
wire n_485;
wire n_2338;
wire newNet_1622;
wire n_4150;
wire n_3730;
wire n_4097;
wire n_884;
wire n_222;
wire n_796;
wire dmem_di_1;
wire newNet_1651;
wire n_3074;
wire n_2777;
wire n_506;
wire n_3552;
wire pmem_d_7;
wire newNet_695;
wire n_1485;
wire n_2601;
wire newNet_848;
wire n_4110;
wire newNet_390;
wire n_2598;
wire n_3527;
wire newNet_1487;
wire n_2083;
wire newNet_721;
wire newNet_335;
wire n_1605;
wire n_606;
wire n_920;
wire n_2766;
wire n_2700;
wire n_158;
wire n_4257;
wire newNet_967;
wire newNet_138;
wire n_1053;
wire newNet_1704;
wire newNet_293;
wire n_894;
wire newNet_1782;
wire GPR_17__0_;
wire newNet_936;
wire newNet_867;
wire n_3766;
wire n_1500;
wire n_624;
wire n_2092;
wire n_2899;
wire n_1659;
wire newNet_882;
wire n_1005;
wire n_1013;
wire n_3467;
wire n_4228;
wire n_727;
wire n_3500;
wire newNet_1565;
wire newNet_607;
wire newNet_504;
wire n_298;
wire n_4386;
wire newNet_285;
wire newNet_177;
wire n_2293;
wire n_4027;
wire newNet_1102;
wire n_3198;
wire newNet_1273;
wire n_2789;
wire n_1320;
wire n_3799;
wire n_3917;
wire newNet_648;
wire newNet_509;
wire n_2065;
wire newNet_705;
wire newNet_811;
wire n_200;
wire n_2671;
wire newNet_1241;
wire n_2487;
wire n_2847;
wire n_1988;
wire n_3116;
wire newNet_1732;
wire n_3164;
wire n_3790;
wire newNet_1275;
wire n_4033;
wire n_2571;
wire newNet_1004;
wire n_35;
wire n_513;
wire n_2884;
wire n_3950;
wire n_2672;
wire dmem_a_0;
wire n_1871;
wire io_do_4;
wire n_2663;
wire newNet_479;
wire n_817;
wire n_2175;
wire n_2;
wire n_954;
wire n_20;
wire n_2141;
wire n_431;
wire newNet_1400;
wire n_477;
wire n_4002;
wire newNet_779;
wire newNet_669;
wire n_2041;
wire newNet_388;
wire n_1069;
wire n_175;
wire n_531;
wire newNet_485;
wire newNet_878;
wire n_4051;
wire newNet_983;
wire newNet_424;
wire n_692;
wire n_3143;
wire n_1643;
wire n_3236;
wire n_2084;
wire n_2947;
wire newNet_1585;
wire n_2453;
wire n_597;
wire n_1666;
wire n_4364;
wire newNet_1175;
wire newNet_1144;
wire n_4060;
wire newNet_1458;
wire n_2723;
wire newNet_588;
wire n_1285;
wire n_2935;
wire n_2912;
wire n_124;
wire n_1627;
wire n_2455;
wire n_95;
wire n_4036;
wire n_3437;
wire n_552;
wire pY_3_;
wire n_3815;
wire n_1923;
wire n_2833;
wire GPR_2__6_;
wire n_3365;
wire n_3861;
wire n_4210;
wire n_1924;
wire newNet_591;
wire GPR_16__3_;
wire newNet_748;
wire n_651;
wire n_4175;
wire newNet_1598;
wire newNet_1482;
wire n_9;
wire n_590;
wire n_3396;
wire n_3788;
wire newNet_941;
wire newNet_899;
wire n_1093;
wire n_2697;
wire n_2415;
wire n_3787;
wire n_2127;
wire n_2375;
wire n_1124;
wire newNet_152;
wire n_4432;
wire n_1566;
wire n_1423;
wire newNet_482;
wire newNet_1315;
wire n_3674;
wire newNet_836;
wire n_522;
wire n_3212;
wire n_2386;
wire n_787;
wire n_3359;
wire n_3026;
wire n_255;
wire n_2350;
wire newNet_1243;
wire newNet_35;
wire n_1422;
wire n_2100;
wire newNet_304;
wire n_1794;
wire newNet_1577;
wire n_2842;
wire newNet_1715;
wire n_1415;
wire n_4561;
wire Rd_0_;
wire n_2357;
wire pZ_4_;
wire newNet_834;
wire newNet_1068;
wire n_3567;
wire n_4083;
wire newNet_240;
wire newNet_1842;
wire n_848;
wire newNet_396;
wire io_sp_5_;
wire n_3362;
wire newNet_1658;
wire newNet_444;
wire n_78;
wire n_2023;
wire newNet_1209;
wire R16_8_;
wire n_3458;
wire newNet_1423;
wire newNet_1042;
wire newNet_412;
wire n_2054;
wire n_2615;
wire n_1190;
wire R16_7_;
wire n_3885;
wire n_3391;
wire newNet_1528;
wire newNet_870;
wire n_4489;
wire n_4221;
wire io_a_2;
wire newNet_1494;
wire n_2167;
wire n_3086;
wire n_499;
wire n_1183;
wire n_2321;
wire n_2816;
wire n_245;
wire n_1249;
wire n_3126;
wire n_3067;
wire n_4276;
wire newNet_96;
wire newNet_1387;
wire newNet_307;
wire n_422;
wire n_4313;
wire newNet_806;
wire n_1621;
wire newNet_1802;
wire n_1741;
wire newNet_407;
wire n_3947;
wire n_4643;
wire newNet_1037;
wire n_3335;
wire n_713;
wire n_2851;
wire newNet_1265;
wire n_2955;
wire n_967;
wire n_3640;
wire newNet_1811;
wire newNet_356;
wire n_833;
wire newNet_87;
wire n_666;
wire dmem_a_7;
wire n_496;
wire n_133;
wire newNet_1294;
wire n_3710;
wire n_3298;
wire n_907;
wire n_2525;
wire newNet_259;
wire n_1469;
wire newNet_68;
wire n_2540;
wire n_3296;
wire n_2653;
wire n_131;
wire n_1546;
wire n_3506;
wire n_4323;
wire newNet_1502;
wire n_2318;
wire n_2166;
wire newNet_437;
wire n_3485;
wire newNet_752;
wire n_814;
wire n_1074;
wire n_1906;
wire n_994;
wire newNet_526;
wire newNet_243;
wire GPR_19__2_;
wire io_di_2;
wire newNet_1634;
wire n_574;
wire n_729;
wire GPR_13__1_;
wire newNet_571;
wire n_3378;
wire n_3419;
wire n_3052;
wire n_3979;
wire n_1526;
wire newNet_281;
wire newNet_443;
wire newNet_1348;
wire newNet_145;
wire n_2189;
wire n_292;
wire n_1158;
wire n_1784;
wire n_2878;
wire n_1004;
wire n_3441;
wire n_3906;
wire newNet_1065;
wire n_471;
wire n_754;
wire n_2378;
wire n_1094;
wire n_1901;
wire newNet_765;
wire n_474;
wire newNet_952;
wire n_3873;
wire n_1295;
wire n_3936;
wire n_1488;
wire n_376;
wire n_1966;
wire n_1692;
wire n_2767;
wire n_1881;
wire newNet_276;
wire newNet_95;
wire n_455;
wire n_2906;
wire n_3324;
wire n_841;
wire newNet_784;
wire newNet_766;
wire newNet_1559;
wire n_2323;
wire n_3076;
wire n_3457;
wire GPR_21__1_;
wire newNet_805;
wire newNet_1805;
wire newNet_1762;
wire newNet_1251;
wire n_2264;
wire n_3603;
wire newNet_1545;
wire n_2803;
wire n_4317;
wire n_193;
wire newNet_1610;
wire n_4370;
wire n_2572;
wire n_2390;
wire PC_4_;
wire n_201;
wire n_143;
wire n_3117;
wire n_4123;
wire n_2071;
wire n_377;
wire newNet_195;
wire n_3623;
wire n_3948;
wire newNet_1744;
wire n_1076;
wire n_3325;
wire GPR_11__7_;
wire n_2108;
wire n_3739;
wire n_3027;
wire newNet_1195;
wire newNet_712;
wire n_71;
wire n_2649;
wire n_2864;
wire newNet_1473;
wire final_adder_mux_R16_278_6_n_11;
wire newNet_249;
wire GPR_15__6_;
wire n_4306;
wire n_1847;
wire R16_10_;
wire n_2259;
wire newNet_171;
wire n_2633;
wire newNet_1378;
wire newNet_672;
wire n_3982;
wire newNet_360;
wire n_4411;
wire newNet_1754;
wire newNet_1016;
wire n_2669;
wire n_2624;
wire n_41;
wire n_3560;
wire n_1713;
wire newNet_476;
wire newNet_1679;
wire n_2640;
wire GPR_9__7_;
wire newNet_462;
wire n_100;
wire n_1853;
wire Rd_1_;
wire n_2014;
wire n_655;
wire n_1840;
wire n_2035;
wire n_1725;
wire n_4231;
wire n_3246;
wire newNet_735;
wire newNet_251;
wire n_1891;
wire n_1677;
wire n_2305;
wire n_4341;
wire n_542;
wire newNet_890;
wire n_4467;
wire n_3727;
wire newNet_1323;
wire n_2556;
wire GPR_16__6_;
wire final_adder_mux_R16_278_6_n_72;
wire n_1805;
wire n_1774;
wire newNet_1385;
wire n_1991;
wire n_1756;
wire newNet_1649;
wire n_783;
wire n_1943;
wire n_2883;
wire newNet_15;
wire GPR_9__3_;
wire n_1184;
wire newNet_34;
wire newNet_530;
wire GPR_3__6_;
wire newNet_687;
wire n_117;
wire n_2534;
wire n_1426;
wire GPR_12__1_;
wire n_3962;
wire newNet_887;
wire newNet_772;
wire n_988;
wire n_2347;
wire final_adder_mux_R16_278_6_n_84;
wire n_4061;
wire GPR_3__5_;
wire n_3426;
wire newNet_1835;
wire n_4474;
wire n_3961;
wire newNet_907;
wire n_2432;
wire n_3176;
wire newNet_1017;
wire n_1135;
wire n_1567;
wire n_3860;
wire n_4208;
wire newNet_1338;
wire n_984;
wire n_834;
wire n_1436;
wire n_2746;
wire newNet_590;
wire newNet_381;
wire n_615;
wire n_1612;
wire n_48;
wire n_3988;
wire n_3341;
wire n_3366;
wire n_1020;
wire newNet_1794;
wire newNet_1586;
wire n_2919;
wire newNet_40;
wire newNet_1642;
wire n_3205;
wire n_367;
wire n_1080;
wire n_440;
wire n_1492;
wire n_774;
wire n_2987;
wire GPR_0__5_;
wire dmem_a_10;
wire n_481;
wire n_726;
wire n_979;
wire n_226;
wire n_1258;
wire n_563;
wire newNet_1139;
wire n_1752;
wire newNet_103;
wire final_adder_mux_R16_278_6_n_63;
wire newNet_161;
wire n_2211;
wire GPR_15__0_;
wire GPR_13__3_;
wire newNet_1630;
wire n_3135;
wire n_3301;
wire GPR_21__0_;
wire pmem_d_15;
wire newNet_1414;
wire n_449;
wire n_3499;
wire newNet_926;
wire n_1715;
wire newNet_1450;
wire pY_8_;
wire n_3520;
wire n_2368;
wire newNet_1445;
wire n_3972;
wire newNet_1130;
wire n_3273;
wire n_4426;
wire n_4217;
wire newNet_159;
wire n_1685;
wire n_3697;
wire n_1709;
wire n_1917;
wire n_2734;
wire newNet_1090;
wire n_770;
wire n_2004;
wire N;
wire newNet_387;
wire newNet_217;
wire newNet_696;
wire n_673;
wire n_1114;
wire n_1579;
wire newNet_947;
wire n_213;
wire n_4518;
wire n_2966;
wire n_1532;
wire newNet_875;
wire n_1813;
wire n_288;
wire n_3159;
wire n_398;
wire n_4157;
wire newNet_203;
wire n_1206;
wire n_1161;
wire n_1501;
wire n_1103;
wire newNet_1522;
wire newNet_333;
wire n_29;
wire newNet_1731;
wire newNet_1309;
wire n_3442;
wire newNet_127;
wire n_706;
wire n_2505;
wire n_344;
wire n_4236;
wire newNet_1552;
wire n_2486;
wire newNet_1101;
wire n_10;
wire newNet_971;
wire n_432;
wire n_1204;
wire final_adder_mux_R16_278_6_n_16;
wire n_3581;
wire newNet_682;
wire n_2497;
wire n_4536;
wire newNet_1678;
wire SP_13_;
wire n_2049;
wire n_876;
wire n_239;
wire pmem_ce;
wire n_1118;
wire n_3826;
wire n_3000;
wire n_3655;
wire n_309;
wire newNet_1764;
wire n_337;
wire n_4609;
wire n_3981;
wire newNet_931;
wire n_3188;
wire n_3253;
wire n_14;
wire n_1381;
wire n_314;
wire n_4204;
wire newNet_45;
wire n_3895;
wire n_3648;
wire newNet_1535;
wire newNet_633;
wire newNet_1797;
wire n_3745;
wire n_2203;
wire pmem_a_5;
wire n_4107;
wire n_761;
wire n_4243;
wire n_4190;
wire n_3613;
wire n_1148;
wire io_do_1;
wire n_4263;
wire newNet_1187;
wire n_3109;
wire n_307;
wire n_2272;
wire newNet_58;
wire n_1593;
wire n_3241;
wire newNet_1616;
wire newNet_1147;
wire n_8;
wire newNet_1035;
wire n_911;
wire newNet_1291;
wire n_3927;
wire newNet_1208;
wire newNet_920;
wire n_3689;
wire dmem_do_4;
wire n_746;
wire newNet_1283;
wire n_380;
wire newNet_1163;
wire n_442;
wire n_1911;
wire newNet_1600;
wire n_900;
wire n_4011;
wire newNet_1088;
wire n_929;
wire newNet_231;
wire newNet_347;
wire n_4074;
wire n_3221;
wire n_3631;
wire n_3834;
wire n_3358;
wire newNet_608;
wire n_1730;
wire GPR_8__4_;
wire n_4448;
wire n_3387;
wire n_2705;
wire n_3776;
wire n_1651;
wire n_1983;
wire final_adder_mux_R16_278_6_n_23;
wire n_2132;
wire n_4237;
wire n_1682;
wire n_1416;
wire n_4440;
wire n_3812;
wire n_2294;
wire n_959;
wire n_3158;
wire n_1372;
wire n_297;
wire n_520;
wire GPR_5__7_;
wire n_3999;
wire n_3411;
wire n_184;
wire n_3602;
wire n_3884;
wire pY_10_;
wire newNet_25;
wire newNet_1863;
wire newNet_578;
wire n_1234;
wire n_2831;
wire n_2546;
wire newNet_1456;
wire n_2440;
wire n_4353;
wire n_3844;
wire n_484;
wire newNet_940;
wire n_3204;
wire n_1691;
wire n_2732;
wire n_854;
wire n_2924;
wire n_157;
wire n_877;
wire newNet_1783;
wire newNet_494;
wire n_1658;
wire n_125;
wire n_1302;
wire n_2239;
wire n_323;
wire n_2753;
wire n_4005;
wire GPR_5__0_;
wire n_1629;
wire newNet_336;
wire newNet_160;
wire n_1354;
wire n_1449;
wire newNet_1829;
wire n_3614;
wire n_724;
wire n_2592;
wire n_2597;
wire n_2778;
wire n_3263;
wire n_3399;
wire n_1619;
wire n_883;
wire newNet_1413;
wire n_1046;
wire PC_8_;
wire n_4151;
wire dmem_di_2;
wire newNet_1284;
wire newNet_1466;
wire n_4094;
wire newNet_1799;
wire newNet_297;
wire n_227;
wire final_adder_mux_R16_278_6_n_38;
wire newNet_1659;
wire newNet_845;
wire n_507;
wire n_1855;
wire n_2701;
wire n_2815;
wire n_223;
wire GPR_13__4_;
wire n_3079;
wire n_2149;
wire n_1012;
wire newNet_286;
wire newNet_139;
wire newNet_1591;
wire n_4385;
wire newNet_1186;
wire n_3274;
wire n_4291;
wire newNet_1363;
wire n_4655;
wire GPR_20__2_;
wire n_4096;
wire n_2664;
wire newNet_881;
wire n_4391;
wire n_2488;
wire n_909;
wire newNet_868;
wire n_2279;
wire n_1054;
wire n_1675;
wire newNet_722;
wire newNet_309;
wire newNet_1426;
wire n_1278;
wire newNet_226;
wire n_1349;
wire n_4014;
wire n_1482;
wire n_4084;
wire newNet_984;
wire n_1513;
wire n_2091;
wire n_97;
wire newNet_1810;
wire newNet_343;
wire n_3262;
wire newNet_771;
wire newNet_1274;
wire n_3791;
wire U_13_;
wire n_3774;
wire n_3165;
wire n_1048;
wire n_115;
wire n_70;
wire newNet_188;
wire n_2956;
wire n_246;
wire n_3924;
wire newNet_777;
wire n_835;
wire newNet_357;
wire n_4131;
wire n_3088;
wire n_2174;
wire newNet_1803;
wire n_1312;
wire newNet_1301;
wire io_do_2;
wire GPR_5__2_;
wire newNet_1686;
wire n_675;
wire n_1930;
wire n_693;
wire n_4634;
wire newNet_423;
wire n_4032;
wire n_3958;
wire n_503;
wire n_1031;
wire final_adder_mux_R16_278_6_n_29;
wire n_1841;
wire n_1970;
wire n_867;
wire n_1267;
wire n_195;
wire n_3805;
wire n_500;
wire newNet_1159;
wire n_2397;
wire newNet_320;
wire n_3482;
wire n_77;
wire n_3132;
wire n_3466;
wire n_739;
wire n_4146;
wire n_2587;
wire n_2117;
wire n_944;
wire n_2187;
wire n_287;
wire n_2139;
wire n_4043;
wire n_1136;
wire n_2859;
wire newNet_321;
wire newNet_112;
wire newNet_169;
wire n_3709;
wire n_3883;
wire n_683;
wire n_4158;
wire n_3290;
wire n_3453;
wire n_2978;
wire n_2233;
wire n_1949;
wire n_1100;
wire n_406;
wire n_2159;
wire newNet_539;
wire n_4311;
wire n_565;
wire n_2462;
wire n_4619;
wire newNet_619;
wire n_69;
wire n_1584;
wire n_3151;
wire n_2834;
wire n_3687;
wire n_4186;
wire n_2694;
wire n_2948;
wire newNet_450;
wire n_825;
wire n_3193;
wire n_461;
wire newNet_274;
wire n_2316;
wire GPR_14__6_;
wire newNet_241;
wire n_3459;
wire newNet_1067;
wire n_3677;
wire n_4573;
wire n_3808;
wire newNet_1316;
wire n_2648;
wire newNet_1231;
wire newNet_65;
wire n_4325;
wire n_3666;
wire n_4562;
wire newNet_819;
wire newNet_36;
wire n_3780;
wire newNet_143;
wire n_4396;
wire n_4166;
wire n_3091;
wire n_3336;
wire newNet_1821;
wire GPR_12__0_;
wire n_2262;
wire newNet_915;
wire n_543;
wire n_2024;
wire newNet_1324;
wire n_1502;
wire n_2053;
wire n_2790;
wire n_2625;
wire n_3007;
wire GPR_0__2_;
wire n_3855;
wire newNet_89;
wire n_3045;
wire n_1326;
wire n_3397;
wire n_3087;
wire n_4230;
wire newNet_835;
wire io_a_3;
wire final_adder_mux_R16_278_6_n_80;
wire n_1620;
wire n_2768;
wire n_607;
wire n_2307;
wire newNet_466;
wire newNet_258;
wire n_2322;
wire n_4380;
wire n_1147;
wire newNet_833;
wire n_2739;
wire n_1527;
wire n_4277;
wire dmem_a_6;
wire newNet_408;
wire n_1964;
wire newNet_1114;
wire n_1545;
wire newNet_563;
wire n_3066;
wire n_2449;
wire newNet_1675;
wire n_4218;
wire newNet_1629;
wire newNet_303;
wire n_1407;
wire newNet_93;
wire n_712;
wire n_1560;
wire newNet_636;
wire newNet_296;
wire GPR_19__1_;
wire n_1182;
wire n_2908;
wire newNet_82;
wire n_132;
wire U_6_;
wire n_4405;
wire newNet_1843;
wire final_adder_mux_R16_278_6_n_13;
wire newNet_1214;
wire newNet_1041;
wire n_4598;
wire newNet_1395;
wire n_130;
wire n_4604;
wire newNet_308;
wire newNet_176;
wire n_2408;
wire n_3297;
wire newNet_1266;
wire n_4039;
wire n_413;
wire newNet_1184;
wire n_690;
wire n_2606;
wire n_1997;
wire n_3142;
wire n_3211;
wire newNet_704;
wire n_4490;
wire GPR_4__4_;
wire newNet_812;
wire n_1897;
wire newNet_1760;
wire newNet_508;
wire newNet_668;
wire n_934;
wire n_3295;
wire n_4406;
wire newNet_949;
wire n_2911;
wire n_3110;
wire n_921;
wire n_2477;
wire n_4227;
wire n_1922;
wire newNet_531;
wire n_795;
wire newNet_1201;
wire n_818;
wire n_3258;
wire n_176;
wire n_1980;
wire n_3465;
wire newNet_1018;
wire n_2852;
wire n_1626;
wire n_1461;
wire n_3537;
wire n_1;
wire newNet_1003;
wire n_955;
wire n_3702;
wire n_3061;
wire newNet_778;
wire n_4526;
wire n_4625;
wire newNet_1608;
wire n_4425;
wire n_2848;
wire n_1783;
wire n_4642;
wire newNet_478;
wire n_2670;
wire newNet_389;
wire GPR_Rd_r_0_;
wire newNet_1647;
wire n_497;
wire n_530;
wire newNet_1809;
wire newNet_1129;
wire newNet_1179;
wire n_21;
wire n_1179;
wire n_3012;
wire n_3652;
wire newNet_1652;
wire newNet_1440;
wire n_1576;
wire pmem_d_14;
wire newNet_1176;
wire n_4220;
wire newNet_718;
wire newNet_417;
wire newNet_1420;
wire n_1335;
wire n_1789;
wire state_1_;
wire n_657;
wire n_2635;
wire n_4176;
wire n_4211;
wire newNet_612;
wire n_2392;
wire n_849;
wire newNet_337;
wire n_1284;
wire n_820;
wire n_2881;
wire newNet_1455;
wire n_1724;
wire n_3331;
wire n_1776;
wire n_2936;
wire newNet_1665;
wire n_2711;
wire n_2456;
wire n_1872;
wire n_3875;
wire newNet_998;
wire newNet_851;
wire newNet_1481;
wire newNet_713;
wire GPR_15__4_;
wire n_3738;
wire n_598;
wire n_430;
wire n_1989;
wire n_551;
wire n_2629;
wire R16_3_;
wire newNet_802;
wire n_2454;
wire n_3069;
wire n_3553;
wire newNet_690;
wire GPR_5__3_;
wire newNet_151;
wire n_1555;
wire n_533;
wire n_3960;
wire n_40;
wire n_4244;
wire n_1099;
wire newNet_1580;
wire n_4624;
wire n_2251;
wire n_3721;
wire newNet_170;
wire newNet_1566;
wire n_3369;
wire n_2249;
wire n_4553;
wire n_2013;
wire newNet_671;
wire n_3222;
wire newNet_1379;
wire newNet_1771;
wire newNet_80;
wire n_985;
wire n_1848;
wire newNet_16;
wire n_2431;
wire n_782;
wire n_3427;
wire newNet_957;
wire n_3528;
wire n_3319;
wire pmem_a_4;
wire n_2795;
wire n_650;
wire n_4359;
wire n_1425;
wire n_2043;
wire newNet_1364;
wire newNet_264;
wire n_3969;
wire final_adder_mux_R16_278_6_n_9;
wire n_3432;
wire n_2086;
wire n_3254;
wire n_4347;
wire n_2555;
wire n_1531;
wire n_4410;
wire n_336;
wire n_3097;
wire n_1336;
wire n_0;
wire n_3042;
wire n_4250;
wire final_adder_mux_R16_278_6_n_22;
wire newNet_1836;
wire n_2745;
wire n_4342;
wire n_3821;
wire newNet_1484;
wire newNet_230;
wire n_7;
wire n_912;
wire n_2306;
wire n_1435;
wire newNet_57;
wire n_2042;
wire n_4209;
wire n_1633;
wire newNet_76;
wire n_971;
wire n_1712;
wire n_1091;
wire n_3983;
wire newNet_1666;
wire final_adder_mux_R16_278_6_n_56;
wire GPR_22__3_;
wire GPR_14__1_;
wire GPR_16__7_;
wire newNet_418;
wire n_82;
wire n_3758;
wire newNet_1570;
wire n_368;
wire n_3312;
wire n_4314;
wire n_1178;
wire n_1990;
wire n_3445;
wire n_771;
wire n_3744;
wire newNet_253;
wire n_989;
wire pY_14_;
wire pX_15_;
wire newNet_1755;
wire newNet_1000;
wire n_475;
wire newNet_1819;
wire n_3989;
wire n_423;
wire n_480;
wire n_2425;
wire n_1613;
wire n_1395;
wire n_2526;
wire newNet_688;
wire newNet_999;
wire newNet_252;
wire n_387;
wire n_2231;
wire n_3342;
wire newNet_751;
wire n_2263;
wire n_3753;
wire n_2214;
wire n_2712;
wire n_2812;
wire newNet_1745;
wire newNet_852;
wire n_2416;
wire n_2652;
wire n_3068;
wire n_3418;
wire newNet_1806;
wire newNet_1070;
wire newNet_1156;
wire n_755;
wire n_2413;
wire n_2185;
wire GPR_9__1_;
wire newNet_282;
wire n_4040;
wire newNet_609;
wire newNet_144;
wire n_443;
wire n_2188;
wire n_3130;
wire n_3019;
wire n_4324;
wire n_4563;
wire newNet_1822;
wire n_1479;
wire SP_14_;
wire n_3127;
wire newNet_1633;
wire n_1900;
wire io_a_0;
wire pZ_12_;
wire n_2990;
wire io_di_1;
wire n_1157;
wire n_1714;
wire newNet_1349;
wire n_1967;
wire n_1146;
wire n_2399;
wire n_3440;
wire n_3053;
wire n_3153;
wire PC_10_;
wire newNet_1080;
wire n_1487;
wire n_4274;
wire n_1606;
wire n_3120;
wire n_4363;
wire newNet_1525;
wire n_291;
wire n_4205;
wire n_275;
wire n_1371;
wire n_194;
wire newNet_953;
wire n_4525;
wire newNet_586;
wire n_842;
wire n_1294;
wire n_301;
wire n_870;
wire newNet_785;
wire newNet_767;
wire n_278;
wire newNet_126;
wire n_3420;
wire newNet_898;
wire newNet_1854;
wire dmem_a_11;
wire newNet_275;
wire newNet_1252;
wire n_2308;
wire newNet_1143;
wire n_4124;
wire n_375;
wire n_3566;
wire n_4645;
wire newNet_600;
wire newNet_1516;
wire n_2377;
wire newNet_1721;
wire n_2345;
wire n_108;
wire n_2407;
wire n_1075;
wire n_142;
wire n_2383;
wire n_3326;
wire n_399;
wire n_806;
wire newNet_557;
wire newNet_1774;
wire newNet_1503;
wire n_1073;
wire n_786;
wire GPR_3__0_;
wire n_1884;
wire final_adder_mux_R16_278_6_n_10;
wire n_1198;
wire n_4667;
wire n_3874;
wire n_2352;
wire n_3949;
wire n_1892;
wire n_2072;
wire n_523;
wire n_3572;
wire n_2531;
wire newNet_620;
wire n_2204;
wire n_1742;
wire n_1250;
wire newNet_358;
wire n_2424;
wire n_2580;
wire newNet_1796;
wire final_adder_mux_R16_278_6_n_19;
wire n_1007;
wire n_2632;
wire n_2872;
wire SP_10_;
wire n_1571;
wire n_4318;
wire n_36;
wire n_3856;
wire newNet_640;
wire n_3001;
wire newNet_747;
wire n_2280;
wire n_260;
wire n_456;
wire n_1348;
wire pmem_d_8;
wire n_4535;
wire n_2324;
wire n_4010;
wire newNet_1164;
wire n_760;
wire n_1638;
wire newNet_736;
wire n_4138;
wire n_1119;
wire n_3937;
wire n_1115;
wire n_1380;
wire newNet_541;
wire GPR_10__1_;
wire n_308;
wire n_265;
wire n_2877;
wire n_3663;
wire n_1971;
wire n_2219;
wire n_3386;
wire n_1753;
wire n_2003;
wire n_2918;
wire n_2317;
wire n_4189;
wire n_901;
wire n_4449;
wire newNet_1099;
wire n_13;
wire newNet_382;
wire n_4419;
wire n_3177;
wire n_1775;
wire n_2133;
wire GPR_2__0_;
wire n_1618;
wire n_3686;
wire newNet_1062;
wire n_747;
wire n_2165;
wire V;
wire n_635;
wire n_928;
wire n_1865;
wire n_47;
wire newNet_794;
wire n_3634;
wire n_2704;
wire n_2809;
wire n_3388;
wire pX_0_;
wire dmem_do_7;
wire n_1460;
wire n_3434;
wire GPR_12__2_;
wire n_2496;
wire newNet_1200;
wire newNet_111;
wire newNet_114;
wire newNet_104;
wire n_669;
wire n_2733;
wire n_1916;
wire n_4431;
wire n_4273;
wire newNet_647;
wire newNet_1553;
wire n_672;
wire GPR_4__5_;
wire newNet_179;
wire GPR_11__0_;
wire n_3104;
wire n_1683;
wire n_2271;
wire n_4339;
wire n_4618;
wire n_2802;
wire n_3998;
wire n_215;
wire n_4597;
wire newNet_1739;
wire n_860;
wire n_564;
wire n_1259;
wire n_441;
wire n_4372;
wire GPR_1__1_;
wire n_740;
wire n_2359;
wire newNet_209;
wire n_738;
wire n_1223;
wire n_3370;
wire n_3515;
wire n_3973;
wire newNet_1341;
wire newNet_131;
wire n_2824;
wire newNet_1234;
wire n_978;
wire newNet_1705;
wire n_2195;
wire final_adder_mux_R16_278_6_n_65;
wire n_2038;
wire n_24;
wire n_212;
wire newNet_37;
wire n_582;
wire n_961;
wire n_3498;
wire n_654;
wire n_156;
wire n_964;
wire n_614;
wire n_3375;
wire newNet_438;
wire Rd_r_3_;
wire n_2989;
wire n_4378;
wire n_2724;
wire newNet_1131;
wire n_3696;
wire n_2367;
wire n_101;
wire n_1640;
wire n_2348;
wire n_343;
wire newNet_1299;
wire newNet_1699;
wire n_54;
wire newNet_972;
wire newNet_395;
wire n_2997;
wire newNet_1308;
wire n_2612;
wire n_3185;
wire n_4015;
wire n_1806;
wire n_3591;
wire newNet_1225;
wire n_3381;
wire n_4075;
wire newNet_372;
wire n_3350;
wire newNet_1059;
wire n_3649;
wire GPR_1__7_;
wire n_3405;
wire newNet_1239;
wire n_1126;
wire newNet_1546;
wire n_1442;
wire newNet_1100;
wire n_3647;
wire n_313;
wire n_2863;
wire n_3521;
wire newNet_723;
wire n_390;
wire n_3894;
wire n_4571;
wire n_3145;
wire GPR_5__4_;
wire n_1770;
wire newNet_568;
wire n_775;
wire newNet_1730;
wire n_1814;
wire n_628;
wire n_1215;
wire n_4392;
wire newNet_946;
wire n_3582;
wire n_1757;
wire n_3189;
wire n_2278;
wire n_2258;
wire newNet_929;
wire n_3703;
wire newNet_298;
wire newNet_1670;
wire newNet_218;
wire n_1169;
wire n_2674;
wire n_4430;
wire newNet_1382;
wire n_2940;
wire newNet_1039;
wire n_1534;
wire GPR_6__4_;
wire n_1095;
wire n_2485;
wire n_3020;
wire n_1340;
wire n_1894;
wire n_2339;
wire newNet_930;
wire newNet_483;
wire n_232;
wire newNet_536;
wire n_2665;
wire n_694;
wire n_4102;
wire n_1602;
wire n_592;
wire n_1561;
wire n_2509;
wire n_611;
wire n_3464;
wire n_4557;
wire n_1641;
wire newNet_973;
wire n_4079;
wire n_1141;
wire newNet_38;
wire newNet_804;
wire n_4020;
wire n_2169;
wire n_3128;
wire newNet_1002;
wire n_3514;
wire n_815;
wire n_3684;
wire newNet_1511;
wire n_3089;
wire newNet_985;
wire newNet_1496;
wire n_1296;
wire newNet_1804;
wire newNet_1653;
wire n_4491;
wire n_1931;
wire n_2457;
wire n_3118;
wire newNet_876;
wire n_1578;
wire newNet_189;
wire n_550;
wire GPR_19__6_;
wire n_247;
wire n_1766;
wire n_2461;
wire n_599;
wire n_318;
wire n_2754;
wire newNet_1168;
wire n_1921;
wire newNet_799;
wire n_1771;
wire newNet_26;
wire n_1467;
wire n_2626;
wire n_2562;
wire n_1764;
wire n_426;
wire n_808;
wire n_2695;
wire n_2879;
wire n_404;
wire n_3100;
wire newNet_1858;
wire n_1101;
wire n_2569;
wire newNet_1161;
wire n_3238;
wire newNet_1177;
wire n_2849;
wire n_4038;
wire n_1173;
wire U_7_;
wire n_3488;
wire n_557;
wire n_4035;
wire n_947;
wire n_3162;
wire n_1008;
wire n_1390;
wire newNet_1409;
wire n_2370;
wire n_262;
wire n_2843;
wire n_1493;
wire n_3824;
wire n_4641;
wire newNet_1109;
wire final_adder_mux_R16_278_6_n_14;
wire newNet_1480;
wire newNet_220;
wire n_2588;
wire newNet_269;
wire n_159;
wire final_adder_mux_R16_278_6_n_53;
wire SP_12_;
wire n_3785;
wire n_3393;
wire n_3352;
wire n_4589;
wire newNet_1848;
wire newNet_119;
wire n_826;
wire n_1283;
wire newNet_801;
wire newNet_3;
wire n_3813;
wire n_3769;
wire n_2314;
wire GPR_4__0_;
wire n_1350;
wire n_3673;
wire n_3065;
wire newNet_1766;
wire n_126;
wire n_183;
wire newNet_257;
wire n_566;
wire n_2021;
wire n_3048;
wire n_1325;
wire n_1122;
wire n_1437;
wire n_4616;
wire n_3615;
wire n_4167;
wire n_1628;
wire n_2160;
wire n_1301;
wire n_3569;
wire n_3601;
wire newNet_47;
wire newNet_1357;
wire n_1548;
wire newNet_1044;
wire newNet_832;
wire n_1831;
wire n_1181;
wire n_2245;
wire n_4366;
wire n_2074;
wire n_715;
wire newNet_1207;
wire n_3653;
wire n_3364;
wire n_424;
wire newNet_1296;
wire newNet_1260;
wire n_1067;
wire newNet_1851;
wire newNet_964;
wire GPR_15__3_;
wire newNet_0;
wire n_1528;
wire n_1886;
wire n_2059;
wire n_2142;
wire n_4602;
wire n_1904;
wire GPR_10__5_;
wire dmem_a_5;
wire newNet_1676;
wire newNet_714;
wire n_4568;
wire n_2814;
wire n_2105;
wire n_2642;
wire n_4264;
wire newNet_503;
wire pY_2_;
wire n_1541;
wire n_2617;
wire newNet_776;
wire n_2355;
wire newNet_939;
wire n_1417;
wire GPR_14__3_;
wire newNet_1425;
wire n_2177;
wire n_459;
wire n_794;
wire io_a_4;
wire newNet_1578;
wire newNet_446;
wire n_3796;
wire newNet_762;
wire n_135;
wire n_3187;
wire n_2953;
wire newNet_1189;
wire n_1402;
wire n_1406;
wire pX_2_;
wire GPR_7__5_;
wire newNet_467;
wire newNet_1077;
wire n_4605;
wire n_3712;
wire n_680;
wire n_935;
wire GPR_21__6_;
wire n_1824;
wire n_4252;
wire n_4153;
wire n_3892;
wire n_812;
wire n_1458;
wire n_1950;
wire n_1016;
wire n_3121;
wire n_1883;
wire n_161;
wire newNet_1369;
wire n_315;
wire n_720;
wire n_4636;
wire n_3150;
wire newNet_1687;
wire newNet_900;
wire n_3259;
wire n_3887;
wire newNet_1123;
wire n_4013;
wire n_2787;
wire newNet_864;
wire n_3940;
wire n_3732;
wire n_2994;
wire n_896;
wire newNet_770;
wire n_1361;
wire newNet_1211;
wire n_878;
wire n_3706;
wire GPR_8__2_;
wire newNet_453;
wire newNet_1464;
wire n_2094;
wire n_514;
wire n_3210;
wire newNet_1393;
wire n_4295;
wire GPR_22__5_;
wire n_3111;
wire n_3804;
wire n_1516;
wire n_2124;
wire n_560;
wire n_886;
wire n_1176;
wire n_4484;
wire n_1448;
wire newNet_1683;
wire n_2439;
wire newNet_733;
wire n_3256;
wire pY_1_;
wire newNet_1788;
wire newNet_75;
wire n_2421;
wire n_3483;
wire pY_5_;
wire newNet_1717;
wire n_1338;
wire n_3957;
wire n_2002;
wire newNet_1432;
wire newNet_344;
wire n_2968;
wire R16_12_;
wire n_4388;
wire newNet_897;
wire n_412;
wire n_3719;
wire newNet_1557;
wire newNet_1713;
wire n_4099;
wire n_1273;
wire newNet_495;
wire n_518;
wire n_2398;
wire n_4415;
wire newNet_1664;
wire n_2238;
wire n_3438;
wire n_3008;
wire n_2717;
wire n_1826;
wire newNet_556;
wire n_4626;
wire U_0_;
wire newNet_1337;
wire n_490;
wire n_995;
wire n_2289;
wire n_2184;
wire n_759;
wire pX_7_;
wire newNet_1524;
wire newNet_859;
wire n_1384;
wire n_1946;
wire n_4113;
wire n_2114;
wire n_1264;
wire n_1583;
wire n_871;
wire n_4305;
wire newNet_1442;
wire GPR_21__3_;
wire n_3549;
wire pZ_14_;
wire newNet_429;
wire n_1040;
wire n_2949;
wire newNet_1599;
wire newNet_869;
wire n_354;
wire newNet_667;
wire n_1218;
wire newNet_1437;
wire n_1038;
wire Rd_r_4_;
wire newNet_527;
wire newNet_1775;
wire n_286;
wire n_3898;
wire n_1199;
wire pY_12_;
wire n_220;
wire n_3646;
wire GPR_20__4_;
wire GPR_10__0_;
wire n_407;
wire n_2257;
wire n_250;
wire n_2927;
wire n_329;
wire newNet_1780;
wire newNet_614;
wire newNet_287;
wire n_3658;
wire newNet_854;
wire newNet_128;
wire n_116;
wire n_2972;
wire newNet_322;
wire n_322;
wire n_3410;
wire final_adder_mux_R16_278_6_n_57;
wire n_2729;
wire n_2827;
wire n_4356;
wire n_2157;
wire n_1329;
wire n_3203;
wire newNet_1448;
wire newNet_1370;
wire n_2982;
wire dmem_di_3;
wire newNet_1119;
wire newNet_410;
wire n_1652;
wire newNet_180;
wire n_575;
wire n_856;
wire newNet_1411;
wire n_16064_BAR;
wire n_2905;
wire newNet_295;
wire n_388;
wire n_1669;
wire n_3219;
wire newNet_1465;
wire n_2775;
wire n_1854;
wire n_4424;
wire n_1687;
wire n_4285;
wire n_1319;
wire n_2028;
wire n_2209;
wire n_2295;
wire newNet_1792;
wire n_396;
wire n_2591;
wire n_4159;
wire newNet_1824;
wire n_4290;
wire n_559;
wire n_2448;
wire n_709;
wire n_1235;
wire n_3078;
wire n_4058;
wire n_2897;
wire io_sp_6_;
wire n_4588;
wire pZ_8_;
wire n_3284;
wire newNet_227;
wire n_864;
wire n_2228;
wire newNet_1623;
wire n_1049;
wire io_re;
wire n_1357;
wire n_1483;
wire newNet_909;
wire n_744;
wire newNet_1763;
wire n_2118;
wire n_4599;
wire newNet_468;
wire n_224;
wire newNet_1259;
wire n_3541;
wire newNet_1300;
wire n_1676;
wire U_9_;
wire n_4658;
wire n_2518;
wire n_4152;
wire n_3264;
wire n_638;
wire n_4665;
wire n_3974;
wire n_1499;
wire n_2080;
wire n_2213;
wire newNet_1438;
wire n_2067;
wire n_345;
wire newNet_694;
wire pmem_d_0;
wire newNet_178;
wire n_969;
wire n_2799;
wire newNet_1813;
wire newNet_585;
wire n_1216;
wire n_3037;
wire n_102;
wire n_1572;
wire n_1863;
wire n_4515;
wire newNet_1098;
wire newNet_840;
wire n_4018;
wire n_1732;
wire n_3836;
wire n_3303;
wire n_444;
wire n_668;
wire n_3524;
wire n_357;
wire n_2406;
wire n_613;
wire n_2511;
wire n_2417;
wire n_1116;
wire n_2342;
wire newNet_488;
wire n_733;
wire newNet_1718;
wire n_1086;
wire newNet_601;
wire newNet_518;
wire n_1377;
wire n_268;
wire n_3497;
wire final_adder_mux_R16_278_6_n_46;
wire newNet_1220;
wire newNet_924;
wire n_3638;
wire n_3237;
wire n_776;
wire newNet_657;
wire n_237;
wire n_214;
wire n_439;
wire n_1671;
wire n_2332;
wire newNet_454;
wire Rd_4_;
wire newNet_1720;
wire pZ_9_;
wire n_2201;
wire n_1610;
wire n_3919;
wire n_2503;
wire n_3587;
wire newNet_1673;
wire newNet_1233;
wire n_3147;
wire newNet_200;
wire n_3556;
wire n_2973;
wire newNet_1142;
wire newNet_813;
wire n_3695;
wire dmem_do_6;
wire n_4269;
wire newNet_1560;
wire n_316;
wire newNet_404;
wire H;
wire n_589;
wire n_850;
wire n_4234;
wire newNet_1475;
wire n_93;
wire GPR_7__6_;
wire newNet_554;
wire n_1815;
wire GPR_6__0_;
wire newNet_263;
wire n_785;
wire n_1956;
wire dmem_do_1;
wire newNet_378;
wire n_4279;
wire newNet_1639;
wire n_2019;
wire newNet_1030;
wire n_3218;
wire newNet_13;
wire n_805;
wire n_3850;
wire n_3571;
wire n_119;
wire n_1318;
wire n_4377;
wire newNet_11;
wire n_3955;
wire n_2728;
wire n_4371;
wire n_88;
wire n_2483;
wire n_1208;
wire n_2969;
wire n_2130;
wire n_2242;
wire newNet_793;
wire newNet_1452;
wire newNet_219;
wire n_335;
wire n_3255;
wire n_2060;
wire n_2655;
wire n_3997;
wire newNet_1082;
wire R16_4_;
wire n_1383;
wire n_3245;
wire n_4081;
wire n_1639;
wire n_2903;
wire newNet_615;
wire n_4265;
wire n_4538;
wire n_3223;
wire newNet_1118;
wire n_2274;
wire newNet_685;
wire newNet_1706;
wire n_1503;
wire newNet_373;
wire n_1936;
wire n_3192;
wire n_4192;
wire n_2329;
wire n_1112;
wire n_3385;
wire newNet_954;
wire newNet_724;
wire newNet_349;
wire n_3920;
wire n_55;
wire newNet_1293;
wire n_2220;
wire n_2178;
wire n_3718;
wire n_4121;
wire n_2871;
wire n_3402;
wire final_adder_mux_R16_278_6_n_66;
wire n_2805;
wire newNet_210;
wire newNet_1307;
wire n_2874;
wire n_3003;
wire newNet_1285;
wire n_970;
wire newNet_90;
wire n_3910;
wire n_2495;
wire n_2479;
wire n_1734;
wire newNet_1253;
wire n_2952;
wire newNet_567;
wire n_3275;
wire newNet_1860;
wire n_3107;
wire n_1225;
wire n_4130;
wire newNet_641;
wire newNet_540;
wire newNet_146;
wire tau_clk;
wire n_2282;
wire GPR_7__7_;
wire n_634;
wire newNet_1132;
wire n_2792;
wire newNet_1697;
wire n_4387;
wire n_3662;
wire newNet_27;
wire n_2703;
wire n_1985;
wire n_2232;
wire newNet_933;
wire n_913;
wire n_3002;
wire newNet_415;
wire n_3548;
wire n_2607;
wire newNet_105;
wire n_973;
wire n_580;
wire n_927;
wire n_2266;
wire n_4072;
wire n_767;
wire n_1750;
wire n_3848;
wire n_3598;
wire n_3995;
wire n_4331;
wire n_4054;
wire newNet_1618;
wire newNet_1571;
wire GPR_7__1_;
wire n_3763;
wire n_544;
wire n_3752;
wire newNet_750;
wire n_1072;
wire n_4631;
wire newNet_1550;
wire newNet_524;
wire n_3343;
wire newNet_1588;
wire newNet_129;
wire newNet_579;
wire n_546;
wire n_2751;
wire n_962;
wire pX_14_;
wire final_adder_mux_R16_278_6_n_59;
wire n_2539;
wire n_1945;
wire n_2685;
wire n_905;
wire n_1060;
wire newNet_1807;
wire n_1418;
wire n_1807;
wire newNet_1124;
wire final_adder_mux_R16_278_6_n_28;
wire n_1022;
wire n_1476;
wire newNet_919;
wire n_3904;
wire n_3546;
wire n_203;
wire n_90;
wire newNet_351;
wire n_2403;
wire n_992;
wire newNet_1504;
wire GPR_15__7_;
wire n_3368;
wire n_4315;
wire newNet_1485;
wire newNet_9;
wire newNet_283;
wire n_781;
wire n_3351;
wire n_294;
wire n_3327;
wire n_671;
wire n_2991;
wire newNet_394;
wire n_2885;
wire n_4067;
wire n_1559;
wire newNet_782;
wire n_2052;
wire n_1972;
wire n_3669;
wire n_3570;
wire n_524;
wire n_458;
wire newNet_1738;
wire final_adder_mux_R16_278_6_n_0;
wire newNet_1342;
wire n_3152;
wire newNet_816;
wire newNet_1325;
wire n_196;
wire n_508;
wire n_3452;
wire n_3621;
wire n_2813;
wire n_3968;
wire n_3986;
wire newNet_741;
wire n_1690;
wire n_379;
wire n_678;
wire newNet_1632;
wire newNet_246;
wire newNet_132;
wire n_1006;
wire n_276;
wire n_1486;
wire n_4233;
wire n_816;
wire n_3095;
wire n_2360;
wire n_4145;
wire n_2769;
wire newNet_1729;
wire newNet_1746;
wire n_752;
wire n_1362;
wire n_1893;
wire n_1474;
wire n_4610;
wire n_1151;
wire newNet_528;
wire n_2504;
wire GPR_22__2_;
wire n_2384;
wire n_2044;
wire n_1580;
wire newNet_1567;
wire n_2545;
wire n_4439;
wire n_3797;
wire GPR_18__6_;
wire n_3505;
wire n_3314;
wire n_1866;
wire newNet_950;
wire n_4304;
wire n_1256;
wire newNet_1009;
wire n_4259;
wire n_1845;
wire n_3725;
wire newNet_430;
wire newNet_1643;
wire n_4441;
wire n_164;
wire n_81;
wire newNet_965;
wire newNet_97;
wire n_4465;
wire pmem_d_9;
wire newNet_650;
wire n_1648;
wire n_248;
wire n_626;
wire newNet_173;
wire n_302;
wire n_1441;
wire n_4206;
wire n_3694;
wire newNet_759;
wire n_4409;
wire n_3428;
wire n_1297;
wire n_1767;
wire n_3133;
wire newNet_1336;
wire n_4344;
wire n_4382;
wire n_1678;
wire newNet_383;
wire n_3859;
wire n_3720;
wire n_3862;
wire n_2073;
wire n_144;
wire n_1388;
wire newNet_831;
wire newNet_1113;
wire newNet_889;
wire n_2773;
wire n_1603;
wire n_1438;
wire n_3768;
wire n_4545;
wire newNet_1051;
wire n_365;
wire n_1466;
wire newNet_1061;
wire n_2303;
wire newNet_1310;
wire n_150;
wire n_836;
wire n_695;
wire n_1912;
wire n_4088;
wire newNet_1383;
wire newNet_84;
wire n_1699;
wire n_2381;
wire n_2532;
wire n_2748;
wire GPR_15__1_;
wire n_4556;
wire n_2760;
wire GPR_21__4_;
wire newNet_278;
wire n_986;
wire n_4202;
wire n_576;
wire n_1368;
wire n_1838;
wire n_2225;
wire newNet_1592;
wire newNet_703;
wire n_1133;
wire newNet_1693;
wire n_1397;
wire n_3163;
wire n_2012;
wire n_1717;
wire final_adder_mux_R16_278_6_n_45;
wire n_46;
wire n_3672;
wire GPR_12__4_;
wire newNet_110;
wire newNet_1092;
wire newNet_1069;
wire n_2143;
wire n_960;
wire final_adder_mux_R16_278_6_n_17;
wire n_4408;
wire n_2194;
wire n_745;
wire newNet_1765;
wire n_1282;
wire n_4122;
wire n_3353;
wire n_3786;
wire newNet_1457;
wire n_4222;
wire newNet_1181;
wire newNet_1663;
wire newNet_2;
wire newNet_247;
wire n_823;
wire newNet_1356;
wire n_4266;
wire n_3049;
wire n_509;
wire newNet_1579;
wire n_1440;
wire n_2327;
wire n_3123;
wire n_3616;
wire n_1272;
wire n_3664;
wire newNet_1712;
wire n_4168;
wire n_3064;
wire n_2022;
wire n_3031;
wire n_1330;
wire n_4438;
wire n_3555;
wire n_4365;
wire n_1106;
wire n_2051;
wire io_do_7;
wire GPR_21__2_;
wire n_3568;
wire n_3578;
wire newNet_1850;
wire n_830;
wire n_3864;
wire SP_15_;
wire newNet_715;
wire n_498;
wire U_11_;
wire newNet_1841;
wire state_2_;
wire newNet_1043;
wire newNet_800;
wire newNet_529;
wire n_2244;
wire U_15_;
wire n_2447;
wire dmem_a_4;
wire newNet_634;
wire n_4003;
wire newNet_1488;
wire n_3299;
wire n_1540;
wire io_we;
wire n_2337;
wire n_4483;
wire newNet_938;
wire newNet_1823;
wire newNet_359;
wire n_1604;
wire newNet_502;
wire n_1504;
wire newNet_46;
wire n_3129;
wire n_1180;
wire n_2176;
wire n_1547;
wire n_3390;
wire n_1021;
wire n_1401;
wire n_1885;
wire n_3094;
wire n_3632;
wire n_205;
wire n_3608;
wire n_3535;
wire n_4374;
wire n_1529;
wire newNet_1727;
wire newNet_763;
wire n_231;
wire newNet_277;
wire n_1823;
wire n_2330;
wire newNet_702;
wire newNet_492;
wire PC_2_;
wire newNet_951;
wire n_4229;
wire GPR_15__2_;
wire n_1743;
wire n_3309;
wire n_2075;
wire newNet_1078;
wire n_1360;
wire n_3675;
wire newNet_406;
wire n_4686;
wire n_855;
wire n_2104;
wire newNet_1024;
wire n_4587;
wire R16_11_;
wire n_4251;
wire io_a_5;
wire n_3209;
wire newNet_1295;
wire n_609;
wire n_1808;
wire n_3513;
wire n_1167;
wire n_3704;
wire newNet_1510;
wire n_2288;
wire n_4590;
wire n_558;
wire n_2673;
wire n_3857;
wire n_1177;
wire n_1958;
wire n_2066;
wire n_556;
wire n_1468;
wire n_681;
wire n_2793;
wire n_3589;
wire n_1396;
wire n_1570;
wire newNet_1242;
wire n_127;
wire n_3021;
wire n_4101;
wire n_1797;
wire GPR_17__5_;
wire n_1533;
wire newNet_1654;
wire newNet_8;
wire n_96;
wire n_1140;
wire n_2470;
wire newNet_1276;
wire n_4021;
wire n_2313;
wire n_427;
wire n_519;
wire n_1341;
wire n_366;
wire n_1405;
wire n_3119;
wire io_sp_2_;
wire n_2627;
wire newNet_1170;
wire newNet_228;
wire n_1951;
wire newNet_1140;
wire n_3014;
wire n_1451;
wire n_1096;
wire n_3144;
wire GPR_14__0_;
wire pY_0_;
wire n_4653;
wire newNet_1064;
wire newNet_1052;
wire n_405;
wire newNet_1857;
wire n_2458;
wire n_273;
wire n_3239;
wire n_1875;
wire n_3101;
wire newNet_1012;
wire n_258;
wire newNet_370;
wire newNet_1169;
wire n_4640;
wire newNet_853;
wire n_1649;
wire n_2722;
wire n_2136;
wire n_3224;
wire newNet_56;
wire newNet_1111;
wire n_659;
wire n_1920;
wire pZ_7_;
wire n_1765;
wire n_1653;
wire n_1494;
wire n_3967;
wire n_1870;
wire n_810;
wire newNet_803;
wire n_1337;
wire n_807;
wire n_512;
wire newNet_1029;
wire n_491;
wire n_3138;
wire R16_2_;
wire n_1661;
wire GPR_16__2_;
wire n_3268;
wire n_3085;
wire n_34;
wire newNet_974;
wire newNet_1244;
wire n_2637;
wire n_4627;
wire newNet_39;
wire n_2493;
wire n_2227;
wire n_3436;
wire newNet_1624;
wire newNet_1001;
wire n_3337;
wire n_1616;
wire n_3747;
wire n_317;
wire newNet_1108;
wire n_1289;
wire n_3773;
wire n_3827;
wire n_4282;
wire n_2036;
wire newNet_549;
wire newNet_181;
wire n_1356;
wire n_2971;
wire n_2561;
wire n_2460;
wire n_4041;
wire n_2836;
wire n_3131;
wire n_299;
wire newNet_481;
wire n_2594;
wire n_2340;
wire io_sp_4_;
wire n_778;
wire newNet_1447;
wire n_2776;
wire n_310;
wire n_1697;
wire n_285;
wire GPR_10__7_;
wire n_3039;
wire newNet_221;
wire n_221;
wire n_45;
wire n_2822;
wire n_2981;
wire newNet_1781;
wire newNet_1412;
wire newNet_435;
wire newNet_847;
wire n_284;
wire newNet_288;
wire n_3050;
wire n_4617;
wire C;
wire newNet_814;
wire newNet_628;
wire n_1196;
wire n_2296;
wire newNet_325;
wire n_2156;
wire n_2866;
wire newNet_1032;
wire newNet_565;
wire dmem_di_4;
wire n_2926;
wire n_3413;
wire n_3363;
wire n_4008;
wire n_2599;
wire n_182;
wire n_4293;
wire n_610;
wire newNet_1786;
wire n_714;
wire n_4258;
wire n_225;
wire newNet_299;
wire newNet_587;
wire n_3938;
wire n_862;
wire n_3798;
wire newNet_469;
wire newNet_164;
wire n_2119;
wire n_2168;
wire SP_6_;
wire n_4320;
wire n_80;
wire n_3043;
wire GPR_Rd_r_7_;
wire n_885;
wire n_2362;
wire newNet_515;
wire n_4073;
wire n_425;
wire n_2570;
wire newNet_1371;
wire n_1000;
wire newNet_1317;
wire n_581;
wire n_505;
wire n_1668;
wire newNet_505;
wire n_2519;
wire pY_15_;
wire n_3731;
wire n_1014;
wire n_76;
wire n_728;
wire n_708;
wire n_4026;
wire n_15;
wire n_1041;
wire n_2898;
wire newNet_445;
wire newNet_384;
wire GPR_20__1_;
wire n_863;
wire n_906;
wire n_272;
wire newNet_1441;
wire GPR_17__1_;
wire newNet_884;
wire n_2000;
wire n_619;
wire newNet_1122;
wire n_3893;
wire newNet_1856;
wire newNet_167;
wire n_837;
wire n_3186;
wire n_3174;
wire n_3711;
wire GPR_23__0_;
wire newNet_1212;
wire n_1754;
wire newNet_198;
wire n_3886;
wire n_3994;
wire n_1265;
wire n_4116;
wire n_4451;
wire n_4637;
wire newNet_519;
wire n_539;
wire newNet_537;
wire newNet_1249;
wire n_2469;
wire n_3439;
wire n_2093;
wire n_2788;
wire newNet_679;
wire n_2085;
wire n_4294;
wire newNet_186;
wire n_3685;
wire n_2702;
wire GPR_4__7_;
wire newNet_1134;
wire n_2358;
wire n_2216;
wire n_721;
wire n_1447;
wire io_do_0;
wire n_1515;
wire newNet_1463;
wire n_162;
wire n_1825;
wire n_3475;
wire newNet_1684;
wire n_4184;
wire newNet_861;
wire n_12;
wire newNet_1493;
wire newNet_1392;
wire GPR_13__6_;
wire n_169;
wire n_895;
wire n_688;
wire n_321;
wire n_1015;
wire n_1370;
wire GPR_23__5_;
wire newNet_452;
wire n_2967;
wire n_1174;
wire n_3876;
wire n_3624;
wire n_567;
wire newNet_613;
wire n_2422;
wire n_924;
wire n_1123;
wire n_3803;
wire n_2873;
wire n_946;
wire newNet_734;
wire n_411;
wire n_1379;
wire n_3956;
wire n_2630;
wire n_3891;
wire n_4120;
wire newNet_1716;
wire n_1938;
wire n_261;
wire n_4098;
wire newNet_960;
wire n_2250;
wire newNet_574;
wire newNet_421;
wire newNet_345;
wire GPR_7__0_;
wire n_2853;
wire n_3941;
wire n_1932;
wire newNet_1688;
wire n_2115;
wire n_2125;
wire newNet_310;
wire n_3899;
wire newNet_1795;
wire n_2841;
wire n_869;
wire n_872;
wire newNet_338;
wire newNet_749;
wire n_64;
wire n_1300;
wire n_3009;
wire n_3846;
wire n_4160;
wire n_1947;
wire n_3384;
wire n_2585;
wire n_4082;
wire n_3408;
wire n_3244;
wire n_4303;
wire newNet_725;
wire n_2256;
wire newNet_1046;
wire n_1205;
wire n_2090;
wire n_3579;
wire n_1582;
wire n_3403;
wire n_438;
wire n_766;
wire n_2243;
wire newNet_1133;
wire GPR_3__7_;
wire newNet_1707;
wire n_2237;
wire n_4104;
wire n_2654;
wire n_3762;
wire newNet_323;
wire n_2001;
wire n_1428;
wire n_3175;
wire n_3863;
wire n_3942;
wire n_3980;
wire n_656;
wire n_1772;
wire rst;
wire n_3996;
wire newNet_1326;
wire newNet_211;
wire n_1755;
wire n_3630;
wire n_3717;
wire n_1777;
wire n_1735;
wire n_3705;
wire n_538;
wire n_2379;
wire n_1594;
wire n_2122;
wire newNet_589;
wire newNet_1335;
wire n_4537;
wire n_2273;
wire n_1382;
wire n_3645;
wire n_11;
wire n_1744;
wire n_4390;
wire n_4520;
wire n_670;
wire n_2829;
wire newNet_1605;
wire n_3265;
wire newNet_348;
wire n_3858;
wire n_4330;
wire n_515;
wire n_1236;
wire n_2494;
wire newNet_658;
wire n_3847;
wire newNet_1812;
wire newNet_564;
wire n_1937;
wire newNet_489;
wire n_2631;
wire n_2984;
wire n_180;
wire n_633;
wire n_2265;
wire n_1009;
wire n_3283;
wire newNet_1519;
wire n_612;
wire n_3911;
wire n_1226;
wire n_3557;
wire newNet_422;
wire n_1113;
wire n_3195;
wire n_2634;
wire newNet_1617;
wire n_1795;
wire n_4423;
wire n_1134;
wire n_56;
wire newNet_1188;
wire n_4450;
wire n_2641;
wire n_2774;
wire n_1117;
wire n_2372;
wire final_adder_mux_R16_278_6_n_25;
wire newNet_1206;
wire n_3597;
wire n_3926;
wire n_2281;
wire newNet_1698;
wire newNet_1286;
wire n_1491;
wire n_1065;
wire n_4119;
wire n_1324;
wire n_3661;
wire U_1_;
wire newNet_67;
wire n_1480;
wire n_2131;
wire n_926;
wire n_1030;
wire n_2752;
wire n_3975;
wire n_3344;
wire n_103;
wire newNet_1097;
wire n_293;
wire n_2759;
wire n_1816;
wire GPR_0__1_;
wire n_1213;
wire n_3372;
wire n_2865;
wire n_3217;
wire n_1257;
wire GPR_19__7_;
wire newNet_1544;
wire n_1877;
wire n_2109;
wire dmem_do_0;
wire GPR_9__4_;
wire n_2315;
wire newNet_1694;
wire n_777;
wire n_3270;
wire newNet_1228;
wire newNet_665;
wire newNet_28;
wire n_963;
wire GPR_22__1_;
wire newNet_693;
wire newNet_1372;
wire n_1475;
wire n_3835;
wire newNet_480;
wire newNet_548;
wire newNet_525;
wire n_3036;
wire n_4059;
wire n_966;
wire n_3525;
wire newNet_1551;
wire newNet_514;
wire newNet_379;
wire n_2199;
wire n_328;
wire n_1785;
wire n_4516;
wire newNet_1107;
wire n_3580;
wire n_3637;
wire n_1573;
wire newNet_921;
wire n_1899;
wire n_1378;
wire n_949;
wire n_2604;
wire n_3496;
wire n_1248;
wire n_3146;
wire n_577;
wire GPR_16__5_;
wire n_252;
wire newNet_1280;
wire newNet_1561;
wire n_1957;
wire GPR_Rd_r_2_;
wire newNet_12;
wire newNet_948;
wire newNet_1194;
wire newNet_1057;
wire newNet_1343;
wire newNet_14;
wire n_648;
wire n_2197;
wire n_1149;
wire n_3939;
wire newNet_1674;
wire pmem_d_2;
wire n_3492;
wire n_1762;
wire n_1830;
wire newNet_133;
wire n_3588;
wire n_1203;
wire n_2614;
wire newNet_98;
wire n_2484;
wire n_2804;
wire n_2502;
wire n_454;
wire newNet_206;
wire n_2512;
wire n_4549;
wire n_4183;
wire n_267;
wire n_4530;
wire n_2369;
wire n_4442;
wire n_3590;
wire n_1089;
wire GPR_5__6_;
wire n_3443;
wire n_87;
wire n_3302;
wire newNet_153;
wire n_1973;
wire n_3921;
wire GPR_6__6_;
wire n_2684;
wire n_3377;
wire n_4235;
wire pmem_d_1;
wire n_174;
wire n_3728;
wire newNet_436;
wire n_4207;
wire n_4191;
wire PC_3_;
wire n_2904;
wire n_3746;
wire n_3040;
wire n_3916;
wire n_2544;
wire GPR_2__1_;
wire newNet_262;
wire n_2045;
wire newNet_1756;
wire newNet_405;
wire n_385;
wire newNet_686;
wire newNet_1490;
wire newNet_1015;
wire newNet_758;
wire n_2011;
wire n_2844;
wire newNet_1362;
wire newNet_172;
wire newNet_906;
wire n_1846;
wire newNet_576;
wire newNet_81;
wire GPR_8__3_;
wire n_3987;
wire newNet_820;
wire n_1150;
wire n_1888;
wire newNet_621;
wire n_987;
wire n_3429;
wire n_4046;
wire newNet_250;
wire n_3693;
wire n_4381;
wire final_adder_mux_R16_278_6_n_3;
wire pmem_a_6;
wire n_2886;
wire n_4464;
wire n_1768;
wire n_2418;
wire GPR_12__5_;
wire n_3609;
wire newNet_55;
wire n_2304;
wire newNet_1011;
wire n_355;
wire n_3526;
wire n_2747;
wire n_4055;
wire n_3276;
wire n_3108;
wire n_1389;
wire n_2718;
wire n_1369;
wire n_3058;
wire n_2186;
wire n_1913;
wire n_1982;
wire newNet_1572;
wire n_1698;
wire newNet_1380;
wire newNet_284;
wire newNet_1311;
wire n_1611;
wire newNet_1112;
wire n_1792;
wire newNet_1072;
wire n_3639;
wire n_1068;
wire n_1071;
wire n_3084;
wire final_adder_mux_R16_278_6_n_51;
wire n_3313;
wire n_4555;
wire n_2666;
wire n_4527;
wire n_4089;
wire n_1907;
wire n_4203;
wire n_625;
wire n_1733;
wire n_2430;
wire n_1751;
wire newNet_1593;
wire newNet_827;
wire n_1679;
wire n_1864;
wire n_2954;
wire n_3328;
wire io_di_7;
wire n_908;
wire newNet_764;
wire n_753;
wire n_3463;
wire newNet_1631;
wire newNet_740;
wire n_547;
wire n_134;
wire n_4603;
wire newNet_350;
wire GPR_0__7_;
wire n_1564;
wire newNet_896;
wire n_545;
wire n_1419;
wire n_483;
wire n_3122;
wire newNet_416;
wire n_3367;
wire n_1303;
wire newNet_1087;
wire GPR_13__5_;
wire n_3051;
wire newNet_1158;
wire n_2761;
wire newNet_1476;
wire n_1159;
wire n_3547;
wire final_adder_mux_R16_278_6_n_36;
wire n_2405;
wire n_4666;
wire newNet_44;
wire newNet_932;
wire n_1085;
wire n_3554;
wire n_4216;
wire newNet_584;
wire n_2029;
wire newNet_1587;
wire n_197;
wire newNet_1254;
wire newNet_918;
wire newNet_1505;
wire n_1837;
wire n_4066;
wire n_1716;
wire n_4245;
wire newNet_1141;
wire GPR_8__0_;
wire n_993;
wire newNet_1808;
wire newNet_78;
wire state_3_;
wire newNet_1091;
wire GPR_5__5_;
wire n_1684;
wire newNet_989;
wire n_1195;
wire n_4349;
wire n_3954;
wire n_1800;
wire newNet_1776;
wire n_4232;
wire n_397;
wire final_adder_mux_R16_278_6_n_1;
wire newNet_1219;
wire n_202;
wire n_525;
wire n_3416;
wire newNet_1558;
wire newNet_955;
wire n_4379;
wire n_2183;
wire n_3071;
wire n_3755;
wire n_3726;
wire n_1558;
wire newNet_1747;
wire n_3518;
wire n_3292;
wire n_3028;
wire newNet_962;
wire n_2750;
wire n_829;
wire newNet_783;
wire n_378;
wire newNet_559;
wire newNet_1728;
wire n_2558;
wire n_4685;
wire n_4611;
wire n_608;
wire n_784;
wire n_732;
wire n_2389;
wire n_3818;
wire newNet_199;
wire n_3321;
wire newNet_235;
wire newNet_1374;
wire newNet_10;
wire n_990;
wire n_980;
wire n_1471;
wire newNet_1740;
wire n_75;
wire n_1090;
wire newNet_1318;
wire n_3315;
wire n_1636;
wire n_3504;
wire newNet_1862;
wire n_4343;
wire newNet_1073;
wire newNet_1381;
wire n_750;
wire n_3345;
wire n_3250;
wire n_2254;
wire n_25;
wire n_3877;
wire final_adder_mux_R16_278_6_n_4;
wire n_4633;
wire final_adder_mux_R16_278_6_n_2;
wire n_701;
wire newNet_1831;
wire n_4646;
wire newNet_83;
wire n_3923;
wire Rd_3_;
wire n_1505;
wire n_410;
wire n_3414;
wire newNet_623;
wire newNet_731;
wire n_1963;
wire n_274;
wire newNet_780;
wire newNet_575;
wire n_326;
wire newNet_1638;
wire newNet_353;
wire n_1459;
wire newNet_774;
wire n_373;
wire newNet_1645;
wire newNet_727;
wire newNet_92;
wire newNet_19;
wire n_3523;
wire n_1617;
wire newNet_769;
wire n_601;
wire newNet_1199;
wire n_4478;
wire newNet_995;
wire n_1034;
wire n_2687;
wire newNet_1084;
wire newNet_1334;
wire n_736;
wire pmem_a_8;
wire n_1721;
wire newNet_961;
wire n_2401;
wire n_1586;
wire newNet_433;
wire n_3354;
wire n_249;
wire n_2854;
wire newNet_256;
wire n_3741;
wire n_3291;
wire n_1708;
wire n_332;
wire n_2492;
wire n_2830;
wire newNet_99;
wire n_165;
wire n_3280;
wire io_di_0;
wire n_3754;
wire n_1736;
wire newNet_237;
wire SP_3_;
wire n_363;
wire n_2382;
wire n_3965;
wire n_3338;
wire n_1130;
wire n_4283;
wire newNet_339;
wire newNet_268;
wire newNet_369;
wire n_3735;
wire newNet_894;
wire n_4522;
wire newNet_365;
wire newNet_1110;
wire newNet_817;
wire n_372;
wire n_2681;
wire n_147;
wire n_1673;
wire n_1232;
wire n_4358;
wire n_3201;
wire newNet_761;
wire n_3562;
wire newNet_883;
wire n_1228;
wire n_3628;
wire newNet_244;
wire n_4240;
wire n_1197;
wire newNet_1255;
wire newNet_261;
wire n_2181;
wire n_2914;
wire n_1914;
wire newNet_594;
wire n_2529;
wire n_4470;
wire n_1553;
wire n_780;
wire n_2650;
wire n_1432;
wire n_1834;
wire n_1139;
wire newNet_29;
wire n_4399;
wire PC_5_;
wire newNet_1778;
wire newNet_660;
wire n_349;
wire n_359;
wire newNet_757;
wire newNet_873;
wire newNet_1321;
wire newNet_260;
wire n_1107;
wire n_44;
wire n_2276;
wire n_537;
wire newNet_821;
wire n_2825;
wire n_1700;
wire n_1681;
wire n_1790;
wire n_1055;
wire n_3512;
wire newNet_1013;
wire n_2743;
wire n_3474;
wire newNet_271;
wire newNet_1327;
wire n_1024;
wire n_4127;
wire n_578;
wire n_383;
wire n_4214;
wire n_1562;
wire newNet_1555;
wire n_152;
wire n_1153;
wire n_4247;
wire n_2162;
wire n_2677;
wire n_838;
wire n_1222;
wire newNet_1816;
wire n_4065;
wire newNet_913;
wire n_1896;
wire n_1719;
wire newNet_788;
wire newNet_385;
wire n_2010;
wire n_4468;
wire newNet_790;
wire newNet_1737;
wire n_3953;
wire n_3644;
wire n_296;
wire n_1399;
wire n_4628;
wire newNet_1360;
wire n_4200;
wire newNet_1582;
wire n_3422;
wire n_1809;
wire n_3449;
wire n_2018;
wire n_2361;
wire n_3852;
wire newNet_879;
wire n_4139;
wire n_1939;
wire newNet_1532;
wire n_3723;
wire newNet_312;
wire newNet_691;
wire n_3585;
wire n_2757;
wire n_3985;
wire n_1464;
wire n_1778;
wire n_3831;
wire n_334;
wire n_3409;
wire n_303;
wire n_257;
wire io_sp_1_;
wire n_1214;
wire newNet_975;
wire n_2137;
wire n_718;
wire n_1575;
wire n_735;
wire n_3838;
wire n_3491;
wire newNet_1063;
wire n_1084;
wire n_2215;
wire n_4170;
wire n_2868;
wire n_621;
wire GPR_2__5_;
wire n_437;
wire n_104;
wire n_4056;
wire n_972;
wire newNet_1267;
wire n_1801;
wire n_1933;
wire n_1521;
wire n_4194;
wire n_4052;
wire n_2962;
wire n_1596;
wire n_3225;
wire newNet_1135;
wire n_916;
wire newNet_1750;
wire n_2636;
wire n_1536;
wire newNet_1454;
wire n_1298;
wire newNet_1691;
wire newNet_205;
wire n_3374;
wire n_2937;
wire GPR_0__4_;
wire n_2740;
wire n_3139;
wire n_1786;
wire newNet_316;
wire newNet_743;
wire n_1063;
wire pX_10_;
wire newNet_922;
wire PC_7_;
wire n_2501;
wire n_3349;
wire n_2481;
wire dmem_di_6;
wire n_2468;
wire n_3480;
wire n_1746;
wire newNet_376;
wire GPR_20__7_;
wire newNet_1222;
wire n_658;
wire newNet_1250;
wire n_4;
wire io_di_5;
wire n_1211;
wire n_3772;
wire n_264;
wire n_3495;
wire n_1986;
wire n_1108;
wire n_269;
wire newNet_797;
wire n_914;
wire newNet_106;
wire n_1710;
wire GPR_20__0_;
wire n_2393;
wire n_1660;
wire newNet_1117;
wire n_217;
wire n_618;
wire n_3912;
wire n_2420;
wire n_2688;
wire newNet_1501;
wire n_57;
wire n_3277;
wire n_3909;
wire n_236;
wire n_743;
wire n_445;
wire n_2922;
wire n_3004;
wire n_3660;
wire n_3155;
wire n_2806;
wire n_587;
wire final_adder_mux_R16_278_6_n_32;
wire n_4336;
wire newNet_1419;
wire n_2930;
wire n_2657;
wire n_639;
wire n_3038;
wire n_3930;
wire n_2290;
wire n_452;
wire newNet_1695;
wire n_4177;
wire n_2284;
wire n_3272;
wire n_3667;
wire n_4332;
wire n_2328;
wire newNet_1603;
wire newNet_1538;
wire n_1861;
wire n_4593;
wire n_3379;
wire n_3306;
wire n_968;
wire n_3635;
wire n_1976;
wire n_1688;
wire n_2542;
wire n_3966;
wire n_2240;
wire newNet_543;
wire n_779;
wire n_2171;
wire newNet_1287;
wire n_1974;
wire n_4614;
wire newNet_1542;
wire newNet_1344;
wire newNet_902;
wire n_3596;
wire newNet_598;
wire n_3243;
wire n_1995;
wire newNet_49;
wire n_2996;
wire n_2781;
wire n_28;
wire n_765;
wire newNet_1190;
wire n_2771;
wire newNet_602;
wire n_181;
wire newNet_1040;
wire newNet_1031;
wire newNet_1346;
wire n_1307;
wire newNet_1568;
wire n_2009;
wire n_348;
wire newNet_1439;
wire n_2785;
wire GPR_10__6_;
wire n_1144;
wire n_1959;
wire n_2107;
wire n_1478;
wire newNet_141;
wire n_4559;
wire n_930;
wire n_3558;
wire n_2709;
wire n_2500;
wire n_2892;
wire newNet_1708;
wire n_4070;
wire n_2268;
wire newNet_1055;
wire n_1081;
wire n_1110;
wire n_925;
wire newNet_1216;
wire n_1780;
wire GPR_11__4_;
wire n_419;
wire n_3993;
wire n_1246;
wire n_1088;
wire newNet_1367;
wire n_1696;
wire GPR_18__7_;
wire n_86;
wire n_1878;
wire newNet_202;
wire n_2202;
wire newNet_1549;
wire newNet_187;
wire n_1070;
wire n_2034;
wire n_4198;
wire GPR_8__5_;
wire n_3149;
wire n_2076;
wire n_2958;
wire newNet_1089;
wire newNet_448;
wire n_50;
wire n_1902;
wire n_3607;
wire n_1323;
wire n_3503;
wire n_2062;
wire newNet_134;
wire n_482;
wire newNet_558;
wire n_865;
wire newNet_315;
wire n_722;
wire n_4161;
wire n_3519;
wire newNet_678;
wire n_3708;
wire newNet_7;
wire newNet_1227;
wire GPR_21__7_;
wire n_3542;
wire n_3093;
wire n_1018;
wire n_3659;
wire n_2096;
wire n_2008;
wire n_188;
wire n_1968;
wire newNet_637;
wire n_3734;
wire n_4638;
wire n_1537;
wire n_843;
wire n_948;
wire newNet_1126;
wire newNet_1859;
wire newNet_61;
wire newNet_162;
wire n_2412;
wire n_951;
wire newNet_155;
wire n_676;
wire n_3678;
wire newNet_895;
wire n_4586;
wire n_3896;
wire n_4651;
wire n_1019;
wire n_879;
wire SP_7_;
wire n_3103;
wire n_3136;
wire n_148;
wire PC_1_;
wire newNet_1398;
wire n_941;
wire n_2543;
wire n_3154;
wire n_4006;
wire n_3819;
wire n_2026;
wire n_898;
wire n_2230;
wire newNet_1533;
wire newNet_577;
wire n_74;
wire n_120;
wire final_adder_mux_R16_278_6_n_77;
wire n_1367;
wire n_3890;
wire newNet_1391;
wire newNet_1120;
wire n_3551;
wire n_2876;
wire n_1275;
wire io_sp_7_;
wire n_851;
wire n_4322;
wire n_1745;
wire newNet_459;
wire n_1934;
wire n_568;
wire newNet_30;
wire newNet_21;
wire newNet_666;
wire n_2058;
wire n_1194;
wire n_4417;
wire newNet_823;
wire n_3888;
wire n_39;
wire n_2921;
wire n_1427;
wire GPR_11__6_;
wire newNet_1830;
wire U_2_;
wire n_2593;
wire newNet_1444;
wire n_1506;
wire n_2207;
wire n_1695;
wire newNet_1449;
wire n_1518;
wire n_4486;
wire n_2557;
wire newNet_123;
wire newNet_1373;
wire final_adder_mux_R16_278_6_n_33;
wire n_3943;
wire GPR_8__1_;
wire newNet_1769;
wire newNet_1594;
wire newNet_324;
wire newNet_222;
wire pY_6_;
wire n_386;
wire n_3168;
wire n_4154;
wire n_2566;
wire n_1439;
wire n_2088;
wire n_1098;
wire newNet_963;
wire n_4111;
wire newNet_675;
wire newNet_326;
wire n_271;
wire n_3041;
wire n_1773;
wire newNet_701;
wire n_65;
wire newNet_70;
wire newNet_289;
wire n_4437;
wire n_2550;
wire n_2221;
wire n_1456;
wire R16_0_;
wire newNet_1312;
wire n_304;
wire n_1170;
wire n_1654;
wire n_3184;
wire n_719;
wire n_4001;
wire newNet_428;
wire n_3070;
wire n_347;
wire n_620;
wire GPR_22__0_;
wire n_2191;
wire newNet_886;
wire final_adder_mux_R16_278_6_n_50;
wire n_3810;
wire n_793;
wire n_1549;
wire newNet_1434;
wire n_2297;
wire newNet_1045;
wire newNet_18;
wire n_1887;
wire n_1254;
wire n_2564;
wire n_1079;
wire n_3477;
wire newNet_1837;
wire n_1291;
wire n_4656;
wire n_320;
wire newNet_77;
wire n_2246;
wire n_3795;
wire newNet_1789;
wire n_4091;
wire newNet_1277;
wire n_3913;
wire n_4547;
wire n_4047;
wire n_3636;
wire newNet_1166;
wire newNet_1155;
wire newNet_1431;
wire n_1066;
wire n_1589;
wire GPR_0__0_;
wire n_2928;
wire n_1769;
wire n_3286;
wire n_880;
wire n_2667;
wire newNet_1096;
wire newNet_655;
wire newNet_290;
wire n_2895;
wire n_3682;
wire n_469;
wire newNet_1248;
wire n_1852;
wire newNet_1518;
wire n_1001;
wire newNet_943;
wire n_4422;
wire pZ_5_;
wire n_402;
wire n_2428;
wire n_2151;
wire n_1241;
wire n_932;
wire newNet_184;
wire n_3016;
wire n_3511;
wire n_3266;
wire newNet_849;
wire n_642;
wire dmem_di_5;
wire n_3610;
wire n_1646;
wire n_1036;
wire newNet_1459;
wire n_516;
wire GPR_3__4_;
wire newNet_709;
wire n_859;
wire n_4443;
wire n_1727;
wire n_3650;
wire n_1793;
wire n_858;
wire n_2762;
wire n_1352;
wire n_2941;
wire newNet_1404;
wire n_4246;
wire GPR_23__7_;
wire U_8_;
wire newNet_1847;
wire newNet_1028;
wire n_3202;
wire newNet_1625;
wire n_3382;
wire n_204;
wire n_3033;
wire n_2579;
wire n_4600;
wire n_3267;
wire n_1316;
wire n_4016;
wire n_198;
wire newNet_1815;
wire GPR_11__2_;
wire n_891;
wire n_2611;
wire newNet_1513;
wire newNet_632;
wire n_2880;
wire n_4591;
wire n_2312;
wire n_465;
wire n_1143;
wire n_4566;
wire n_2050;
wire newNet_1777;
wire n_4684;
wire n_1703;
wire newNet_1428;
wire n_3462;
wire n_1632;
wire newNet_493;
wire n_3216;
wire n_230;
wire n_2523;
wire n_2575;
wire n_2196;
wire newNet_1106;
wire GPR_20__5_;
wire n_2182;
wire n_4022;
wire n_3714;
wire n_661;
wire n_696;
wire n_2959;
wire n_1601;
wire newNet_844;
wire GPR_18__3_;
wire n_2736;
wire n_3232;
wire U_4_;
wire n_2069;
wire n_2459;
wire n_1281;
wire n_4373;
wire GPR_11__3_;
wire n_3563;
wire n_3600;
wire newNet_866;
wire newNet_1637;
wire n_371;
wire n_1104;
wire newNet_1217;
wire n_1342;
wire newNet_583;
wire n_1556;
wire n_4400;
wire newNet_842;
wire newNet_371;
wire n_1359;
wire newNet_471;
wire n_3870;
wire SP_8_;
wire n_3160;
wire newNet_1682;
wire n_417;
wire n_4199;
wire n_2727;
wire newNet_775;
wire n_4328;
wire n_2618;
wire newNet_229;
wire n_1120;
wire n_2975;
wire newNet_516;
wire n_1495;
wire n_171;
wire n_649;
wire n_3022;
wire n_2123;
wire n_4368;
wire newNet_1058;
wire n_3577;
wire io_sp_0_;
wire n_495;
wire n_1411;
wire n_3865;
wire n_1288;
wire n_2320;
wire n_2931;
wire n_4144;
wire newNet_1328;
wire n_1927;
wire n_555;
wire n_1876;
wire n_2344;
wire n_2586;
wire n_99;
wire n_1880;
wire n_2353;
wire n_1542;
wire n_1952;
wire n_1763;
wire n_4663;
wire n_1375;
wire n_2334;
wire newNet_1022;
wire n_3538;
wire n_3841;
wire newNet_1852;
wire newNet_20;
wire n_3029;
wire n_2675;
wire n_1165;
wire n_2017;
wire n_3881;
wire n_18;
wire newNet_212;
wire newNet_1726;
wire n_173;
wire n_1168;
wire n_1332;
wire n_3226;
wire n_981;
wire newNet_1497;
wire newNet_1180;
wire newNet_986;
wire newNet_501;
wire newNet_1355;
wire n_824;
wire n_4136;
wire newNet_717;
wire n_2144;
wire n_1385;
wire newNet_744;
wire n_4421;
wire n_2692;
wire n_251;
wire n_2491;
wire n_3030;
wire n_3617;
wire final_adder_mux_R16_278_6_n_24;
wire n_492;
wire newNet_991;
wire n_594;
wire newNet_622;
wire n_3082;
wire n_3671;
wire n_4403;
wire n_3533;
wire newNet_456;
wire n_3063;
wire n_585;
wire n_4620;
wire n_2845;
wire newNet_1826;
wire n_4171;
wire n_591;
wire newNet_1298;
wire newNet_402;
wire n_2395;
wire n_2901;
wire newNet_43;
wire newNet_1736;
wire n_2690;
wire n_327;
wire n_1262;
wire newNet_756;
wire n_4224;
wire n_2198;
wire n_4254;
wire n_1404;
wire n_2605;
wire n_1595;
wire newNet_148;
wire n_4389;
wire n_600;
wire n_2450;
wire n_1998;
wire n_1245;
wire newNet_440;
wire n_4028;
wire newNet_1008;
wire n_3194;
wire n_2444;
wire n_4034;
wire newNet_1150;
wire pX_9_;
wire GPR_18__5_;
wire n_3339;
wire n_3392;
wire newNet_1573;
wire newNet_1609;
wire newNet_1205;
wire n_2371;
wire n_2658;
wire n_2983;
wire n_1720;
wire n_2446;
wire n_2112;
wire newNet_916;
wire n_137;
wire n_3112;
wire n_1828;
wire n_3782;
wire newNet_1408;
wire n_129;
wire n_1400;
wire n_241;
wire n_3400;
wire n_2515;
wire n_4479;
wire n_3320;
wire n_2706;
wire n_3531;
wire n_2438;
wire n_4280;
wire newNet_1779;
wire newNet_912;
wire n_1791;
wire n_4044;
wire newNet_79;
wire n_4471;
wire n_2828;
wire GPR_4__3_;
wire n_2180;
wire n_3627;
wire n_331;
wire n_3749;
wire n_189;
wire n_1431;
wire n_2938;
wire newNet_413;
wire n_647;
wire newNet_818;
wire n_1193;
wire n_353;
wire n_1172;
wire newNet_292;
wire n_2680;
wire newNet_874;
wire n_3489;
wire n_1839;
wire n_3448;
wire n_4071;
wire n_2429;
wire GPR_7__3_;
wire dmem_we;
wire n_4248;
wire n_3964;
wire n_3278;
wire n_2366;
wire n_1779;
wire n_2820;
wire n_1565;
wire n_1833;
wire newNet_1515;
wire n_395;
wire newNet_1662;
wire newNet_1034;
wire n_2235;
wire n_3059;
wire n_4201;
wire n_1056;
wire n_763;
wire newNet_1014;
wire newNet_604;
wire n_2535;
wire n_2616;
wire n_478;
wire n_2676;
wire n_3932;
wire n_1915;
wire newNet_214;
wire n_1718;
wire newNet_279;
wire n_3113;
wire newNet_201;
wire n_151;
wire newNet_140;
wire n_1037;
wire newNet_789;
wire n_1152;
wire n_1484;
wire n_527;
wire newNet_1322;
wire n_4287;
wire n_4215;
wire newNet_1361;
wire n_3902;
wire n_2749;
wire n_4355;
wire GPR_18__1_;
wire newNet_791;
wire n_4302;
wire n_1637;
wire n_3952;
wire n_3516;
wire GPR_0__6_;
wire n_1707;
wire n_300;
wire newNet_1319;
wire n_3740;
wire n_3992;
wire n_1510;
wire n_561;
wire GPR_19__4_;
wire n_2517;
wire newNet_572;
wire newNet_534;
wire n_1239;
wire n_1457;
wire newNet_1562;
wire n_418;
wire n_1131;
wire newNet_234;
wire n_3757;
wire n_3172;
wire n_2255;
wire n_2530;
wire n_809;
wire n_3322;
wire n_1869;
wire newNet_582;
wire n_190;
wire n_665;
wire newNet_732;
wire n_170;
wire newNet_1388;
wire newNet_726;
wire newNet_1495;
wire n_3878;
wire n_3346;
wire newNet_1470;
wire n_3692;
wire n_3944;
wire n_2708;
wire n_2686;
wire n_3417;
wire newNet_1757;
wire newNet_958;
wire newNet_798;
wire n_991;
wire n_3251;
wire n_2046;
wire n_2134;
wire final_adder_mux_R16_278_6_n_5;
wire n_166;
wire GPR_4__2_;
wire newNet_522;
wire n_3423;
wire n_2027;
wire newNet_599;
wire n_1552;
wire n_2241;
wire newNet_1507;
wire newNet_368;
wire n_1121;
wire n_4521;
wire newNet_1333;
wire newNet_1832;
wire newNet_1160;
wire n_3724;
wire pmem_a_7;
wire n_2902;
wire newNet_856;
wire newNet_781;
wire newNet_1256;
wire newNet_1048;
wire n_2620;
wire n_2128;
wire n_827;
wire newNet_893;
wire n_3509;
wire n_2537;
wire newNet_364;
wire n_3594;
wire n_325;
wire n_312;
wire n_4629;
wire n_1926;
wire n_4106;
wire newNet_742;
wire n_3355;
wire newNet_1071;
wire newNet_1613;
wire n_2855;
wire newNet_352;
wire U_3_;
wire n_2716;
wire n_2993;
wire newNet_1074;
wire newNet_236;
wire newNet_122;
wire n_146;
wire n_1994;
wire newNet_267;
wire n_364;
wire dmem_do_3;
wire S;
wire n_2283;
wire newNet_1230;
wire n_2583;
wire n_3929;
wire n_4178;
wire n_2356;
wire n_3576;
wire newNet_1543;
wire n_3005;
wire newNet_901;
wire newNet_1236;
wire GPR_8__7_;
wire newNet_1574;
wire n_2082;
wire newNet_542;
wire n_1207;
wire n_3866;
wire newNet_545;
wire newNet_245;
wire newNet_330;
wire newNet_48;
wire newNet_42;
wire n_58;
wire n_2656;
wire newNet_903;
wire PC_6_;
wire n_1975;
wire n_2077;
wire newNet_639;
wire newNet_107;
wire n_631;
wire n_975;
wire n_1217;
wire n_3643;
wire n_4335;
wire newNet_434;
wire final_adder_mux_R16_278_6_n_15;
wire n_764;
wire n_3908;
wire n_4268;
wire n_2541;
wire n_453;
wire newNet_52;
wire dmem_a_12;
wire n_3406;
wire n_1689;
wire n_2061;
wire n_2913;
wire newNet_1288;
wire n_2974;
wire newNet_1701;
wire newNet_393;
wire n_235;
wire n_3595;
wire n_1862;
wire n_3931;
wire n_3242;
wire U_5_;
wire newNet_1696;
wire n_1614;
wire n_3830;
wire n_219;
wire newNet_1619;
wire newNet_1793;
wire n_51;
wire newNet_1121;
wire n_1002;
wire n_4560;
wire n_751;
wire n_4078;
wire pY_4_;
wire newNet_1281;
wire n_1446;
wire n_4558;
wire n_643;
wire n_1111;
wire n_2891;
wire n_2867;
wire n_85;
wire n_4532;
wire newNet_1191;
wire newNet_192;
wire newNet_656;
wire n_279;
wire n_4117;
wire n_4063;
wire newNet_822;
wire n_1023;
wire newNet_1539;
wire n_931;
wire n_2056;
wire n_1398;
wire newNet_829;
wire n_3817;
wire newNet_1709;
wire newNet_1148;
wire newNet_643;
wire n_636;
wire n_4585;
wire n_1477;
wire n_4539;
wire newNet_603;
wire newNet_1105;
wire n_2950;
wire n_2472;
wire n_3540;
wire n_4057;
wire n_3305;
wire n_2643;
wire n_1087;
wire n_2033;
wire newNet_1569;
wire n_3559;
wire n_4567;
wire n_2986;
wire newNet_1725;
wire GPR_19__0_;
wire n_4278;
wire n_2161;
wire pmem_d_3;
wire n_4149;
wire n_1247;
wire n_4197;
wire n_2200;
wire newNet_118;
wire n_632;
wire n_2786;
wire n_207;
wire n_2106;
wire newNet_1479;
wire newNet_1418;
wire n_3502;
wire n_1977;
wire n_3329;
wire final_adder_mux_R16_278_6_n_27;
wire pZ_13_;
wire n_3606;
wire n_4534;
wire newNet_1741;
wire final_adder_mux_R16_278_6_n_40;
wire n_1987;
wire n_2510;
wire newNet_1268;
wire n_2267;
wire n_1220;
wire n_1802;
wire n_536;
wire n_32;
wire n_3771;
wire n_263;
wire newNet_925;
wire n_3700;
wire n_1520;
wire n_1200;
wire final_adder_mux_R16_278_6_n_71;
wire n_4445;
wire newNet_100;
wire n_915;
wire n_1078;
wire n_758;
wire n_4514;
wire n_436;
wire n_1644;
wire newNet_1748;
wire pX_4_;
wire n_2772;
wire GPR_17__3_;
wire n_3490;
wire n_2095;
wire n_1083;
wire newNet_555;
wire n_105;
wire newNet_54;
wire n_4594;
wire n_801;
wire n_917;
wire newNet_1167;
wire n_3493;
wire n_1905;
wire n_1064;
wire newNet_1197;
wire newNet_683;
wire n_2698;
wire newNet_473;
wire n_2302;
wire n_27;
wire n_3371;
wire newNet_208;
wire newNet_1345;
wire n_4472;
wire n_1391;
wire n_333;
wire newNet_377;
wire n_1255;
wire n_548;
wire newNet_1692;
wire n_2758;
wire n_1212;
wire newNet_22;
wire n_1737;
wire newNet_1204;
wire n_3148;
wire n_4541;
wire n_94;
wire n_3494;
wire newNet_680;
wire newNet_311;
wire n_216;
wire n_1961;
wire n_1311;
wire n_1535;
wire n_2720;
wire n_4650;
wire final_adder_mux_R16_278_6_n_60;
wire n_1450;
wire n_572;
wire n_700;
wire n_2349;
wire newNet_1767;
wire n_446;
wire n_1663;
wire newNet_1224;
wire n_3141;
wire n_1655;
wire newNet_976;
wire n_2508;
wire newNet_1221;
wire newNet_455;
wire n_3825;
wire n_4529;
wire n_3586;
wire newNet_1735;
wire n_1109;
wire n_3837;
wire n_4019;
wire newNet_1606;
wire GPR_Rd_r_1_;
wire n_2482;
wire n_3;
wire n_3294;
wire newNet_1838;
wire n_1290;
wire n_4000;
wire n_2208;
wire n_3880;
wire n_2846;
wire n_857;
wire n_3469;
wire n_1445;
wire n_4420;
wire n_259;
wire n_1851;
wire n_1240;
wire n_17;
wire n_887;
wire n_3605;
wire newNet_1644;
wire n_1662;
wire n_2298;
wire n_2113;
wire n_4292;
wire n_2364;
wire newNet_885;
wire n_3651;
wire n_2860;
wire newNet_223;
wire n_43;
wire n_2563;
wire n_1351;
wire n_3683;
wire n_2150;
wire newNet_1589;
wire n_4615;
wire n_1940;
wire newNet_1081;
wire n_4169;
wire newNet_1768;
wire newNet_427;
wire n_2565;
wire n_554;
wire n_627;
wire newNet_1095;
wire n_33;
wire n_4569;
wire n_1358;
wire n_1343;
wire n_270;
wire newNet_1306;
wire n_4109;
wire n_3811;
wire n_2190;
wire n_2170;
wire newNet_908;
wire n_873;
wire newNet_968;
wire newNet_629;
wire n_1306;
wire n_4297;
wire n_4551;
wire n_163;
wire n_2451;
wire n_400;
wire n_2437;
wire newNet_1278;
wire n_3412;
wire n_573;
wire n_757;
wire n_4444;
wire n_4193;
wire n_1187;
wire n_831;
wire n_3106;
wire newNet_708;
wire n_1686;
wire n_1873;
wire n_187;
wire newNet_1007;
wire n_358;
wire n_468;
wire n_1984;
wire n_145;
wire n_1050;
wire newNet_1368;
wire newNet_62;
wire n_3024;
wire n_2929;
wire GPR_16__1_;
wire n_4659;
wire n_352;
wire n_3765;
wire n_2222;
wire n_1726;
wire newNet_1247;
wire newNet_935;
wire n_3816;
wire n_792;
wire n_1230;
wire n_821;
wire n_1827;
wire n_933;
wire n_4360;
wire newNet_1462;
wire n_4090;
wire n_1310;
wire n_4053;
wire n_4135;
wire newNet_977;
wire newNet_942;
wire n_4592;
wire n_2331;
wire newNet_1210;
wire newNet_327;
wire newNet_1433;
wire n_2896;
wire n_2942;
wire n_136;
wire n_1859;
wire newNet_1151;
wire n_394;
wire n_3622;
wire n_2007;
wire newNet_447;
wire n_1960;
wire newNet_517;
wire newNet_1655;
wire n_890;
wire n_3801;
wire n_4630;
wire n_3304;
wire newNet_196;
wire n_2068;
wire n_2835;
wire newNet_677;
wire n_2961;
wire n_4683;
wire n_1969;
wire newNet_1700;
wire n_1470;
wire n_1490;
wire n_3137;
wire n_1017;
wire n_339;
wire n_844;
wire n_904;
wire GPR_9__5_;
wire newNet_185;
wire n_940;
wire n_63;
wire n_723;
wire newNet_270;
wire n_4321;
wire newNet_1218;
wire n_3733;
wire n_3233;
wire newNet_1486;
wire n_4155;
wire n_283;
wire n_697;
wire n_1694;
wire newNet_154;
wire n_4009;
wire n_1263;
wire n_2721;
wire newNet_1240;
wire n_1376;
wire n_3928;
wire n_734;
wire n_3530;
wire newNet_1270;
wire n_2691;
wire n_4023;
wire n_2589;
wire newNet_1787;
wire newNet_1196;
wire newNet_824;
wire n_199;
wire n_4128;
wire n_3161;
wire n_2875;
wire newNet_420;
wire newNet_1825;
wire final_adder_mux_R16_278_6_n_34;
wire n_1027;
wire n_2782;
wire newNet_699;
wire n_1042;
wire n_504;
wire SP_1_;
wire n_3905;
wire n_1274;
wire newNet_1492;
wire n_2341;
wire newNet_1390;
wire n_3454;
wire newNet_1417;
wire n_686;
wire n_593;
wire newNet_1469;
wire n_4416;
wire n_689;
wire newNet_1410;
wire newNet_165;
wire n_2275;
wire newNet_1671;
wire n_1670;
wire n_1473;
wire newNet_1556;
wire pX_11_;
wire n_111;
wire n_73;
wire n_1935;
wire n_121;
wire n_569;
wire newNet_458;
wire n_1366;
wire n_280;
wire n_679;
wire newNet_1443;
wire newNet_31;
wire n_118;
wire n_3840;
wire n_3543;
wire n_897;
wire n_2471;
wire n_1747;
wire n_16;
wire n_4114;
wire n_2951;
wire newNet_863;
wire n_2467;
wire newNet_1714;
wire n_3629;
wire n_489;
wire n_1517;
wire n_1171;
wire n_1166;
wire n_4436;
wire newNet_792;
wire newNet_616;
wire n_3670;
wire n_4402;
wire n_2644;
wire n_2103;
wire n_4077;
wire newNet_990;
wire newNet_6;
wire n_4309;
wire n_2693;
wire n_2374;
wire n_705;
wire n_1832;
wire n_2516;
wire newNet_500;
wire n_3849;
wire n_2639;
wire n_2490;
wire newNet_595;
wire io_do_5;
wire n_2145;
wire n_2621;
wire newNet_1407;
wire n_1665;
wire newNet_1429;
wire n_3532;
wire n_1581;
wire newNet_475;
wire n_3169;
wire newNet_1669;
wire newNet_987;
wire newNet_69;
wire n_4329;
wire n_3083;
wire n_1647;
wire n_66;
wire n_1331;
wire newNet_1262;
wire newNet_1;
wire pY_9_;
wire newNet_213;
wire n_3062;
wire n_2179;
wire newNet_266;
wire newNet_1498;
wire n_4080;
wire n_3897;
wire newNet_1183;
wire newNet_1050;
wire newNet_994;
wire newNet_980;
wire newNet_552;
wire GPR_0__3_;
wire n_4485;
wire n_2445;
wire newNet_147;
wire n_428;
wire newNet_1506;
wire newNet_300;
wire n_517;
wire GPR_6__7_;
wire n_1403;
wire n_3784;
wire n_1465;
wire n_4253;
wire n_3471;
wire newNet_566;
wire n_254;
wire n_646;
wire n_4179;
wire n_2443;
wire newNet_1354;
wire n_4639;
wire n_3285;
wire n_238;
wire n_791;
wire R16_15_;
wire GPR_20__6_;
wire n_1588;
wire n_4223;
wire newNet_1136;
wire n_3656;
wire n_1132;
wire n_998;
wire n_3618;
wire n_2791;
wire n_242;
wire newNet_700;
wire n_240;
wire n_2020;
wire n_4281;
wire n_3486;
wire n_403;
wire n_4601;
wire n_4350;
wire n_2856;
wire n_3783;
wire newNet_1581;
wire newNet_1297;
wire n_4064;
wire n_3707;
wire GPR_2__7_;
wire n_3713;
wire n_4181;
wire newNet_1125;
wire n_2524;
wire n_464;
wire newNet_809;
wire n_660;
wire n_1953;
wire newNet_642;
wire n_2404;
wire n_4103;
wire newNet_490;
wire pmem_d_10;
wire n_1287;
wire n_319;
wire n_4162;
wire newNet_135;
wire n_3023;
wire n_3092;
wire Rd_r_1_;
wire n_617;
wire n_1879;
wire newNet_86;
wire n_3851;
wire n_4584;
wire n_1523;
wire newNet_1403;
wire n_2576;
wire newNet_1427;
wire n_2311;
wire n_1496;
wire n_1590;
wire n_295;
wire n_1704;
wire newNet_1626;
wire newNet_1375;
wire newNet_839;
wire n_2039;
wire n_416;
wire newNet_649;
wire newNet_1527;
wire n_3215;
wire n_579;
wire n_588;
wire n_2410;
wire newNet_1814;
wire n_370;
wire n_3208;
wire n_4429;
wire n_2396;
wire GPR_4__1_;
wire newNet_512;
wire n_1280;
wire n_1322;
wire newNet_1719;
wire newNet_945;
wire n_3124;
wire n_3401;
wire n_3918;
wire GPR_17__4_;
wire newNet_403;
wire newNet_1451;
wire n_3871;
wire n_1105;
wire n_4397;
wire GPR_1__4_;
wire newNet_815;
wire newNet_1422;
wire n_4286;
wire newNet_535;
wire n_172;
wire n_703;
wire newNet_1171;
wire n_2735;
wire newNet_1027;
wire newNet_470;
wire n_2596;
wire n_2619;
wire newNet_663;
wire dmem_a_3;
wire n_4621;
wire n_4143;
wire n_493;
wire newNet_1512;
wire n_1142;
wire GPR_19__3_;
wire n_4519;
wire n_2819;
wire n_346;
wire n_938;
wire SP_2_;
wire n_4664;
wire n_1412;
wire GPR_11__5_;
wire GPR_3__3_;
wire newNet_1079;
wire newNet_1021;
wire n_2057;
wire n_3227;
wire newNet_1749;
wire n_664;
wire n_479;
wire SP_4_;
wire n_1598;
wire newNet_745;
wire newNet_1791;
wire newNet_738;
wire n_2882;
wire n_160;
wire GPR_16__4_;
wire n_2985;
wire n_2135;
wire newNet_1540;
wire n_1978;
wire n_4062;
wire newNet_193;
wire newNet_684;
wire newNet_414;
wire n_2480;
wire newNet_1530;
wire R16_9_;
wire GPR_2__4_;
wire n_2285;
wire newNet_314;
wire newNet_1508;
wire n_616;
wire newNet_1137;
wire newNet_651;
wire n_3748;
wire newNet_1758;
wire n_1462;
wire newNet_318;
wire n_4261;
wire n_1591;
wire newNet_653;
wire n_1842;
wire n_2499;
wire n_584;
wire n_1867;
wire n_4595;
wire n_2707;
wire n_3991;
wire newNet_101;
wire n_640;
wire n_2755;
wire newNet_1269;
wire newNet_846;
wire newNet_1359;
wire n_305;
wire n_1077;
wire n_179;
wire newNet_113;
wire newNet_53;
wire newNet_1526;
wire GPR_2__2_;
wire n_977;
wire n_549;
wire n_1244;
wire n_1577;
wire n_2261;
wire n_1252;
wire newNet_611;
wire n_1849;
wire n_2945;
wire n_535;
wire newNet_1690;
wire n_772;
wire n_1554;
wire n_1919;
wire n_3380;
wire newNet_374;
wire newNet_1085;
wire n_4334;
wire n_2870;
wire n_3854;
wire n_789;
wire n_3907;
wire n_3191;
wire n_1803;
wire n_918;
wire n_2916;
wire n_2659;
wire n_4085;
wire newNet_157;
wire n_828;
wire n_3833;
wire n_391;
wire n_4413;
wire SP_0_;
wire newNet_1223;
wire newNet_618;
wire n_435;
wire n_4012;
wire pX_1_;
wire n_3056;
wire newNet_1115;
wire newNet_108;
wire newNet_150;
wire pX_13_;
wire n_3032;
wire n_2063;
wire n_6;
wire newNet_331;
wire n_974;
wire n_2638;
wire n_1201;
wire n_511;
wire n_2725;
wire n_3593;
wire newNet_1602;
wire n_3105;
wire n_2387;
wire n_37;
wire n_154;
wire n_4238;
wire pZ_6_;
wire GPR_6__3_;
wire newNet_1075;
wire PC_9_;
wire GPR_12__6_;
wire n_2032;
wire newNet_158;
wire GPR_Rd_r_5_;
wire n_653;
wire n_3970;
wire n_2210;
wire n_141;
wire newNet_400;
wire newNet_914;
wire n_361;
wire n_3901;
wire n_2006;
wire n_748;
wire n_3737;
wire n_1339;
wire n_4574;
wire n_2346;
wire n_2960;
wire n_3157;
wire newNet_116;
wire newNet_51;
wire n_853;
wire GPR_9__6_;
wire n_1748;
wire n_528;
wire n_2939;
wire n_2551;
wire n_637;
wire newNet_904;
wire n_360;
wire n_447;
wire n_2610;
wire n_4004;
wire n_3823;
wire n_2890;
wire newNet_23;
wire n_450;
wire n_234;
wire n_3214;
wire n_3914;
wire n_3099;
wire newNet_625;
wire GPR_10__4_;
wire n_2373;
wire newNet_624;
wire n_4531;
wire GPR_23__6_;
wire newNet_1547;
wire newNet_41;
wire n_1229;
wire n_1192;
wire n_3006;
wire n_644;
wire n_3575;
wire newNet_474;
wire n_52;
wire newNet_66;
wire final_adder_mux_R16_278_6_n_12;
wire newNet_207;
wire newNet_121;
wire newNet_1474;
wire n_3178;
wire n_1454;
wire newNet_1332;
wire final_adder_mux_R16_278_6_n_30;
wire n_3249;
wire n_2964;
wire n_2783;
wire n_3925;
wire n_4196;
wire newNet_635;
wire newNet_1607;
wire n_4172;
wire newNet_1536;
wire newNet_1229;
wire n_218;
wire newNet_1053;
wire newNet_392;
wire n_2236;
wire n_716;
wire n_3407;
wire newNet_1049;
wire n_3760;
wire n_4367;
wire n_2965;
wire n_3308;
wire newNet_137;
wire GPR_7__2_;
wire n_4118;
wire n_630;
wire n_2808;
wire n_731;
wire n_1270;
wire n_2977;
wire newNet_1329;
wire newNet_544;
wire n_2932;
wire n_4533;
wire newNet_204;
wire n_3665;
wire n_253;
wire newNet_461;
wire newNet_431;
wire newNet_1394;
wire n_3800;
wire n_1981;
wire newNet_94;
wire n_623;
wire n_3701;
wire pZ_11_;
wire newNet_1724;
wire newNet_1521;
wire n_1607;
wire newNet_1005;
wire n_3282;
wire newNet_1019;
wire n_381;
wire n_1507;
wire n_2608;
wire n_2087;
wire n_1996;
wire newNet_197;
wire newNet_959;
wire final_adder_mux_R16_278_6_n_6;
wire n_3751;
wire n_4635;
wire n_3933;
wire n_4524;
wire newNet_592;
wire n_3756;
wire n_2797;
wire newNet_1563;
wire newNet_581;
wire n_3013;
wire n_2319;
wire pmem_a_3;
wire n_2434;
wire newNet_439;
wire newNet_1584;
wire n_1238;
wire newNet_363;
wire n_4446;
wire n_4141;
wire n_1782;
wire newNet_1128;
wire n_2710;
wire n_3323;
wire newNet_1033;
wire n_2400;
wire n_2252;
wire newNet_1376;
wire n_39083_BAR;
wire n_167;
wire GPR_3__1_;
wire n_1032;
wire GPR_1__5_;
wire n_674;
wire n_1706;
wire newNet_1203;
wire n_369;
wire newNet_698;
wire n_982;
wire final_adder_mux_R16_278_6_n_43;
wire newNet_17;
wire n_3430;
wire n_1965;
wire n_1909;
wire n_691;
wire newNet_367;
wire n_1723;
wire newNet_1289;
wire n_1615;
wire n_3173;
wire n_2365;
wire n_3455;
wire n_4105;
wire n_2380;
wire n_2520;
wire newNet_1257;
wire n_2414;
wire newNet_596;
wire n_4271;
wire newNet_1471;
wire n_3508;
wire n_2538;
wire n_138;
wire io_di_4;
wire n_3054;
wire n_2507;
wire n_769;
wire GPR_17__7_;
wire n_1511;
wire newNet_1612;
wire n_1345;
wire n_2900;
wire n_1393;
wire newNet_1636;
wire n_3421;
wire pmem_d_12;
wire n_330;
wire n_1430;
wire n_2714;
wire n_2731;
wire newNet_239;
wire newNet_142;
wire newNet_354;
wire n_4348;
wire n_4480;
wire GPR_18__2_;
wire newNet_506;
wire n_3510;
wire n_3574;
wire n_211;
wire final_adder_mux_R16_278_6_n_68;
wire n_2248;
wire n_4354;
wire n_2549;
wire newNet_969;
wire n_3690;
wire n_460;
wire n_1373;
wire n_4126;
wire n_2427;
wire newNet_399;
wire n_521;
wire newNet_1752;
wire newNet_1489;
wire n_2016;
wire newNet_1282;
wire newNet_755;
wire n_3867;
wire n_209;
wire n_42;
wire newNet_1235;
wire n_1057;
wire GPR_Rd_r_6_;
wire n_1929;
wire newNet_1751;
wire n_2683;
wire newNet_1352;
wire n_4025;
wire n_4284;
wire n_1155;
wire GPR_20__3_;
wire n_4308;
wire n_1137;
wire n_342;
wire n_2081;
wire n_1760;
wire n_2527;
wire newNet_1026;
wire n_3963;
wire newNet_1818;
wire n_3976;
wire n_1429;
wire newNet_1798;
wire newNet_570;
wire n_3626;
wire newNet_254;
wire GPR_9__0_;
wire n_4326;
wire n_3807;
wire n_3318;
wire n_1860;
wire n_3764;
wire SP_9_;
wire n_4345;
wire n_1026;
wire final_adder_mux_R16_278_6_n_7;
wire n_206;
wire n_3424;
wire newNet_1702;
wire n_2770;
wire n_3583;
wire newNet_1833;
wire n_1836;
wire n_2738;
wire n_3779;
wire n_4466;
wire newNet_892;
wire n_540;
wire n_3691;
wire n_472;
wire n_3476;
wire U_12_;
wire n_1701;
wire n_1156;
wire n_1434;
wire n_2554;
wire n_1634;
wire dmem_do_2;
wire pmem_a_1;
wire GPR_4__6_;
wire n_725;
wire n_109;
wire pZ_10_;
wire newNet_1723;
wire n_2679;
wire newNet_786;
wire pmem_d_4;
wire n_2363;
wire newNet_871;
wire newNet_215;
wire final_adder_mux_R16_278_6_n_39;
wire n_3447;
wire n_1481;
wire n_762;
wire io_sp_3_;
wire newNet_273;
wire newNet_646;
wire newNet_605;
wire n_2536;
wire n_4301;
wire n_282;
wire n_3536;
wire n_340;
wire newNet_442;
wire newNet_1271;
wire newNet_305;
wire n_2660;
wire GPR_2__3_;
wire newNet_507;
wire n_4428;
wire n_3114;
wire n_415;
wire n_338;
wire n_3361;
wire n_604;
wire n_4212;
wire n_2910;
wire n_4272;
wire newNet_630;
wire n_3565;
wire n_4024;
wire n_4668;
wire final_adder_mux_R16_278_6_n_86;
wire newNet_1104;
wire n_4031;
wire n_4219;
wire newNet_1640;
wire newNet_1215;
wire n_570;
wire n_4156;
wire n_408;
wire n_698;
wire n_4682;
wire n_2037;
wire n_3269;
wire n_4606;
wire newNet_1402;
wire n_952;
wire n_3234;
wire n_228;
wire n_1293;
wire n_4661;
wire newNet_1416;
wire n_1025;
wire n_2699;
wire n_3770;
wire n_1286;
wire n_3200;
wire newNet_850;
wire n_3330;
wire newNet_808;
wire n_922;
wire n_2229;
wire io_a_1;
wire n_3230;
wire n_2205;
wire newNet_491;
wire n_4182;
wire n_1544;
wire n_819;
wire n_4226;
wire final_adder_mux_R16_278_6_n_83;
wire pZ_1_;
wire n_1625;
wire n_4435;
wire final_adder_mux_R16_278_6_n_18;
wire newNet_719;
wire n_4398;
wire n_3729;
wire n_4173;
wire newNet_1172;
wire n_4125;
wire newNet_1853;
wire n_22;
wire n_939;
wire n_177;
wire n_3444;
wire n_1788;
wire newNet_1627;
wire n_4142;
wire n_663;
wire newNet_1672;
wire newNet_569;
wire n_2351;
wire newNet_1421;
wire n_741;
wire n_2391;
wire n_420;
wire n_2521;
wire n_602;
wire n_704;
wire n_3716;
wire n_2957;
wire n_4564;
wire n_1497;
wire n_1043;
wire newNet_746;
wire pmem_d_13;
wire n_2466;
wire n_1874;
wire n_488;
wire newNet_1734;
wire n_4275;
wire n_2818;
wire newNet_638;
wire n_3356;
wire n_1630;
wire n_1127;
wire newNet_1770;
wire n_702;
wire n_1954;
wire n_463;
wire newNet_1056;
wire n_2573;
wire dmem_a_9;
wire newNet_1182;
wire n_4289;
wire SP_5_;
wire n_1409;
wire n_4241;
wire newNet_1461;
wire n_3743;
wire io_do_6;
wire newNet_1668;
wire newNet_265;
wire n_1344;
wire newNet_1313;
wire newNet_1499;
wire n_553;
wire newNet_838;
wire n_2861;
wire n_1530;
wire newNet_1305;
wire dmem_di_7;
wire newNet_1800;
wire GPR_18__0_;
wire newNet_1263;
wire n_2933;
wire newNet_486;
wire newNet_498;
wire n_1597;
wire newNet_981;
wire n_2146;
wire n_2613;
wire n_2078;
wire n_1623;
wire newNet_190;
wire n_596;
wire n_1162;
wire n_874;
wire n_1334;
wire n_4256;
wire n_711;
wire dmem_a_2;
wire newNet_997;
wire newNet_978;
wire n_3433;
wire newNet_409;
wire n_3010;
wire newNet_1353;
wire n_243;
wire n_2513;
wire newNet_1006;
wire n_3311;
wire n_1817;
wire n_401;
wire n_4137;
wire n_1608;
wire newNet_1453;
wire newNet_1165;
wire n_2796;
wire n_3333;
wire newNet_1828;
wire GPR_1__2_;
wire n_3025;
wire newNet_988;
wire n_1413;
wire newNet_115;
wire n_2452;
wire n_1568;
wire newNet_233;
wire n_1268;
wire newNet_496;
wire final_adder_mux_R16_278_6_n_21;
wire n_3657;
wire n_3394;
wire final_adder_mux_R16_278_6_n_26;
wire newNet_302;
wire n_790;
wire n_3633;
wire n_3611;
wire n_3228;
wire newNet_1149;
wire n_4418;
wire n_1125;
wire n_139;
wire n_583;
wire n_3035;
wire newNet_551;
wire n_3435;
wire newNet_1845;
wire newNet_993;
wire newNet_1844;
wire n_1796;
wire n_3080;
wire newNet_1595;
wire newNet_934;
wire newNet_795;
wire newNet_1406;
wire n_822;
wire n_1394;
wire n_2173;
wire n_3792;
wire GPR_1__0_;
wire n_1925;
wire newNet_85;
wire n_2164;
wire newNet_1389;
wire n_122;
wire newNet_560;
wire n_1231;
wire n_457;
wire newNet_1152;
wire n_1277;
wire n_4583;
wire newNet_510;
wire n_23;
wire n_3487;
wire n_3166;
wire n_3517;
wire Rd_r_2_;
wire n_2811;
wire n_2713;
wire n_2602;
wire newNet_182;
wire newNet_4;
wire newNet_32;
wire GPR_17__2_;
wire newNet_1192;
wire n_1539;
wire newNet_1157;
wire n_3820;
wire n_1092;
wire n_2763;
wire n_2559;
wire n_3945;
wire n_3073;
wire n_4338;
wire newNet_825;
wire n_4093;
wire newNet_1710;
wire n_2837;
wire n_1305;
wire n_62;
wire newNet_1661;
wire n_155;
wire newNet_1656;
wire n_510;
wire n_3879;
wire n_3096;
wire n_311;
wire n_965;
wire n_4644;
wire n_1321;
wire n_3207;
wire newNet_573;
wire n_1186;
wire n_687;
wire n_2552;
wire n_4299;
wire n_2335;
wire n_1224;
wire n_3125;
wire n_1799;
wire n_1941;
wire newNet_928;
wire GPR_22__6_;
wire n_2595;
wire n_30;
wire n_2102;
wire newNet_523;
wire n_4048;
wire n_4612;
wire n_2887;
wire n_943;
wire n_799;
wire n_3789;
wire n_3046;
wire newNet_664;
wire n_1508;
wire newNet_136;
wire n_532;
wire n_4187;
wire n_501;
wire newNet_168;
wire n_3468;
wire n_3347;
wire newNet_125;
wire n_112;
wire n_1189;
wire n_1821;
wire final_adder_mux_R16_278_6_n_75;
wire n_1365;
wire n_3260;
wire GPR_22__4_;
wire newNet_1047;
wire newNet_855;
wire n_2801;
wire n_3544;
wire n_4622;
wire n_2120;
wire n_882;
wire n_1315;
wire GPR_13__7_;
wire n_1472;
wire n_2998;
wire n_2325;
wire n_1524;
wire n_3252;
wire newNet_340;
wire n_3197;
wire n_4296;
wire n_2647;
wire n_3376;
wire n_3479;
wire n_4045;
wire n_3990;
wire n_1251;
wire n_3293;
wire n_956;
wire n_4572;
wire n_1664;
wire n_2299;
wire GPR_14__5_;
wire n_1309;
wire newNet_737;
wire n_4488;
wire n_2943;
wire n_2923;
wire n_3288;
wire n_1979;
wire newNet_1010;
wire n_3843;
wire GPR_3__2_;
wire n_60;
wire n_3529;
wire newNet_1279;
wire newNet_72;
wire n_2129;
wire n_1656;
wire newNet_1839;
wire n_186;
wire n_1444;
wire n_2464;
wire newNet_1680;
wire n_2893;
wire newNet_1094;
wire n_289;
wire n_4310;
wire n_2474;
wire n_2498;
wire newNet_1477;
wire n_4632;
wire n_1843;
wire n_2622;
wire n_893;
wire newNet_1491;
wire n_2568;
wire n_2286;
wire newNet_710;
wire newNet_224;
wire pZ_2_;
wire n_2832;
wire n_1051;
wire n_1522;
wire n_832;
wire newNet_1621;
wire n_1033;
wire newNet_1820;
wire n_384;
wire n_3470;
wire newNet_830;
wire n_1587;
wire n_67;
wire n_4384;
wire newNet_880;
wire n_3018;
wire n_3620;
wire n_999;
wire n_2223;
wire n_3829;
wire n_2857;
wire n_2476;
wire n_2153;
wire n_2426;
wire n_2291;
wire newNet_513;
wire GPR_21__5_;
wire n_845;
wire newNet_673;
wire newNet_328;
wire n_3599;
wire n_4140;
wire n_3182;
wire n_2590;
wire n_2154;
wire newNet_175;
wire newNet_532;
wire n_2436;
wire n_4361;
wire n_1243;
wire n_429;
wire n_3736;
wire n_467;
wire newNet_1784;
wire newNet_626;
wire n_1858;
wire n_2823;
wire n_1850;
wire newNet_1483;
wire newNet_426;
wire n_3680;
wire n_2917;
wire n_2098;
wire R16_13_;
wire n_4100;
wire newNet_1246;
wire n_2064;
wire newNet_905;
wire newNet_1436;
wire n_1138;
wire newNet_707;
wire n_4086;
wire n_1810;
wire newNet_120;
wire final_adder_mux_R16_278_6_n_69;
wire n_730;
wire newNet_1520;
wire n_2651;
wire n_2915;
wire newNet_130;
wire newNet_24;
wire n_2300;
wire n_1328;
wire n_4337;
wire n_210;
wire newNet_1076;
wire newNet_1086;
wire n_2270;
wire newNet_117;
wire newNet_63;
wire n_3075;
wire newNet_1601;
wire io_sel_1_;
wire n_362;
wire n_4487;
wire newNet_1677;
wire n_3654;
wire n_3822;
wire newNet_739;
wire n_2354;
wire newNet_1500;
wire n_341;
wire n_541;
wire newNet_593;
wire GPR_13__2_;
wire n_652;
wire n_451;
wire n_737;
wire newNet_1590;
wire n_4327;
wire n_749;
wire n_3098;
wire newNet_124;
wire newNet_149;
wire n_4307;
wire newNet_375;
wire n_2015;
wire pmem_d_6;
wire n_2807;
wire newNet_730;
wire n_3915;
wire n_3761;
wire n_1453;
wire n_534;
wire n_4333;
wire newNet_1261;
wire n_256;
wire newNet_1038;
wire newNet_460;
wire n_3179;
wire n_2963;
wire newNet_1537;
wire newNet_1397;
wire newNet_272;
wire n_2645;
wire newNet_1817;
wire n_3307;
wire Z;
wire n_1740;
wire n_92;
wire newNet_1554;
wire newNet_670;
wire n_2780;
wire n_233;
wire newNet_1703;
wire newNet_1331;
wire newNet_1290;
wire n_53;
wire n_3248;
wire n_1154;
wire n_107;
wire n_1781;
wire n_2193;
wire n_645;
wire newNet_1340;
wire newNet_1548;
wire n_2784;
wire n_3592;
wire n_1082;
wire n_797;
wire n_1387;
wire n_1202;
wire GPR_12__7_;
wire newNet_174;
wire newNet_1576;
wire n_2394;
wire newNet_1103;
wire n_3641;
wire dmem_do_5;
wire n_2765;
wire newNet_917;
wire newNet_891;
wire GPR_13__0_;
wire n_1729;
wire n_622;
wire n_3481;
wire pmem_d_5;
wire n_3199;
wire n_2031;
wire n_3404;
wire final_adder_mux_R16_278_6_n_31;
wire n_2309;
wire n_4076;
wire newNet_449;
wire n_1145;
wire newNet_1790;
wire n_3699;
wire n_290;
wire n_26;
wire n_641;
wire n_1895;
wire newNet_1541;
wire newNet_1358;
wire n_1635;
wire n_2869;
wire n_4596;
wire n_2409;
wire n_1918;
wire newNet_464;
wire n_1260;
wire n_4447;
wire n_2756;
wire n_1868;
wire pmem_a_0;
wire newNet_1733;
wire n_2988;
wire newNet_313;
wire n_1962;
wire n_773;
wire n_3946;
wire n_2600;
wire newNet_1193;
wire n_3316;
wire n_1999;
wire n_83;
wire newNet_645;
wire n_2269;
wire newNet_652;
wire newNet_317;
wire n_1210;
wire newNet_74;
wire n_4050;
wire newNet_877;
wire n_3698;
wire n_208;
wire newNet_610;
wire final_adder_mux_R16_278_6_n_62;
wire n_4260;
wire n_2433;
wire n_434;
wire n_4134;
wire newNet_654;
wire newNet_661;
wire n_1642;
wire T;
wire n_3584;
wire newNet_109;
wire newNet_255;
wire n_1804;
wire n_4433;
wire n_3832;
wire newNet_1226;
wire newNet_432;
wire R16_5_;
wire newNet_754;
wire n_2260;
wire n_2800;
wire n_1787;
wire newNet_50;
wire n_1209;
wire n_1812;
wire GPR_5__1_;
wire n_2326;
wire n_1722;
wire n_1299;
wire newNet_681;
wire n_1557;
wire n_847;
wire n_1253;
wire n_2110;
wire n_919;
wire pY_13_;
wire GPR_11__1_;
wire GPR_8__6_;
wire n_2888;
wire n_1667;
wire n_881;
wire n_266;
wire n_976;
wire n_2689;
wire newNet_1646;
wire newNet_631;
wire n_389;
wire U_10_;
wire n_4543;
wire newNet_1258;
wire n_936;
wire n_3373;
wire n_2218;
wire io_di_6;
wire final_adder_mux_R16_278_6_n_42;
wire n_3461;
wire n_3180;
wire R16_1_;
wire n_1739;
wire newNet_923;
wire n_3348;
wire n_2662;
wire newNet_872;
wire n_983;
wire n_1550;
wire n_1680;
wire n_2682;
wire n_4351;
wire n_3977;
wire newNet_280;
wire newNet_1320;
wire n_3156;
wire n_3767;
wire newNet_659;
wire newNet_398;
wire newNet_216;
wire n_393;
wire newNet_1154;
wire GPR_23__3_;
wire n_4412;
wire n_2817;
wire n_2553;
wire newNet_411;
wire n_3971;
wire n_742;
wire n_3271;
wire n_2047;
wire GPR_14__7_;
wire newNet_1517;
wire newNet_294;
wire n_140;
wire n_3213;
wire n_3057;
wire newNet_597;
wire n_1061;
wire n_529;
wire n_3573;
wire n_2385;
wire n_902;
wire n_1058;
wire n_4129;
wire n_2442;
wire n_1992;
wire n_1942;
wire n_1421;
wire GPR_18__4_;
wire n_1835;
wire n_3839;
wire newNet_937;
wire newNet_1657;
wire n_3190;
wire n_3742;
wire n_3561;
wire newNet_1743;
wire newNet_1351;
wire n_2388;
wire n_3900;
wire n_4393;
wire n_351;
wire newNet_720;
wire newNet_1529;
wire newNet_1759;
wire newNet_768;
wire n_2577;
wire n_2277;
wire R16_14_;
wire n_3425;
wire n_3869;
wire newNet_1127;
wire n_1028;
wire n_4375;
wire newNet_1054;
wire n_1903;
wire n_374;
wire newNet_910;
wire n_1191;
wire n_3317;
wire final_adder_mux_R16_278_6_n_20;
wire newNet_1722;
wire n_3310;
wire GPR_1__3_;
wire n_2376;
wire n_1433;
wire n_1928;
wire n_4195;
wire n_1563;
wire n_3922;
wire newNet_1365;
wire n_473;
wire newNet_1366;
wire n_4148;
wire n_1185;
wire n_3140;
wire n_1035;
wire newNet_729;
wire GPR_23__2_;
wire n_4340;
wire n_1414;
wire n_4239;
wire newNet_1753;
wire newNet_966;
wire n_4346;
wire n_3501;
wire pmem_a_2;
wire n_2528;
wire n_4163;
wire n_3446;
wire n_2798;
wire newNet_1386;
wire n_3206;
wire newNet_787;
wire n_4249;
wire n_2678;
wire newNet_1347;
wire newNet_956;
wire n_3017;
wire n_3507;
wire n_803;
wire newNet_1861;
wire n_110;
wire n_2730;
wire newNet_1377;
wire n_2253;
wire n_717;
wire n_382;
wire n_168;
wire n_996;
wire newNet_1472;
wire n_2995;
wire io_di_3;
wire newNet_1509;
wire newNet_1531;
wire newNet_1198;
wire n_1221;
wire GPR_Rd_r_4_;
wire newNet_580;
wire n_3951;
wire n_4473;
wire n_2609;
wire GPR_6__2_;
wire newNet_232;
wire newNet_1772;
wire n_888;
wire n_244;
wire n_191;
wire newNet_1840;
wire n_1705;
wire n_2140;
wire n_277;
wire n_3415;
wire n_3750;
wire n_1819;
wire newNet_1834;
wire n_4270;
wire newNet_301;
wire n_840;
wire n_1489;
wire n_2040;
wire n_306;
wire newNet_366;
wire U_14_;
wire newNet_1583;
wire n_3722;
wire newNet_484;
wire n_2402;
wire n_149;
wire final_adder_mux_R16_278_6_n_8;
wire n_1599;
wire n_4523;
wire n_2548;
wire n_3431;
wire n_1711;
wire n_1392;
wire n_1129;
wire n_2741;
wire newNet_1611;
wire pmem_a_9;
wire n_1749;
wire n_1889;
wire n_595;
wire n_788;
wire n_3759;
wire n_3055;
wire n_2126;
wire n_2581;
wire n_3550;
wire n_3625;
wire n_852;
wire n_1512;
wire n_3451;
wire n_2744;
wire pmem_d_11;
wire n_3522;
wire n_1424;
wire newNet_520;
wire n_3300;
wire n_2715;
wire n_1898;
wire n_839;
wire newNet_1145;
wire newNet_1604;
wire n_3484;
wire n_1237;
wire GPR_14__4_;
wire newNet_362;
wire newNet_1597;
wire n_3802;
wire newNet_156;
wire n_677;
wire n_4242;
wire n_1227;
wire newNet_697;
wire newNet_59;
wire n_4369;
wire n_756;
wire n_4068;
wire n_2696;
wire n_476;
wire n_1346;
wire n_3984;
wire n_3473;
wire n_3281;
wire n_1890;
wire n_768;
wire n_813;
wire newNet_1083;
wire n_4319;
wire newNet_1635;
wire n_1908;
wire n_1188;
wire newNet_1405;
wire newNet_1185;
wire newNet_992;
wire newNet_1330;
wire n_3604;
wire newNet_728;
wire newNet_238;
wire n_804;
wire n_4623;
wire n_1622;
wire newNet_1116;
wire final_adder_mux_R16_278_6_n_74;
wire newNet_191;
wire newNet_499;
wire n_2646;
wire newNet_1025;
wire newNet_361;
wire newNet_1681;
wire n_4255;
wire newNet_837;
wire n_4288;
wire newNet_711;
wire n_4482;
wire n_3853;
wire newNet_380;
wire n_1408;
wire newNet_477;
wire newNet_996;
wire newNet_472;
wire n_3060;
wire newNet_1314;
wire n_4404;
wire newNet_1173;
wire final_adder_mux_R16_278_6_n_41;
wire n_2976;
wire newNet_397;
wire GPR_Rd_r_3_;
wire GPR_16__0_;
wire n_2089;
wire n_3715;
wire newNet_355;
wire n_1761;
wire newNet_1060;
wire n_2301;
wire n_1645;
wire n_1163;
wire newNet_753;
wire GPR_9__2_;
wire n_1569;
wire n_802;
wire n_710;
wire newNet_911;
wire newNet_88;
wire n_3357;
wire n_3668;
wire newNet_1146;
wire n_3334;
wire n_1410;
wire n_3778;
wire newNet_1667;
wire n_667;
wire n_3279;
wire n_662;
wire n_4069;
wire n_2850;
wire newNet_796;
wire n_1269;
wire newNet_550;
wire n_3395;
wire pX_8_;
wire io_do_3;
wire n_2489;
wire n_3793;
wire n_4037;
wire n_2737;
wire n_3781;
wire GPR_12__3_;
wire n_1333;
wire newNet_773;
wire newNet_533;
wire n_3011;
wire GPR_1__6_;
wire n_2533;
wire newNet_1292;
wire n_4352;
wire newNet_982;
wire n_3828;
wire n_1609;
wire n_3688;
wire n_699;
wire n_2742;
wire newNet_1846;
wire n_1993;
wire n_2623;
wire n_2514;
wire n_1551;
wire newNet_1036;
wire n_3383;
wire n_3034;
wire n_2172;
wire newNet_1801;
wire n_3619;
wire newNet_1264;
wire newNet_497;
wire n_4607;
wire dmem_a_8;
wire newNet_1596;
wire newNet_487;
wire newNet_391;
wire GPR_23__4_;
wire n_1463;
wire n_1702;
wire n_3081;
wire dmem_a_1;
wire newNet_841;
wire n_462;
wire n_3679;
wire GPR_15__5_;
wire newNet_1401;
wire n_605;
wire GPR_6__1_;
wire n_562;
wire n_923;
wire n_1420;
wire newNet_441;
wire n_3676;
wire pX_3_;
wire n_1498;
wire n_3102;
wire n_2779;
wire n_2097;
wire newNet_1575;
wire n_2934;
wire n_3360;
wire n_4401;
wire newNet_1650;
wire n_1317;
wire n_889;
wire n_1525;
wire final_adder_mux_R16_278_6_n_48;
wire pX_12_;
wire newNet_1138;
wire n_4017;
wire newNet_1399;
wire newNet_1020;
wire n_4662;
wire n_1574;
wire n_1955;
wire n_2826;
wire n_2522;
wire n_414;
wire n_1600;
wire n_1128;
wire n_2661;
wire n_3090;
wire newNet_1742;
wire n_4213;
wire n_953;
wire n_1910;
wire newNet_810;
wire n_2441;
wire n_4517;
wire n_3231;
wire n_4434;
wire n_2726;
wire newNet_553;
wire n_3235;
wire n_409;
wire n_3077;
wire n_1624;
wire n_1592;
wire newNet_692;
wire n_866;
wire n_2578;
wire n_4029;
wire newNet_843;
wire newNet_386;
wire n_3978;
wire n_470;
wire pX_6_;
wire n_1818;
wire n_1631;
wire n_448;
wire GPR_17__6_;
wire newNet_248;
wire n_4164;
wire newNet_419;
wire newNet_970;
wire newNet_242;
wire n_421;
wire newNet_1424;
wire n_4174;
wire n_4049;
wire n_3809;
wire newNet_163;
wire n_38;
wire n_4395;
wire n_4225;
wire n_2101;
wire newNet_1628;
wire n_494;
wire n_433;
wire n_2574;
wire newNet_644;
wire n_3868;
wire n_2055;
wire n_3814;
wire newNet_1174;
wire n_3539;
wire n_2506;
wire n_603;
wire n_178;
wire n_3134;
wire n_586;
wire newNet_807;
wire n_4376;
wire pX_5_;
wire newNet_1232;
wire pZ_3_;
wire newNet_1514;
wire n_2333;
wire n_4657;
wire n_1242;
wire newNet_979;
wire n_4112;
wire newNet_760;
wire n_5;
wire n_875;
wire n_957;
wire n_2435;
wire newNet_71;
wire n_4133;
wire n_3460;
wire n_1455;
wire newNet_463;
wire newNet_401;
wire newNet_676;
wire n_487;
wire n_2862;
wire n_2465;
wire newNet_617;
wire n_2192;
wire n_3478;
wire newNet_1478;
wire n_1292;
wire n_2473;
wire newNet_225;
wire n_1829;
wire n_1657;
wire n_3261;
wire n_84;
wire GPR_7__4_;
wire n_892;
wire n_1261;
wire n_3240;
wire n_4300;
wire newNet_465;
wire n_1738;
wire n_1443;
wire n_899;
wire n_2560;
wire newNet_1468;
wire n_185;
wire n_3247;
wire newNet_457;
wire n_2070;
wire n_2419;
wire newNet_1093;
wire newNet_888;
wire n_113;
wire n_2668;
wire n_1844;
wire newNet_944;
wire n_571;
wire newNet_547;
wire n_153;
wire n_3287;
wire n_2206;
wire n_59;
wire n_2894;
wire newNet_1827;
wire newNet_1066;
wire n_128;
wire n_3229;
wire n_2152;
wire n_1052;
wire n_3183;
wire n_3842;
wire n_4087;
wire newNet_1384;
wire n_2224;
wire newNet_858;
wire dmem_di_0;
wire n_2463;
wire n_350;
wire n_229;
wire n_4383;
wire final_adder_mux_R16_278_6_n_78;
wire n_846;
wire n_3612;
wire n_1857;
wire newNet_1785;
wire newNet_606;
wire n_2292;
wire n_1353;
wire n_1811;
wire n_392;
wire n_1308;
wire newNet_102;
wire n_2944;
wire newNet_334;
wire n_3794;
wire n_1097;
wire newNet_1564;
wire n_2147;
wire n_3115;
wire newNet_1614;
wire n_3681;
wire n_910;
wire n_4362;
wire newNet_1620;
wire newNet_706;
wire n_3882;
wire n_2567;
wire newNet_538;
wire n_1059;
wire n_2111;
wire newNet_33;
wire n_3220;
wire newNet_1245;
wire GPR_19__5_;
wire newNet_291;
wire n_2858;
wire newNet_1153;
wire newNet_1435;
wire n_2247;
wire n_3777;
wire n_2025;
wire n_4357;
wire n_466;
wire newNet_425;
wire n_4092;
wire n_2475;
wire n_1314;
wire n_942;
wire Rd_r_0_;
wire n_1327;
wire n_3564;
wire n_4565;
wire newNet_1272;
wire n_3903;
wire n_1543;
wire n_2310;
wire n_684;
wire n_1538;
wire newNet_329;
wire n_281;
wire n_49;
wire n_4108;
wire n_2840;
wire pmem_a_10;
wire newNet_561;
wire n_2764;
wire n_4030;
wire n_2212;
wire n_2099;
wire newNet_60;
wire final_adder_mux_R16_278_6_n_54;
wire newNet_1415;
wire newNet_826;
wire newNet_716;
wire newNet_306;
wire n_4647;
wire n_106;
wire n_2838;
wire GPR_6__5_;
wire newNet_1396;
wire n_2163;
wire n_2603;
wire newNet_1660;
wire newNet_511;
wire newNet_64;
wire n_2411;
wire n_1276;
wire n_123;
wire n_3170;
wire GPR_23__1_;
wire n_3934;
wire newNet_860;
wire pZ_15_;
wire n_1728;
wire n_4649;
wire n_1364;
wire n_945;
wire n_3456;
wire newNet_1534;
wire n_3047;
wire n_2909;
wire n_1374;
wire newNet_865;
wire newNet_91;
wire n_31;
wire n_950;
wire newNet_332;
wire n_91;
wire n_1882;
wire n_72;
wire newNet_1238;
wire n_2336;
wire n_1509;
wire n_2121;
wire n_79;
wire n_4613;
wire n_1029;
wire n_1820;
wire n_903;
wire n_1693;
wire n_19;
wire n_1386;
wire n_1011;
wire n_1798;
wire n_2079;
wire n_1758;
wire n_2005;
wire newNet_194;
wire n_3889;
wire n_3072;
wire n_1672;
wire n_1003;
wire n_1164;
wire n_1304;
wire n_3642;
wire n_3545;
wire n_2946;
wire n_4188;
wire n_2584;
wire n_3872;
wire n_2343;
wire n_3196;
wire SP_11_;
wire n_4298;
wire newNet_1523;
wire n_1219;
wire n_1044;
wire n_4654;
wire newNet_1304;
wire n_1102;
wire n_1010;
wire n_798;
wire n_526;
wire pY_11_;
wire n_4007;
wire n_2920;
wire newNet_341;

// Start cells
NAND2_Z01 g59270 ( .a(n_1775), .b(n_464), .o(n_1853) );
BUF_X2 newInst_1154 ( .a(newNet_1153), .o(newNet_1154) );
NAND2_Z01 g59214 ( .a(n_1847), .b(n_267), .o(n_1903) );
BUF_X2 newInst_1859 ( .a(newNet_1858), .o(newNet_1859) );
BUF_X2 newInst_540 ( .a(newNet_539), .o(newNet_540) );
BUF_X2 newInst_224 ( .a(newNet_223), .o(newNet_224) );
NAND2_Z01 g61016 ( .a(n_121), .b(n_59), .o(n_166) );
BUF_X2 newInst_378 ( .a(newNet_115), .o(newNet_378) );
NOR3_Z1 g59034 ( .a(n_964), .b(n_1869), .c(n_963), .o(n_2084) );
BUF_X2 newInst_1472 ( .a(newNet_710), .o(newNet_1472) );
NAND3_Z1 g59198 ( .a(n_1644), .b(n_1834), .c(n_854), .o(n_1970) );
NAND2_Z01 g35209 ( .a(n_3321), .b(n_3296), .o(n_3451) );
BUF_X2 newInst_785 ( .a(newNet_784), .o(newNet_785) );
INV_X1 g35053 ( .a(n_3526), .o(Rd_4_) );
fflopd GPR_reg_20__7_ ( .CK(newNet_1170), .D(n_3156), .Q(GPR_20__7_) );
NAND4_Z2 g35186 ( .a(n_3389), .b(n_3406), .c(n_3401), .d(n_3398), .o(n_4644) );
NAND2_Z01 g59323 ( .a(n_1700), .b(n_4545), .o(n_1790) );
NAND4_Z1 g58980 ( .a(n_1015), .b(n_1881), .c(n_1889), .d(n_1759), .o(n_2127) );
NAND2_Z01 g58058 ( .a(n_2886), .b(n_2229), .o(n_2924) );
BUF_X2 newInst_1211 ( .a(newNet_1210), .o(newNet_1211) );
NOR2_Z1 g60603 ( .a(n_323), .b(n_189), .o(n_516) );
BUF_X2 newInst_1284 ( .a(newNet_1283), .o(newNet_1284) );
BUF_X2 newInst_369 ( .a(newNet_368), .o(newNet_369) );
NOR2_Z1 g60602 ( .a(n_334), .b(n_184), .o(n_517) );
BUF_X2 newInst_410 ( .a(newNet_409), .o(newNet_410) );
XOR2_X1 g58943 ( .a(n_2111), .b(n_288), .o(n_2164) );
NAND2_Z01 g60559 ( .a(n_392), .b(n_390), .o(n_547) );
BUF_X2 newInst_667 ( .a(newNet_547), .o(newNet_667) );
BUF_X2 newInst_1368 ( .a(newNet_1367), .o(newNet_1368) );
AND2_X1 g58511 ( .a(n_2567), .b(n_2205), .o(n_2585) );
NAND2_Z01 g57703 ( .a(n_3139), .b(n_2240), .o(n_3166) );
AND2_X1 g34511 ( .a(n_3994), .b(n_3995), .o(n_4034) );
NAND2_Z01 g58652 ( .a(n_2353), .b(n_1930), .o(n_2458) );
BUF_X2 newInst_1275 ( .a(newNet_1274), .o(newNet_1275) );
NAND2_Z02 g58913 ( .a(n_2160), .b(n_1172), .o(n_2209) );
BUF_X2 newInst_1107 ( .a(newNet_1106), .o(newNet_1107) );
BUF_X2 newInst_1048 ( .a(newNet_1047), .o(newNet_1048) );
BUF_X2 newInst_1821 ( .a(newNet_1820), .o(newNet_1821) );
BUF_X2 newInst_1168 ( .a(newNet_1167), .o(newNet_1168) );
AND2_X1 g60106 ( .a(n_839), .b(n_172), .o(n_1016) );
NAND4_Z1 g34089 ( .a(n_4256), .b(n_4237), .c(n_4343), .d(n_4143), .o(n_4388) );
NAND2_Z01 g58721 ( .a(n_2207), .b(GPR_22__2_), .o(n_2386) );
AND2_X1 g58359 ( .a(n_2657), .b(n_2139), .o(n_2712) );
NAND2_Z01 g58037 ( .a(n_2907), .b(n_2263), .o(n_2948) );
NAND2_Z01 g35221 ( .a(n_3354), .b(pmem_d_3), .o(n_3447) );
NAND2_Z01 g59504 ( .a(n_1556), .b(n_901), .o(n_1616) );
AND2_X1 g58405 ( .a(n_2657), .b(n_2199), .o(n_2663) );
AND2_X1 g57747 ( .a(n_3115), .b(n_2204), .o(n_3124) );
BUF_X2 newInst_693 ( .a(newNet_167), .o(newNet_693) );
NOR2_Z1 g60800 ( .a(n_177), .b(SP_13_), .o(n_314) );
AND2_X1 g58518 ( .a(n_2567), .b(n_2140), .o(n_2578) );
NAND2_Z01 g34803 ( .a(n_3582), .b(GPR_0__2_), .o(n_3760) );
NAND2_Z01 g58694 ( .a(n_2210), .b(GPR_1__1_), .o(n_2412) );
NAND2_Z01 g59352 ( .a(n_1731), .b(n_854), .o(n_1761) );
AND2_X1 g58368 ( .a(n_2656), .b(n_2156), .o(n_2703) );
BUF_X2 newInst_1465 ( .a(newNet_1464), .o(newNet_1465) );
BUF_X2 newInst_173 ( .a(newNet_172), .o(newNet_173) );
NAND2_Z01 g60503 ( .a(n_361), .b(GPR_5__6_), .o(n_643) );
NAND2_Z01 g60085 ( .a(n_786), .b(n_221), .o(n_1052) );
BUF_X2 newInst_108 ( .a(newNet_107), .o(newNet_108) );
XNOR2_X1 final_adder_mux_R16_278_6_g413 ( .a(n_4450), .b(n_4434), .o(final_adder_mux_R16_278_6_n_36) );
INV_X1 g61054 ( .a(SP_5_), .o(n_98) );
XOR2_X1 final_adder_mux_R16_278_6_g373 ( .a(final_adder_mux_R16_278_6_n_74), .b(final_adder_mux_R16_278_6_n_30), .o(R16_11_) );
AND2_X1 g58107 ( .a(n_2850), .b(n_2157), .o(n_2905) );
AND2_X1 g34351 ( .a(n_4178), .b(n_4042), .o(n_4183) );
NAND2_Z01 g34132 ( .a(n_4164), .b(GPR_Rd_r_2_), .o(n_4376) );
NOR2_Z1 g34375 ( .a(n_4125), .b(n_4072), .o(n_4166) );
NOR2_Z1 g59583 ( .a(n_1529), .b(n_4639), .o(n_1548) );
NAND2_Z01 g60726 ( .a(n_200), .b(GPR_12__4_), .o(n_412) );
NOR2_Z1 g34426 ( .a(n_4088), .b(n_3514), .o(n_4111) );
NAND4_Z1 g34586 ( .a(n_3748), .b(n_3651), .c(n_3677), .d(n_3747), .o(n_3974) );
BUF_X2 newInst_1474 ( .a(newNet_650), .o(newNet_1474) );
NAND2_Z01 g59058 ( .a(n_1902), .b(n_4596), .o(n_2049) );
INV_X1 g35514 ( .a(pY_4_), .o(n_3214) );
NAND2_Z01 g58769 ( .a(n_2202), .b(GPR_5__5_), .o(n_2331) );
NOR2_Z1 g35433 ( .a(n_3236), .b(pmem_d_3), .o(n_3287) );
NOR2_Z1 g59117 ( .a(n_1891), .b(n_87), .o(n_1992) );
BUF_X2 newInst_644 ( .a(newNet_643), .o(newNet_644) );
NAND2_Z01 g60236 ( .a(n_598), .b(GPR_15__0_), .o(n_909) );
NAND2_Z01 g58352 ( .a(n_2648), .b(n_2304), .o(n_2719) );
NAND2_Z01 g34937 ( .a(n_3543), .b(n_3294), .o(n_3638) );
NAND2_Z01 g58642 ( .a(n_2358), .b(pZ_3_), .o(n_2454) );
NAND2_Z01 g58536 ( .a(n_2529), .b(pY_15_), .o(n_2561) );
NAND2_Z01 g58899 ( .a(n_2158), .b(GPR_12__0_), .o(n_2183) );
NAND2_Z01 g60366 ( .a(n_486), .b(state_1_), .o(n_845) );
NAND2_Z01 g58051 ( .a(n_2894), .b(n_2376), .o(n_2931) );
NAND2_Z01 g34859 ( .a(n_3635), .b(GPR_14__0_), .o(n_3704) );
NAND2_Z01 g60552 ( .a(n_371), .b(GPR_21__6_), .o(n_554) );
NAND2_Z01 g59066 ( .a(n_1875), .b(n_4565), .o(n_2041) );
INV_X1 g35390 ( .a(n_3299), .o(n_3298) );
NAND2_Z01 g59460 ( .a(n_1614), .b(n_230), .o(n_1669) );
NOR4_Z1 g34478 ( .a(n_3460), .b(n_4657), .c(n_3963), .d(n_4664), .o(n_4064) );
NAND2_Z01 g58589 ( .a(n_2482), .b(n_1621), .o(n_2509) );
NAND2_Z01 g34506 ( .a(n_4646), .b(n_4645), .o(n_4039) );
INV_X1 g34370 ( .a(n_4613), .o(n_4162) );
XOR2_X1 g59733 ( .a(n_1306), .b(n_121), .o(n_1397) );
AND2_X1 g60810 ( .a(n_164), .b(SP_2_), .o(n_359) );
NAND2_Z01 g59646 ( .a(io_do_6), .b(n_1418), .o(n_1475) );
NAND4_Z1 g60134 ( .a(n_643), .b(n_554), .c(n_692), .d(n_537), .o(n_998) );
fflopd GPR_reg_21__2_ ( .CK(newNet_1150), .D(n_2762), .Q(GPR_21__2_) );
BUF_X2 newInst_1006 ( .a(newNet_1005), .o(newNet_1006) );
BUF_X2 newInst_20 ( .a(newNet_19), .o(newNet_20) );
NAND4_Z1 g57912 ( .a(n_1914), .b(n_2516), .c(n_2988), .d(n_2046), .o(n_3027) );
NAND2_Z01 g59079 ( .a(n_1871), .b(n_4605), .o(n_2028) );
BUF_X2 newInst_1166 ( .a(newNet_1165), .o(newNet_1166) );
BUF_X2 newInst_926 ( .a(newNet_925), .o(newNet_926) );
NAND2_Z01 g60499 ( .a(Rd_4_), .b(n_340), .o(n_647) );
NAND4_Z1 g58485 ( .a(n_297), .b(n_50), .c(n_2569), .d(n_239), .o(n_2611) );
NAND3_Z1 g34643 ( .a(n_3448), .b(n_3558), .c(n_3310), .o(n_3917) );
fflopd GPR_reg_17__6_ ( .CK(newNet_1380), .D(n_3083), .Q(GPR_17__6_) );
NOR3_Z1 g59300 ( .a(n_1704), .b(n_1358), .c(n_1311), .o(n_1827) );
XNOR2_X1 g59814 ( .a(n_1216), .b(pmem_d_2), .o(n_1343) );
NOR2_Z1 g60616 ( .a(n_459), .b(n_197), .o(n_591) );
NAND2_Z01 g58470 ( .a(n_2380), .b(n_2586), .o(n_2626) );
INV_X1 g60950 ( .a(n_198), .o(n_197) );
NOR2_Z1 g59018 ( .a(n_1974), .b(n_1919), .o(n_2091) );
NAND3_Z1 g58970 ( .a(n_262), .b(n_1938), .c(n_265), .o(n_2136) );
BUF_X2 newInst_1583 ( .a(newNet_1582), .o(newNet_1583) );
BUF_X2 newInst_1376 ( .a(newNet_1375), .o(newNet_1376) );
NAND2_Z01 g60915 ( .a(n_113), .b(pY_7_), .o(n_226) );
BUF_X2 newInst_700 ( .a(newNet_574), .o(newNet_700) );
NAND2_Z01 final_adder_mux_R16_278_6_g368 ( .a(final_adder_mux_R16_278_6_n_80), .b(final_adder_mux_R16_278_6_n_4), .o(final_adder_mux_R16_278_6_n_81) );
BUF_X2 newInst_647 ( .a(newNet_646), .o(newNet_647) );
NOR2_Z1 g58527 ( .a(n_2551), .b(n_579), .o(n_2570) );
NAND2_Z01 g57941 ( .a(n_2966), .b(n_2339), .o(n_3001) );
NAND2_Z01 g59830 ( .a(n_1217), .b(pX_7_), .o(n_1313) );
fflopd GPR_reg_22__6_ ( .CK(newNet_1074), .D(n_3074), .Q(GPR_22__6_) );
NAND2_Z01 g60574 ( .a(n_357), .b(pY_14_), .o(n_537) );
NAND2_Z01 g35111 ( .a(n_3457), .b(n_3290), .o(n_3495) );
INV_X1 g35109 ( .a(n_3490), .o(n_3489) );
BUF_X2 newInst_298 ( .a(newNet_297), .o(newNet_298) );
NAND2_Z01 g58632 ( .a(n_2354), .b(pX_2_), .o(n_2470) );
INV_X1 g61072 ( .a(pX_9_), .o(n_80) );
NOR2_Z1 g59728 ( .a(n_1355), .b(io_sel_1_), .o(n_1414) );
NOR2_Z1 g34275 ( .a(n_4163), .b(n_3238), .o(n_4258) );
NAND4_Z1 g58137 ( .a(n_2125), .b(n_2544), .c(n_2823), .d(n_2042), .o(n_2876) );
BUF_X2 newInst_1017 ( .a(newNet_1016), .o(newNet_1017) );
BUF_X2 newInst_10 ( .a(newNet_9), .o(newNet_10) );
NAND2_Z01 g60252 ( .a(n_605), .b(n_4686), .o(n_961) );
NAND2_Z01 g59684 ( .a(n_1317), .b(n_4665), .o(n_1441) );
NAND2_Z01 g58764 ( .a(n_2202), .b(GPR_5__0_), .o(n_2336) );
BUF_X2 newInst_216 ( .a(newNet_215), .o(newNet_216) );
BUF_X2 newInst_168 ( .a(newNet_167), .o(newNet_168) );
fflopd Z_reg ( .CK(newNet_348), .D(n_3193), .Q(Z) );
NOR2_Z1 g59359 ( .a(n_1701), .b(n_1631), .o(n_1754) );
NOR3_Z1 g58063 ( .a(n_1863), .b(n_2835), .c(n_1009), .o(n_2921) );
AND2_X1 g35241 ( .a(n_4487), .b(pmem_d_1), .o(n_4632) );
NOR2_Z1 g35212 ( .a(n_3364), .b(n_3338), .o(n_3438) );
BUF_X2 newInst_1243 ( .a(newNet_1242), .o(newNet_1243) );
NOR2_Z2 g60989 ( .a(pmem_d_9), .b(pmem_d_3), .o(n_183) );
NAND2_Z01 g35403 ( .a(pY_9_), .b(pY_8_), .o(n_3306) );
NAND2_Z01 g60223 ( .a(n_588), .b(GPR_7__3_), .o(n_922) );
NAND2_Z01 g34770 ( .a(n_3628), .b(GPR_19__4_), .o(n_3795) );
BUF_X2 newInst_19 ( .a(newNet_18), .o(newNet_19) );
NAND4_Z1 g59449 ( .a(n_1340), .b(n_1479), .c(n_1611), .d(n_772), .o(n_1673) );
NAND2_Z02 g58919 ( .a(n_2154), .b(n_1172), .o(n_2203) );
AND2_X1 g35236 ( .a(n_3347), .b(n_4684), .o(n_3431) );
XOR2_X1 g59497 ( .a(n_1531), .b(n_48), .o(n_1631) );
BUF_X2 newInst_488 ( .a(newNet_487), .o(newNet_488) );
NAND2_Z01 g59023 ( .a(n_1977), .b(n_1447), .o(n_2079) );
BUF_X2 newInst_197 ( .a(newNet_196), .o(newNet_197) );
NAND2_Z01 g60877 ( .a(pY_0_), .b(pY_1_), .o(n_280) );
NAND2_Z01 g57842 ( .a(n_3034), .b(n_2322), .o(n_3068) );
INV_X1 g61029 ( .a(pX_6_), .o(n_123) );
NAND2_Z01 g60679 ( .a(n_237), .b(n_268), .o(n_472) );
BUF_X2 newInst_340 ( .a(newNet_339), .o(newNet_340) );
NAND2_Z01 g60263 ( .a(n_584), .b(GPR_18__6_), .o(n_883) );
AND2_X1 g58370 ( .a(n_2657), .b(n_2214), .o(n_2701) );
NAND2_Z01 g35033 ( .a(n_3524), .b(n_3503), .o(n_3540) );
BUF_X2 newInst_1701 ( .a(newNet_1700), .o(newNet_1701) );
NAND2_Z01 g35080 ( .a(n_3495), .b(n_3268), .o(n_3505) );
BUF_X2 newInst_1290 ( .a(newNet_1289), .o(newNet_1290) );
NAND2_Z01 g59399 ( .a(n_1647), .b(n_1375), .o(n_1716) );
AND3_X1 g58066 ( .a(n_2552), .b(n_2893), .c(n_2673), .o(n_2919) );
fflopd U_reg_7_ ( .CK(newNet_365), .D(n_3183), .Q(U_7_) );
INV_X1 g34983 ( .a(n_3563), .o(n_3562) );
NAND2_Z01 g59745 ( .a(n_1314), .b(n_185), .o(n_1377) );
fflopd pX_reg_11_ ( .CK(newNet_272), .D(n_2952), .Q(pX_11_) );
NAND3_Z1 g59182 ( .a(N), .b(n_1827), .c(n_41), .o(n_1925) );
NAND2_Z01 g34260 ( .a(n_4176), .b(pX_3_), .o(n_4273) );
NAND2_Z01 g58774 ( .a(n_2201), .b(GPR_6__2_), .o(n_2326) );
NAND2_Z01 g57808 ( .a(n_3078), .b(n_1387), .o(n_3099) );
INV_X2 newInst_375 ( .a(newNet_374), .o(newNet_375) );
NOR2_Z1 g35061 ( .a(n_3507), .b(pX_7_), .o(n_4515) );
NAND2_Z01 g34706 ( .a(n_3629), .b(GPR_3__6_), .o(n_3859) );
BUF_X2 newInst_1671 ( .a(newNet_1670), .o(newNet_1671) );
NAND2_Z01 g60129 ( .a(n_780), .b(pmem_d_3), .o(n_1031) );
BUF_X2 newInst_42 ( .a(newNet_41), .o(newNet_42) );
BUF_X2 newInst_716 ( .a(newNet_715), .o(newNet_716) );
XOR2_X1 g58613 ( .a(n_2274), .b(pmem_d_9), .o(n_2485) );
BUF_X2 newInst_808 ( .a(newNet_807), .o(newNet_808) );
NAND2_Z01 g34887 ( .a(n_3564), .b(pX_1_), .o(n_3676) );
INV_X1 drc_bufs35587 ( .a(n_4684), .o(n_3200) );
BUF_X2 newInst_102 ( .a(newNet_101), .o(newNet_102) );
NAND2_Z01 g59392 ( .a(n_1648), .b(dmem_di_3), .o(n_1723) );
NAND2_Z01 g34950 ( .a(n_3549), .b(U_11_), .o(n_3612) );
NAND2_Z01 g34603 ( .a(n_3788), .b(n_3669), .o(n_3956) );
NAND2_Z02 g58910 ( .a(n_2161), .b(n_1203), .o(n_2212) );
INV_X1 g35230 ( .a(n_3424), .o(n_3425) );
NAND2_Z01 g57830 ( .a(n_3046), .b(n_2440), .o(n_3083) );
NAND2_Z01 g59940 ( .a(n_1109), .b(pmem_d_1), .o(n_1184) );
INV_Z1 g16807 ( .a(GPR_5__1_), .o(n_4402) );
NAND2_Z02 g58959 ( .a(n_2115), .b(n_1211), .o(n_2157) );
NOR2_Z1 g59297 ( .a(n_1773), .b(rst), .o(n_1828) );
NAND2_Z01 g34617 ( .a(n_3895), .b(n_3483), .o(n_3943) );
BUF_X2 newInst_1108 ( .a(newNet_1107), .o(newNet_1108) );
NOR2_Z1 g35254 ( .a(n_3315), .b(pZ_10_), .o(n_4519) );
BUF_X2 newInst_233 ( .a(newNet_232), .o(newNet_233) );
NAND2_X2 g58905 ( .a(n_2129), .b(n_2113), .o(n_2217) );
NAND2_Z01 g58590 ( .a(n_2461), .b(pX_3_), .o(n_2508) );
AND2_X1 g34249 ( .a(n_4188), .b(state_2_), .o(n_4284) );
INV_X1 g61083 ( .a(n_4615), .o(n_69) );
BUF_X2 newInst_1385 ( .a(newNet_961), .o(newNet_1385) );
NAND4_Z1 g59550 ( .a(n_1354), .b(n_1496), .c(n_1480), .d(n_496), .o(n_1578) );
NAND2_Z01 g35368 ( .a(n_4659), .b(n_3220), .o(n_3347) );
BUF_X2 newInst_530 ( .a(newNet_529), .o(newNet_530) );
BUF_X2 newInst_1219 ( .a(newNet_1218), .o(newNet_1219) );
NAND2_Z01 g59051 ( .a(n_18), .b(n_4572), .o(n_2056) );
NOR2_Z1 g35136 ( .a(n_4639), .b(n_4641), .o(io_re) );
NOR2_Z1 g35042 ( .a(n_3517), .b(n_4629), .o(n_3531) );
NAND2_Z01 g34348 ( .a(n_4161), .b(n_4574), .o(n_4186) );
BUF_X2 newInst_883 ( .a(newNet_882), .o(newNet_883) );
BUF_X2 newInst_1678 ( .a(newNet_660), .o(newNet_1678) );
XOR2_X1 g35015 ( .a(n_4517), .b(pY_8_), .o(n_4589) );
BUF_X2 newInst_241 ( .a(newNet_240), .o(newNet_241) );
BUF_X2 newInst_1798 ( .a(newNet_1797), .o(newNet_1798) );
BUF_X2 newInst_1564 ( .a(newNet_1563), .o(newNet_1564) );
BUF_X2 newInst_901 ( .a(newNet_338), .o(newNet_901) );
NAND2_Z01 g60548 ( .a(n_21), .b(Rd_r_1_), .o(n_558) );
NOR2_Z1 g34964 ( .a(n_3511), .b(n_3550), .o(n_3635) );
NAND2_Z01 g34960 ( .a(n_3536), .b(pY_4_), .o(n_3602) );
XOR2_X1 g59453 ( .a(n_1626), .b(n_106), .o(n_1670) );
NAND2_Z01 g34082 ( .a(n_4164), .b(GPR_Rd_r_1_), .o(n_4391) );
NAND2_Z01 g34544 ( .a(n_3916), .b(n_3920), .o(pmem_a_9) );
NAND2_Z01 g60924 ( .a(n_114), .b(pX_12_), .o(n_219) );
NAND2_Z01 g58783 ( .a(n_2200), .b(GPR_7__3_), .o(n_2317) );
BUF_X2 newInst_1633 ( .a(newNet_1632), .o(newNet_1633) );
XOR2_X1 g60831 ( .a(PC_5_), .b(pmem_d_8), .o(n_300) );
NAND2_Z01 g60696 ( .a(pY_1_), .b(n_249), .o(n_442) );
NAND2_Z01 g58466 ( .a(n_2413), .b(n_2591), .o(n_2630) );
fflopd GPR_reg_10__1_ ( .CK(newNet_1762), .D(n_2787), .Q(GPR_10__1_) );
NAND2_Z01 g59617 ( .a(n_1414), .b(io_di_3), .o(n_1510) );
AND2_X1 g58521 ( .a(n_2564), .b(n_587), .o(n_2576) );
NAND2_Z01 g58994 ( .a(n_2058), .b(n_4597), .o(n_2112) );
BUF_X2 newInst_1686 ( .a(newNet_1685), .o(newNet_1686) );
AND2_X1 g34193 ( .a(n_4324), .b(n_4626), .o(n_4330) );
NAND2_Z01 g58307 ( .a(n_2686), .b(n_2395), .o(n_2763) );
NAND2_Z01 g34833 ( .a(n_3568), .b(GPR_22__1_), .o(n_3730) );
fflopd GPR_reg_8__2_ ( .CK(newNet_723), .D(n_2737), .Q(GPR_8__2_) );
BUF_X2 newInst_23 ( .a(newNet_22), .o(newNet_23) );
NAND3_Z1 g34443 ( .a(n_3671), .b(n_4050), .c(n_3798), .o(n_4096) );
INV_X2 newInst_281 ( .a(newNet_280), .o(newNet_281) );
NAND3_Z1 g58130 ( .a(n_1233), .b(n_2790), .c(n_1076), .o(n_2883) );
BUF_X2 newInst_1278 ( .a(newNet_1277), .o(newNet_1278) );
NAND2_Z01 g60072 ( .a(n_841), .b(io_do_4), .o(n_1062) );
XNOR2_X1 g59047 ( .a(n_1903), .b(n_379), .o(n_2062) );
NAND3_Z1 g34551 ( .a(n_3833), .b(n_3835), .c(n_3834), .o(n_4008) );
BUF_X2 newInst_415 ( .a(newNet_414), .o(newNet_415) );
BUF_X2 newInst_1223 ( .a(newNet_1006), .o(newNet_1223) );
INV_X1 g35499 ( .a(pX_5_), .o(n_3228) );
NAND2_Z01 g59121 ( .a(n_1899), .b(n_1729), .o(n_1990) );
NAND2_Z01 g34737 ( .a(n_3625), .b(GPR_1__5_), .o(n_3828) );
NAND2_Z01 g34334 ( .a(n_4161), .b(n_4571), .o(n_4200) );
NOR2_Z1 g60809 ( .a(n_248), .b(n_182), .o(n_360) );
BUF_X2 newInst_1170 ( .a(newNet_1169), .o(newNet_1170) );
NAND2_Z01 g58479 ( .a(n_2578), .b(n_2223), .o(n_2615) );
AND2_X1 g59342 ( .a(n_381), .b(n_1695), .o(n_1775) );
NOR2_Z1 g58483 ( .a(n_2573), .b(n_579), .o(n_2613) );
NAND2_Z01 g34112 ( .a(n_4335), .b(n_4348), .o(n_4430) );
AND2_X1 g59575 ( .a(n_1466), .b(pmem_d_1), .o(n_1554) );
BUF_X2 newInst_1124 ( .a(newNet_1123), .o(newNet_1124) );
BUF_X2 newInst_1113 ( .a(newNet_1112), .o(newNet_1113) );
NAND2_Z01 g34319 ( .a(n_4166), .b(n_4549), .o(n_4214) );
BUF_X2 newInst_454 ( .a(newNet_453), .o(newNet_454) );
AND2_X1 g59279 ( .a(io_do_6), .b(n_1764), .o(n_1836) );
NOR2_Z1 g34995 ( .a(n_3510), .b(n_3553), .o(n_3587) );
BUF_X2 newInst_1063 ( .a(newNet_1062), .o(newNet_1063) );
XOR2_X1 final_adder_mux_R16_278_6_g391 ( .a(final_adder_mux_R16_278_6_n_56), .b(final_adder_mux_R16_278_6_n_40), .o(R16_5_) );
NAND2_Z01 g58797 ( .a(n_2195), .b(U_10_), .o(n_2303) );
BUF_X2 newInst_473 ( .a(newNet_472), .o(newNet_473) );
fflopd GPR_reg_0__4_ ( .CK(newNet_1790), .D(n_2922), .Q(GPR_0__4_) );
NAND2_Z01 g58845 ( .a(n_2139), .b(GPR_11__6_), .o(n_2262) );
NAND2_Z01 g60336 ( .a(n_566), .b(pmem_d_0), .o(n_794) );
fflopd GPR_reg_10__5_ ( .CK(newNet_1728), .D(n_3021), .Q(GPR_10__5_) );
NOR2_Z1 g34272 ( .a(n_4613), .b(n_3265), .o(n_4261) );
BUF_X2 newInst_1839 ( .a(newNet_1838), .o(newNet_1839) );
BUF_X2 newInst_248 ( .a(newNet_174), .o(newNet_248) );
XOR2_X1 g60393 ( .a(n_295), .b(n_266), .o(n_753) );
INV_X1 g59127 ( .a(n_1971), .o(n_1972) );
NAND2_Z01 g60412 ( .a(n_347), .b(GPR_11__4_), .o(n_734) );
fflopd GPR_reg_17__1_ ( .CK(newNet_1410), .D(n_2772), .Q(GPR_17__1_) );
NOR2_Z2 g35455 ( .a(pmem_d_5), .b(pmem_d_4), .o(n_3275) );
NAND2_Z01 g34792 ( .a(n_3599), .b(GPR_5__3_), .o(n_3773) );
NOR2_Z1 g59422 ( .a(io_do_7), .b(n_29), .o(n_1702) );
AND2_X1 g35123 ( .a(n_3466), .b(pZ_5_), .o(n_3488) );
NAND4_Z1 g59205 ( .a(n_1427), .b(n_1561), .c(n_1837), .d(n_1327), .o(n_1906) );
fflopd GPR_reg_4__1_ ( .CK(newNet_922), .D(n_2746), .Q(GPR_4__1_) );
NAND2_Z01 g35327 ( .a(pZ_2_), .b(n_3199), .o(n_3342) );
BUF_X2 newInst_908 ( .a(newNet_907), .o(newNet_908) );
fflopd GPR_reg_3__0_ ( .CK(newNet_977), .D(n_2624), .Q(GPR_3__0_) );
BUF_X2 newInst_874 ( .a(newNet_873), .o(newNet_874) );
BUF_X2 newInst_1 ( .a(newNet_0), .o(newNet_1) );
NOR2_Z1 g59718 ( .a(n_1343), .b(n_850), .o(n_1408) );
BUF_X2 newInst_1780 ( .a(newNet_1779), .o(newNet_1780) );
BUF_X2 newInst_443 ( .a(newNet_372), .o(newNet_443) );
NOR2_Z1 g60813 ( .a(n_250), .b(n_258), .o(n_357) );
BUF_X2 newInst_314 ( .a(newNet_313), .o(newNet_314) );
NAND2_Z01 g34779 ( .a(n_3571), .b(GPR_20__3_), .o(n_3786) );
NOR4_Z1 g34210 ( .a(n_3970), .b(n_3971), .c(n_4286), .d(n_3954), .o(n_4316) );
BUF_X2 newInst_1766 ( .a(newNet_1765), .o(newNet_1766) );
XNOR2_X1 g60862 ( .a(n_4450), .b(n_4434), .o(n_329) );
INV_X1 g35492 ( .a(pmem_d_12), .o(n_3233) );
BUF_X2 newInst_543 ( .a(newNet_542), .o(newNet_543) );
NAND2_Z01 g60424 ( .a(n_380), .b(GPR_4__2_), .o(n_722) );
NAND2_Z01 g60187 ( .a(n_663), .b(n_662), .o(n_966) );
XNOR2_X1 g60672 ( .a(n_279), .b(pX_2_), .o(n_477) );
NAND2_Z01 g57714 ( .a(n_3125), .b(n_2364), .o(n_3153) );
XOR2_X1 g34197 ( .a(n_4307), .b(SP_12_), .o(n_4326) );
BUF_X2 newInst_1694 ( .a(newNet_721), .o(newNet_1694) );
fflopd GPR_reg_6__4_ ( .CK(newNet_813), .D(n_2926), .Q(GPR_6__4_) );
NAND2_Z01 g58835 ( .a(n_2159), .b(GPR_10__1_), .o(n_2272) );
BUF_X2 newInst_1307 ( .a(newNet_1306), .o(newNet_1307) );
BUF_X2 newInst_881 ( .a(newNet_880), .o(newNet_881) );
BUF_X2 newInst_573 ( .a(newNet_572), .o(newNet_573) );
NAND2_Z01 g60979 ( .a(n_86), .b(n_52), .o(n_147) );
NAND2_Z01 g60443 ( .a(n_342), .b(GPR_19__1_), .o(n_703) );
AND2_X1 g59978 ( .a(n_4583), .b(n_1035), .o(n_1162) );
BUF_X2 newInst_1143 ( .a(newNet_1142), .o(newNet_1143) );
BUF_X2 newInst_828 ( .a(newNet_827), .o(newNet_828) );
NAND3_Z1 g59255 ( .a(n_1487), .b(n_1748), .c(n_303), .o(n_1857) );
NOR2_Z1 g34406 ( .a(n_4610), .b(n_3764), .o(n_4132) );
AND2_X1 g60104 ( .a(n_859), .b(io_do_5), .o(n_1048) );
NAND2_Z01 g59838 ( .a(n_1207), .b(n_1168), .o(n_1312) );
NOR2_Z1 g59169 ( .a(n_1893), .b(pY_14_), .o(n_1977) );
NAND2_Z01 g34854 ( .a(n_3568), .b(GPR_22__0_), .o(n_3709) );
XOR2_X1 g58413 ( .a(n_2641), .b(n_1769), .o(n_2687) );
AND2_X1 g59874 ( .a(n_1207), .b(n_473), .o(n_1253) );
BUF_X2 newInst_1496 ( .a(newNet_1495), .o(newNet_1496) );
AND2_X1 g59854 ( .a(n_1218), .b(rst), .o(n_1308) );
AND2_X1 g59365 ( .a(n_1698), .b(n_1269), .o(n_1748) );
INV_X2 newInst_1597 ( .a(newNet_27), .o(newNet_1597) );
NAND2_Z01 g60432 ( .a(n_353), .b(GPR_8__2_), .o(n_714) );
NOR4_Z1 g58986 ( .a(n_1725), .b(n_1758), .c(n_2000), .d(n_1013), .o(n_2121) );
BUF_X2 newInst_1134 ( .a(newNet_1133), .o(newNet_1134) );
BUF_X2 newInst_148 ( .a(newNet_147), .o(newNet_148) );
NAND2_Z01 g60706 ( .a(n_198), .b(GPR_17__4_), .o(n_432) );
NOR2_Z1 g59635 ( .a(n_1405), .b(n_1080), .o(n_1494) );
NOR2_Z1 g35359 ( .a(n_3297), .b(pmem_d_0), .o(n_3327) );
BUF_X2 newInst_398 ( .a(newNet_322), .o(newNet_398) );
BUF_X2 newInst_953 ( .a(newNet_952), .o(newNet_953) );
XOR2_X1 g59499 ( .a(n_1575), .b(n_83), .o(n_1629) );
NAND4_Z1 g59983 ( .a(n_512), .b(n_783), .c(n_757), .d(n_497), .o(n_1145) );
BUF_X2 newInst_940 ( .a(newNet_939), .o(newNet_940) );
NAND2_Z01 g59317 ( .a(n_4), .b(n_4537), .o(n_1796) );
NOR2_Z1 g34243 ( .a(n_4182), .b(n_4178), .o(n_4290) );
BUF_X2 newInst_1195 ( .a(newNet_1194), .o(newNet_1195) );
NAND2_Z01 g58744 ( .a(n_2204), .b(GPR_3__0_), .o(n_2363) );
BUF_X2 newInst_362 ( .a(newNet_300), .o(newNet_362) );
BUF_X2 newInst_133 ( .a(newNet_132), .o(newNet_133) );
INV_X1 g58314 ( .a(n_2752), .o(n_2751) );
BUF_X2 newInst_269 ( .a(newNet_268), .o(newNet_269) );
NAND2_Z01 g59561 ( .a(n_10), .b(n_594), .o(n_1565) );
fflopd pY_reg_4_ ( .CK(newNet_148), .D(n_3027), .Q(pY_4_) );
NOR3_Z1 g35096 ( .a(n_3433), .b(n_3465), .c(n_3455), .o(n_3497) );
AND2_X1 g57732 ( .a(n_3115), .b(n_2158), .o(n_3140) );
fflopd GPR_reg_14__1_ ( .CK(newNet_1572), .D(n_2779), .Q(GPR_14__1_) );
NAND2_Z01 g34098 ( .a(n_4367), .b(n_4366), .o(n_4440) );
NAND2_Z01 g57923 ( .a(n_2986), .b(n_2294), .o(n_3022) );
NAND2_Z01 g57931 ( .a(n_2976), .b(n_2441), .o(n_3014) );
NAND2_Z01 g35420 ( .a(n_3262), .b(state_0_), .o(n_4561) );
BUF_X2 newInst_190 ( .a(newNet_189), .o(newNet_190) );
BUF_X2 newInst_94 ( .a(newNet_93), .o(newNet_94) );
NAND2_Z01 g58039 ( .a(n_2905), .b(n_2184), .o(n_2946) );
NOR2_Z1 g59769 ( .a(n_1310), .b(rst), .o(n_1384) );
NOR2_Z1 g59651 ( .a(n_1451), .b(n_314), .o(n_1487) );
INV_X1 g59960 ( .a(n_1170), .o(n_1169) );
INV_X1 g34633 ( .a(n_4564), .o(n_3927) );
NOR2_Z1 g34325 ( .a(n_4612), .b(n_3477), .o(n_4209) );
NAND2_Z01 g59967 ( .a(n_984), .b(n_340), .o(n_1171) );
INV_X1 drc_bufs35524 ( .a(n_4616), .o(n_3206) );
BUF_X2 newInst_1805 ( .a(newNet_1804), .o(newNet_1805) );
fflopd SP_reg_12_ ( .CK(newNet_549), .D(n_1859), .Q(SP_12_) );
NAND2_Z01 g34711 ( .a(n_3625), .b(GPR_1__6_), .o(n_3854) );
NAND2_Z01 g58847 ( .a(n_2139), .b(GPR_11__7_), .o(n_2260) );
BUF_X2 newInst_1570 ( .a(newNet_1569), .o(newNet_1570) );
BUF_X2 newInst_1024 ( .a(newNet_1023), .o(newNet_1024) );
NAND2_Z01 g34828 ( .a(n_3575), .b(GPR_8__1_), .o(n_3735) );
BUF_X2 newInst_1235 ( .a(newNet_1234), .o(newNet_1235) );
NAND2_Z01 g59082 ( .a(n_1875), .b(n_4567), .o(n_2025) );
NOR2_Z1 g60638 ( .a(n_462), .b(n_250), .o(n_577) );
BUF_X2 newInst_1085 ( .a(newNet_1084), .o(newNet_1085) );
BUF_X2 newInst_1735 ( .a(newNet_1734), .o(newNet_1735) );
AND2_X1 g61010 ( .a(PC_0_), .b(PC_1_), .o(n_171) );
NOR2_Z1 g59862 ( .a(n_1219), .b(n_378), .o(n_1264) );
NAND2_Z01 g59338 ( .a(io_do_3), .b(n_1696), .o(n_1778) );
NOR2_Z1 g34880 ( .a(n_3565), .b(n_3229), .o(n_3683) );
NAND2_Z01 g60508 ( .a(n_380), .b(GPR_4__7_), .o(n_638) );
NAND4_Z1 g59668 ( .a(n_1065), .b(n_1289), .c(n_1366), .d(n_1060), .o(n_1460) );
INV_X2 newInst_422 ( .a(newNet_421), .o(newNet_422) );
NAND2_Z01 g34944 ( .a(n_3536), .b(GPR_20__2_), .o(n_3618) );
AND2_X1 g60077 ( .a(n_848), .b(n_44), .o(n_1058) );
BUF_X2 newInst_1627 ( .a(newNet_1626), .o(newNet_1627) );
BUF_X1 mybuffer0 ( .o(io_a_0), .a(pmem_d_0) );
NAND4_Z1 g58656 ( .a(n_1503), .b(n_1808), .c(n_2180), .d(n_1502), .o(n_2446) );
fflopd GPR_reg_19__1_ ( .CK(newNet_1317), .D(n_2769), .Q(GPR_19__1_) );
fflopd PC_reg_2_ ( .CK(newNet_640), .D(n_2278), .Q(PC_2_) );
BUF_X2 newInst_1528 ( .a(newNet_1527), .o(newNet_1528) );
BUF_X2 newInst_1515 ( .a(newNet_945), .o(newNet_1515) );
BUF_X2 newInst_1744 ( .a(newNet_1743), .o(newNet_1744) );
XOR2_X1 g60387 ( .a(n_468), .b(pY_3_), .o(n_759) );
NAND2_Z01 g35280 ( .a(pZ_15_), .b(n_3199), .o(n_3395) );
BUF_X2 newInst_534 ( .a(newNet_533), .o(newNet_534) );
NOR3_Z1 g60668 ( .a(n_4560), .b(n_130), .c(state_2_), .o(n_564) );
BUF_X2 newInst_227 ( .a(newNet_226), .o(newNet_227) );
NAND2_Z01 g35445 ( .a(n_3212), .b(n_3254), .o(n_3282) );
BUF_X2 newInst_1523 ( .a(newNet_1522), .o(newNet_1523) );
NAND2_Z01 g59924 ( .a(n_1120), .b(n_147), .o(n_1193) );
AND2_X1 g58502 ( .a(n_2567), .b(n_2214), .o(n_2595) );
NAND2_Z01 g60842 ( .a(n_128), .b(state_1_), .o(n_340) );
INV_Z1 g16795 ( .a(n_4464), .o(n_4411) );
INV_X1 g35515 ( .a(pmem_d_15), .o(n_3213) );
NAND2_Z01 g59510 ( .a(n_1562), .b(n_207), .o(n_1627) );
NAND2_Z01 g59398 ( .a(n_1647), .b(n_1189), .o(n_1717) );
BUF_X2 newInst_160 ( .a(newNet_159), .o(newNet_160) );
NOR2_Z1 g59106 ( .a(n_1901), .b(n_77), .o(n_2003) );
AND2_X1 g58116 ( .a(n_2850), .b(n_2208), .o(n_2896) );
NAND2_Z01 g34141 ( .a(n_4325), .b(n_4623), .o(n_4367) );
NAND3_Z1 g59799 ( .a(n_93), .b(n_1201), .c(SP_13_), .o(n_1327) );
NAND2_Z01 g35421 ( .a(pmem_d_3), .b(pmem_d_2), .o(n_3297) );
NAND2_Z01 g60423 ( .a(n_374), .b(GPR_12__3_), .o(n_723) );
BUF_X2 newInst_1194 ( .a(newNet_1193), .o(newNet_1194) );
BUF_X2 newInst_740 ( .a(newNet_29), .o(newNet_740) );
NAND2_Z01 g59160 ( .a(n_55), .b(n_1877), .o(n_1940) );
AND2_X1 g35219 ( .a(n_3413), .b(n_3252), .o(n_4530) );
AND4_X1 g60149 ( .a(n_4662), .b(n_4661), .c(n_4556), .d(n_296), .o(n_984) );
XOR2_X1 final_adder_mux_R16_278_6_g388 ( .a(final_adder_mux_R16_278_6_n_59), .b(final_adder_mux_R16_278_6_n_41), .o(R16_6_) );
NAND4_Z1 g60004 ( .a(n_831), .b(n_923), .c(n_878), .d(n_887), .o(n_1125) );
NAND2_Z01 g58291 ( .a(n_2705), .b(n_2236), .o(n_2779) );
NAND4_Z1 g60153 ( .a(n_670), .b(n_744), .c(n_650), .d(n_728), .o(n_982) );
NAND2_Z01 g35275 ( .a(U_5_), .b(n_3275), .o(n_3400) );
BUF_X2 newInst_710 ( .a(newNet_709), .o(newNet_710) );
NAND4_Z1 g34073 ( .a(n_4227), .b(n_4267), .c(n_4389), .d(n_4134), .o(dmem_a_8) );
AND2_X1 g58264 ( .a(n_2752), .b(n_2206), .o(n_2803) );
AND2_X1 g34405 ( .a(n_4089), .b(n_4635), .o(n_4133) );
NAND2_Z01 g34728 ( .a(n_3628), .b(GPR_18__5_), .o(n_3837) );
NAND2_Z01 g58242 ( .a(n_2755), .b(n_2216), .o(n_2825) );
AND2_X1 final_adder_mux_R16_278_6_g436 ( .a(n_4446), .b(n_4430), .o(final_adder_mux_R16_278_6_n_13) );
NAND2_Z01 g58622 ( .a(n_2358), .b(pZ_1_), .o(n_2475) );
NAND2_Z01 g60878 ( .a(io_do_2), .b(n_4652), .o(n_246) );
NAND2_Z01 g60584 ( .a(io_do_7), .b(n_22), .o(n_528) );
NAND2_Z01 g59402 ( .a(n_1223), .b(n_1650), .o(n_1714) );
NAND2_Z01 g34812 ( .a(n_3637), .b(n_3270), .o(n_3751) );
NAND4_Z1 g60148 ( .a(n_542), .b(n_559), .c(n_624), .d(n_722), .o(n_985) );
NAND2_Z01 g58321 ( .a(n_2674), .b(n_2335), .o(n_2744) );
XOR2_X1 g35077 ( .a(n_3494), .b(n_3323), .o(n_3514) );
fflopd GPR_Rd_r_reg_1_ ( .CK(newNet_1862), .D(io_do_1), .Q(GPR_Rd_r_1_) );
XOR2_X1 g59903 ( .a(n_1120), .b(n_319), .o(n_1227) );
NAND3_Z1 g58358 ( .a(n_218), .b(n_2612), .c(n_119), .o(n_2713) );
BUF_X2 newInst_1418 ( .a(newNet_663), .o(newNet_1418) );
XOR2_X1 g34252 ( .a(n_4172), .b(SP_6_), .o(n_4281) );
AND2_X1 g60827 ( .a(n_162), .b(io_do_2), .o(n_348) );
NAND2_Z01 g60492 ( .a(n_360), .b(GPR_1__7_), .o(n_654) );
AND2_X1 g58380 ( .a(n_2656), .b(n_2209), .o(n_2691) );
NAND2_Z01 g35305 ( .a(n_3289), .b(pY_3_), .o(n_3371) );
BUF_X2 newInst_706 ( .a(newNet_705), .o(newNet_706) );
AND2_X1 g58542 ( .a(n_2528), .b(n_587), .o(n_2556) );
BUF_X2 newInst_270 ( .a(newNet_269), .o(newNet_270) );
NAND2_Z01 g35329 ( .a(pZ_3_), .b(n_3199), .o(n_3340) );
NAND2_Z01 g34152 ( .a(n_4325), .b(n_4626), .o(n_4356) );
fflopd GPR_reg_16__6_ ( .CK(newNet_1433), .D(n_3084), .Q(GPR_16__6_) );
BUF_X2 newInst_766 ( .a(newNet_733), .o(newNet_766) );
BUF_X2 newInst_550 ( .a(newNet_525), .o(newNet_550) );
NAND3_Z1 g58339 ( .a(n_2457), .b(n_2654), .c(n_2110), .o(n_2730) );
NOR4_Z1 g34216 ( .a(n_4187), .b(n_4189), .c(n_4260), .d(n_4106), .o(n_4310) );
fflopd Rd_r_reg_4_ ( .CK(newNet_575), .D(n_951), .Q(Rd_r_4_) );
NAND4_Z1 g59540 ( .a(n_1301), .b(n_1511), .c(n_1510), .d(n_1074), .o(n_1588) );
BUF_X2 newInst_742 ( .a(newNet_741), .o(newNet_742) );
XOR2_X1 g60871 ( .a(n_4438), .b(n_4422), .o(n_322) );
NOR4_Z1 g34242 ( .a(n_4020), .b(n_4032), .c(n_4168), .d(n_3808), .o(n_4291) );
NAND2_Z01 g60750 ( .a(n_203), .b(SP_0_), .o(n_392) );
BUF_X2 newInst_896 ( .a(newNet_895), .o(newNet_896) );
NOR2_Z1 g59863 ( .a(n_1165), .b(io_do_3), .o(n_1263) );
INV_Z1 g16800 ( .a(n_4555), .o(n_4417) );
NAND2_Z01 g60562 ( .a(n_299), .b(n_228), .o(n_617) );
NAND2_Z01 g59177 ( .a(n_1872), .b(n_1390), .o(n_1930) );
NAND2_Z01 g60317 ( .a(n_600), .b(pX_7_), .o(n_809) );
INV_X1 g34439 ( .a(n_4099), .o(n_4100) );
NAND3_Z1 g57647 ( .a(n_1845), .b(n_3182), .c(n_1435), .o(n_3193) );
BUF_X2 newInst_1053 ( .a(newNet_1052), .o(newNet_1053) );
BUF_X2 newInst_501 ( .a(newNet_500), .o(newNet_501) );
NAND2_Z01 g60525 ( .a(n_374), .b(GPR_14__4_), .o(n_621) );
AND2_X1 g57998 ( .a(n_2940), .b(n_2210), .o(n_2973) );
XOR2_X1 g35380 ( .a(pZ_0_), .b(pmem_d_0), .o(n_3313) );
BUF_X2 newInst_1514 ( .a(newNet_1513), .o(newNet_1514) );
NOR2_Z1 g60207 ( .a(n_730), .b(n_4413), .o(n_938) );
NAND2_Z01 g57985 ( .a(n_2942), .b(n_2196), .o(n_2987) );
NAND2_Z01 g58302 ( .a(n_2696), .b(n_2420), .o(n_2768) );
BUF_X2 newInst_758 ( .a(newNet_757), .o(newNet_758) );
NAND2_Z01 g60881 ( .a(n_4616), .b(pmem_d_7), .o(n_244) );
BUF_X2 newInst_421 ( .a(newNet_420), .o(newNet_421) );
AND2_X1 g58271 ( .a(n_2752), .b(n_2153), .o(n_2796) );
NAND2_Z01 g34704 ( .a(n_3573), .b(U_6_), .o(n_3861) );
NOR2_Z1 g60114 ( .a(n_862), .b(rst), .o(n_1012) );
NAND4_Z1 g34566 ( .a(n_3861), .b(n_3863), .c(n_3864), .d(n_3664), .o(n_3994) );
AND2_X1 g58390 ( .a(n_2657), .b(n_2204), .o(n_2678) );
BUF_X2 newInst_131 ( .a(newNet_130), .o(newNet_131) );
NAND2_Z01 g59919 ( .a(n_1021), .b(n_245), .o(n_1221) );
NAND3_Z1 g60120 ( .a(n_4531), .b(n_857), .c(n_81), .o(n_1007) );
BUF_X2 newInst_755 ( .a(newNet_754), .o(newNet_755) );
AND2_X1 g59792 ( .a(n_1267), .b(pmem_d_7), .o(n_1332) );
NAND3_Z1 g59529 ( .a(n_1387), .b(n_1485), .c(H), .o(n_1598) );
AND2_X1 g58384 ( .a(n_2657), .b(n_2207), .o(n_2684) );
NAND2_Z01 g34487 ( .a(n_4036), .b(n_4561), .o(n_4054) );
INV_X1 g61102 ( .a(n_4657), .o(n_50) );
NOR2_Z1 g59884 ( .a(n_1191), .b(n_1196), .o(n_1243) );
INV_X1 g59236 ( .a(n_1871), .o(n_1870) );
fflopd PC_reg_7_ ( .CK(newNet_609), .D(n_2282), .Q(PC_7_) );
INV_X1 g61041 ( .a(pZ_6_), .o(n_111) );
NOR4_Z1 g34126 ( .a(n_4217), .b(n_4252), .c(n_4305), .d(n_4117), .o(n_4381) );
NAND2_Z01 g58559 ( .a(n_2505), .b(pZ_14_), .o(n_2539) );
BUF_X2 newInst_1757 ( .a(newNet_1756), .o(newNet_1757) );
BUF_X2 newInst_1741 ( .a(newNet_1740), .o(newNet_1741) );
NAND2_Z01 g34759 ( .a(n_3581), .b(GPR_16__4_), .o(n_3806) );
NOR2_Z1 g60028 ( .a(n_938), .b(n_4473), .o(n_1101) );
NAND4_Z1 g34583 ( .a(n_3693), .b(n_3774), .c(n_3773), .d(n_3772), .o(n_3977) );
NAND2_Z01 g60683 ( .a(n_200), .b(GPR_9__5_), .o(n_454) );
AND2_X1 g60593 ( .a(n_333), .b(n_254), .o(n_522) );
NAND2_Z01 g35261 ( .a(U_13_), .b(n_3275), .o(n_3411) );
AND2_X1 g59636 ( .a(n_1417), .b(n_90), .o(n_1493) );
AND2_X1 g34411 ( .a(n_4079), .b(n_4088), .o(n_4127) );
BUF_X2 newInst_1092 ( .a(newNet_1091), .o(newNet_1092) );
BUF_X2 newInst_937 ( .a(newNet_289), .o(newNet_937) );
BUF_X2 newInst_565 ( .a(newNet_564), .o(newNet_565) );
INV_X1 drc_bufs35539 ( .a(n_3201), .o(n_3198) );
BUF_X2 newInst_934 ( .a(newNet_933), .o(newNet_934) );
BUF_X2 newInst_601 ( .a(newNet_44), .o(newNet_601) );
AND3_X1 g59655 ( .a(n_80), .b(n_1390), .c(n_100), .o(n_1486) );
NOR2_Z1 g34472 ( .a(n_3207), .b(n_4039), .o(n_4070) );
NAND2_Z01 g60549 ( .a(n_358), .b(GPR_0__5_), .o(n_557) );
XNOR2_X1 g59452 ( .a(n_1627), .b(pmem_d_9), .o(n_1694) );
NAND2_Z01 g58096 ( .a(n_2851), .b(n_2218), .o(n_2917) );
NAND2_Z01 g60258 ( .a(n_585), .b(GPR_23__0_), .o(n_888) );
NAND2_Z01 g57837 ( .a(n_3039), .b(n_2373), .o(n_3073) );
INV_X1 drc_bufs35590 ( .a(n_3209), .o(n_4643) );
NAND2_Z01 g59559 ( .a(n_1527), .b(SP_2_), .o(n_1567) );
XOR2_X1 final_adder_mux_R16_278_6_g382 ( .a(final_adder_mux_R16_278_6_n_65), .b(final_adder_mux_R16_278_6_n_43), .o(R16_8_) );
INV_X1 g60948 ( .a(n_202), .o(n_201) );
NAND4_Z1 g59157 ( .a(n_4621), .b(n_4619), .c(n_1776), .d(n_4623), .o(n_1943) );
BUF_X2 newInst_438 ( .a(newNet_437), .o(newNet_438) );
BUF_X2 newInst_875 ( .a(newNet_874), .o(newNet_875) );
BUF_X2 newInst_110 ( .a(newNet_109), .o(newNet_110) );
NAND2_Z01 g60239 ( .a(n_591), .b(GPR_22__3_), .o(n_906) );
fflopd PC_reg_6_ ( .CK(newNet_617), .D(n_2), .Q(PC_6_) );
BUF_X2 newInst_1064 ( .a(newNet_405), .o(newNet_1064) );
AND2_X1 g58824 ( .a(n_2163), .b(n_587), .o(n_2281) );
BUF_X2 newInst_685 ( .a(newNet_684), .o(newNet_685) );
NAND2_Z01 g58552 ( .a(n_2495), .b(pY_11_), .o(n_2545) );
BUF_X2 newInst_86 ( .a(newNet_85), .o(newNet_86) );
BUF_X2 newInst_1555 ( .a(newNet_1554), .o(newNet_1555) );
BUF_X2 newInst_1455 ( .a(newNet_1454), .o(newNet_1455) );
BUF_X2 newInst_117 ( .a(newNet_116), .o(newNet_117) );
NOR2_Z2 g35029 ( .a(n_3467), .b(Rd_4_), .o(n_3551) );
BUF_X2 newInst_1408 ( .a(newNet_1407), .o(newNet_1408) );
NAND2_Z01 g58665 ( .a(n_2213), .b(GPR_17__5_), .o(n_2441) );
fflopd GPR_reg_13__0_ ( .CK(newNet_1613), .D(n_2636), .Q(GPR_13__0_) );
BUF_X2 newInst_591 ( .a(newNet_590), .o(newNet_591) );
fflopd GPR_reg_10__2_ ( .CK(newNet_1751), .D(n_2786), .Q(GPR_10__2_) );
BUF_X2 newInst_1264 ( .a(newNet_1263), .o(newNet_1264) );
BUF_X2 newInst_866 ( .a(newNet_865), .o(newNet_866) );
NOR2_Z1 g35169 ( .a(n_3428), .b(pX_4_), .o(n_3463) );
NAND3_Z1 g59531 ( .a(n_1336), .b(n_1572), .c(n_427), .o(n_1596) );
BUF_X2 newInst_1149 ( .a(newNet_1148), .o(newNet_1149) );
BUF_X2 newInst_1488 ( .a(newNet_1487), .o(newNet_1488) );
NAND2_Z01 g58549 ( .a(n_2521), .b(pZ_10_), .o(n_2548) );
NOR2_Z1 g35332 ( .a(n_3306), .b(n_3222), .o(n_4523) );
BUF_X2 newInst_1816 ( .a(newNet_1815), .o(newNet_1816) );
BUF_X2 newInst_1328 ( .a(newNet_1327), .o(newNet_1328) );
INV_X1 g35486 ( .a(U_0_), .o(n_3239) );
BUF_X2 newInst_555 ( .a(newNet_554), .o(newNet_555) );
BUF_X2 newInst_679 ( .a(newNet_381), .o(newNet_679) );
NAND2_Z01 g58041 ( .a(n_2903), .b(n_2226), .o(n_2944) );
NOR2_Z1 g59720 ( .a(n_1347), .b(pmem_d_7), .o(n_1407) );
INV_X1 g35487 ( .a(pmem_d_9), .o(n_3238) );
NAND2_Z01 g60515 ( .a(n_380), .b(GPR_4__6_), .o(n_631) );
NAND2_Z01 g59172 ( .a(n_1896), .b(n_476), .o(n_1934) );
AND2_X1 g57754 ( .a(n_3115), .b(n_571), .o(n_3131) );
NAND2_Z01 g57708 ( .a(n_3133), .b(n_2423), .o(n_3161) );
fflopd pZ_reg_7_ ( .CK(newNet_56), .D(n_3186), .Q(pZ_7_) );
NAND2_Z01 g59694 ( .a(io_do_1), .b(n_1353), .o(n_1436) );
NAND2_Z01 g59278 ( .a(n_63), .b(n_1766), .o(n_1850) );
NAND2_Z01 g34736 ( .a(n_3633), .b(pZ_13_), .o(n_3829) );
XOR2_X1 g35050 ( .a(n_3508), .b(pZ_7_), .o(n_3533) );
BUF_X2 newInst_1387 ( .a(newNet_1386), .o(newNet_1387) );
NAND2_Z01 g60409 ( .a(n_371), .b(GPR_21__7_), .o(n_737) );
NAND2_Z01 g60400 ( .a(n_414), .b(n_397), .o(n_746) );
NOR4_Z1 g59806 ( .a(n_504), .b(n_1146), .c(n_1143), .d(n_493), .o(n_1322) );
NAND2_Z01 g59280 ( .a(n_63), .b(n_1765), .o(n_1835) );
NAND2_Z01 g35171 ( .a(n_3198), .b(n_3269), .o(n_3461) );
NAND2_Z01 g60762 ( .a(n_195), .b(pmem_d_9), .o(n_461) );
NAND2_Z01 g58814 ( .a(n_2181), .b(n_1803), .o(n_2362) );
AND2_X1 g57901 ( .a(n_3009), .b(n_2204), .o(n_3037) );
fflopd GPR_reg_18__7_ ( .CK(newNet_1335), .D(n_3161), .Q(GPR_18__7_) );
NOR2_Z1 g34433 ( .a(n_4088), .b(n_3314), .o(n_4104) );
NOR2_Z1 g34311 ( .a(n_4159), .b(n_4044), .o(n_4222) );
NOR3_Z1 g60659 ( .a(n_116), .b(n_253), .c(n_125), .o(n_486) );
NAND2_Z01 g58720 ( .a(n_2207), .b(GPR_22__1_), .o(n_2387) );
NAND2_Z01 g35328 ( .a(pZ_4_), .b(n_3199), .o(n_3341) );
NAND2_Z01 g58574 ( .a(n_2459), .b(n_2031), .o(n_2522) );
NOR4_Z1 g34458 ( .a(n_3755), .b(n_3969), .c(n_4047), .d(n_3723), .o(n_4084) );
XOR2_X1 g35365 ( .a(pY_1_), .b(pmem_d_1), .o(n_3324) );
BUF_X2 newInst_1359 ( .a(newNet_556), .o(newNet_1359) );
NOR2_Z1 g60970 ( .a(n_4634), .b(n_4633), .o(n_195) );
NAND2_Z01 g57829 ( .a(n_3047), .b(n_2434), .o(n_3084) );
NOR2_Z1 g34389 ( .a(n_4084), .b(n_3469), .o(n_4149) );
NAND2_Z01 g58800 ( .a(n_2195), .b(U_13_), .o(n_2300) );
NOR2_Z1 g60617 ( .a(n_459), .b(n_182), .o(n_590) );
XOR2_X1 g59553 ( .a(n_1526), .b(n_65), .o(n_1600) );
AND2_X1 g34180 ( .a(n_4324), .b(pmem_d_0), .o(n_4336) );
BUF_X2 newInst_651 ( .a(newNet_650), .o(newNet_651) );
NAND4_Z1 g58349 ( .a(n_2567), .b(n_2657), .c(n_2656), .d(n_1535), .o(n_2721) );
BUF_X2 newInst_128 ( .a(newNet_127), .o(newNet_128) );
NAND2_Z01 final_adder_mux_R16_278_6_g426 ( .a(n_4449), .b(n_4433), .o(final_adder_mux_R16_278_6_n_22) );
NAND2_Z01 g34945 ( .a(n_3554), .b(PC_9_), .o(n_3617) );
XOR2_X1 g34462 ( .a(n_4055), .b(pZ_9_), .o(n_4080) );
NAND2_Z01 g59692 ( .a(n_1372), .b(n_1273), .o(n_1438) );
BUF_X2 newInst_588 ( .a(newNet_587), .o(newNet_588) );
BUF_X2 newInst_1142 ( .a(newNet_891), .o(newNet_1142) );
BUF_X2 newInst_1779 ( .a(newNet_1778), .o(newNet_1779) );
BUF_X2 newInst_847 ( .a(newNet_846), .o(newNet_847) );
BUF_X2 newInst_1074 ( .a(newNet_1073), .o(newNet_1074) );
INV_X1 g61113 ( .a(io_do_1), .o(n_39) );
INV_X1 g35462 ( .a(state_3_), .o(n_3262) );
NAND2_Z01 g60709 ( .a(n_198), .b(GPR_17__5_), .o(n_429) );
NAND2_Z01 g60213 ( .a(n_574), .b(GPR_10__0_), .o(n_932) );
BUF_X2 newInst_1851 ( .a(newNet_1850), .o(newNet_1851) );
BUF_X2 newInst_638 ( .a(newNet_637), .o(newNet_638) );
NAND4_Z1 g34593 ( .a(n_3710), .b(n_3712), .c(n_3709), .d(n_3711), .o(n_3967) );
BUF_X2 newInst_857 ( .a(newNet_856), .o(newNet_857) );
NAND4_Z1 g60140 ( .a(n_538), .b(n_707), .c(n_708), .d(n_704), .o(n_992) );
INV_X1 g34980 ( .a(n_3574), .o(n_3573) );
BUF_X2 newInst_1546 ( .a(newNet_1545), .o(newNet_1546) );
BUF_X2 newInst_0 ( .a(tau_clk), .o(newNet_0) );
XOR2_X1 g59674 ( .a(n_1389), .b(pmem_d_3), .o(n_1483) );
BUF_X2 newInst_1774 ( .a(newNet_1773), .o(newNet_1774) );
NAND2_Z03 g34221 ( .a(n_4284), .b(n_3440), .o(n_4556) );
NAND2_Z01 g60891 ( .a(n_4557), .b(n_119), .o(n_237) );
BUF_X2 newInst_1606 ( .a(newNet_1605), .o(newNet_1606) );
NAND2_Z01 g60485 ( .a(n_357), .b(pY_11_), .o(n_661) );
NAND2_Z01 g59136 ( .a(n_1872), .b(n_1282), .o(n_1962) );
NAND2_Z01 g59073 ( .a(n_1871), .b(n_4599), .o(n_2034) );
AND2_X1 g60745 ( .a(n_103), .b(n_250), .o(n_397) );
BUF_X2 newInst_795 ( .a(newNet_277), .o(newNet_795) );
AND2_X1 g59405 ( .a(n_64), .b(n_1649), .o(n_1711) );
NAND4_Z1 g59545 ( .a(n_788), .b(n_1299), .c(n_1504), .d(n_1077), .o(n_1583) );
NAND2_Z01 g58249 ( .a(n_2756), .b(n_2193), .o(n_2818) );
INV_X1 g61030 ( .a(PC_5_), .o(n_122) );
BUF_X2 newInst_615 ( .a(newNet_614), .o(newNet_615) );
BUF_X2 newInst_481 ( .a(newNet_480), .o(newNet_481) );
AND2_X1 g60329 ( .a(n_589), .b(n_43), .o(n_799) );
NAND2_Z01 g60215 ( .a(n_590), .b(GPR_6__2_), .o(n_930) );
NAND2_Z01 g60905 ( .a(PC_0_), .b(pmem_d_3), .o(n_266) );
NAND2_Z01 g58288 ( .a(n_2709), .b(n_2258), .o(n_2782) );
NAND2_Z01 g34146 ( .a(n_4317), .b(n_4625), .o(n_4362) );
NAND4_Z1 g59532 ( .a(n_824), .b(n_826), .c(n_1471), .d(n_913), .o(n_1595) );
NAND2_Z01 g58146 ( .a(n_2820), .b(n_2296), .o(n_2867) );
NAND2_Z02 g34379 ( .a(n_4643), .b(n_4092), .o(n_4612) );
BUF_X2 newInst_180 ( .a(newNet_179), .o(newNet_180) );
NAND2_Z01 g58900 ( .a(n_2155), .b(GPR_14__4_), .o(n_2182) );
NAND2_Z01 g34645 ( .a(n_4539), .b(n_3768), .o(n_3915) );
INV_X2 newInst_516 ( .a(newNet_515), .o(newNet_516) );
NOR2_Z1 g34605 ( .a(n_3736), .b(n_3668), .o(n_3955) );
XOR2_X1 g59289 ( .a(io_do_0), .b(n_1695), .o(n_1832) );
BUF_X2 newInst_460 ( .a(newNet_459), .o(newNet_460) );
NAND2_Z01 g34769 ( .a(n_3599), .b(GPR_5__4_), .o(n_3796) );
BUF_X2 newInst_1617 ( .a(newNet_1616), .o(newNet_1617) );
BUF_X2 newInst_675 ( .a(newNet_674), .o(newNet_675) );
XOR2_X1 final_adder_mux_R16_278_6_g379 ( .a(final_adder_mux_R16_278_6_n_68), .b(final_adder_mux_R16_278_6_n_44), .o(R16_9_) );
BUF_X2 newInst_1713 ( .a(newNet_1712), .o(newNet_1713) );
NAND2_Z01 g34845 ( .a(n_3585), .b(GPR_13__1_), .o(n_3718) );
NOR2_Z4 g58452 ( .a(n_2609), .b(n_1580), .o(n_2656) );
BUF_X2 newInst_763 ( .a(newNet_762), .o(newNet_763) );
BUF_X2 newInst_380 ( .a(newNet_379), .o(newNet_380) );
BUF_X2 newInst_338 ( .a(newNet_337), .o(newNet_338) );
BUF_X2 newInst_67 ( .a(newNet_66), .o(newNet_67) );
NOR2_Z1 g59431 ( .a(n_1646), .b(n_603), .o(n_1688) );
BUF_X2 newInst_1749 ( .a(newNet_1748), .o(newNet_1749) );
BUF_X2 newInst_77 ( .a(newNet_51), .o(newNet_77) );
NAND4_Z1 g58279 ( .a(n_1330), .b(n_2175), .c(n_2643), .d(n_1333), .o(n_2789) );
BUF_X2 newInst_631 ( .a(newNet_186), .o(newNet_631) );
NAND2_Z01 g34692 ( .a(n_3590), .b(pY_15_), .o(n_3873) );
BUF_X2 newInst_1643 ( .a(newNet_1642), .o(newNet_1643) );
AND2_X1 g59241 ( .a(n_1825), .b(n_850), .o(n_1865) );
NOR2_Z1 g35133 ( .a(n_3468), .b(n_4651), .o(n_3474) );
BUF_X2 newInst_1156 ( .a(newNet_1155), .o(newNet_1156) );
NAND2_Z01 g59756 ( .a(n_1312), .b(io_do_5), .o(n_1368) );
NAND2_Z01 g60439 ( .a(n_360), .b(GPR_3__1_), .o(n_707) );
NOR2_Z1 g60310 ( .a(n_616), .b(n_126), .o(n_866) );
NAND2_Z01 g59776 ( .a(n_1268), .b(n_331), .o(n_1354) );
NAND2_Z01 g35350 ( .a(n_3285), .b(n_3243), .o(n_3355) );
NAND2_Z01 g60426 ( .a(n_361), .b(GPR_5__5_), .o(n_720) );
NAND2_Z01 g60730 ( .a(n_178), .b(n_4534), .o(n_409) );
NAND2_Z01 g60566 ( .a(n_467), .b(pZ_3_), .o(n_616) );
NAND2_Z01 g34204 ( .a(io_do_4), .b(n_4177), .o(n_4322) );
NAND2_Z01 g58852 ( .a(n_2158), .b(GPR_12__5_), .o(n_2255) );
NAND2_Z01 g58151 ( .a(n_2814), .b(n_2252), .o(n_2862) );
BUF_X2 newInst_1751 ( .a(newNet_1750), .o(newNet_1751) );
NAND2_Z01 g34176 ( .a(n_4325), .b(n_4471), .o(n_4340) );
XOR2_X1 g59371 ( .a(io_do_1), .b(n_1664), .o(n_1767) );
NAND2_Z01 g34398 ( .a(n_3208), .b(pZ_6_), .o(n_4140) );
NAND2_Z01 g59828 ( .a(n_1171), .b(dmem_di_7), .o(n_1296) );
NAND2_Z01 g60783 ( .a(n_166), .b(n_262), .o(n_320) );
fflopd U_reg_10_ ( .CK(newNet_440), .D(n_2869), .Q(U_10_) );
INV_X1 g59740 ( .a(n_1387), .o(n_1386) );
NAND2_Z01 g59482 ( .a(n_27), .b(n_753), .o(n_1643) );
NAND2_Z01 g34863 ( .a(n_3584), .b(GPR_21__0_), .o(n_3700) );
BUF_X2 newInst_1730 ( .a(newNet_1729), .o(newNet_1730) );
NAND2_Z01 g34750 ( .a(n_3197), .b(GPR_23__5_), .o(n_3815) );
NAND2_Z01 g34616 ( .a(n_3896), .b(n_3481), .o(n_3944) );
NAND2_Z01 g57712 ( .a(n_3128), .b(n_2389), .o(n_3155) );
NAND4_Z1 g59667 ( .a(n_1070), .b(n_1291), .c(n_1368), .d(n_1069), .o(n_1461) );
NAND2_Z01 g57692 ( .a(n_3158), .b(n_2215), .o(n_3174) );
NAND2_Z01 g58599 ( .a(n_2479), .b(n_1959), .o(n_2496) );
BUF_X2 newInst_560 ( .a(newNet_559), .o(newNet_560) );
NOR2_Z1 g60641 ( .a(n_348), .b(io_do_3), .o(n_576) );
NAND2_Z01 g34308 ( .a(n_4166), .b(n_4545), .o(n_4225) );
BUF_X2 newInst_1321 ( .a(newNet_1320), .o(newNet_1321) );
NAND2_Z01 g58603 ( .a(n_2459), .b(n_1953), .o(n_2492) );
XOR2_X1 g60160 ( .a(n_593), .b(SP_4_), .o(n_976) );
INV_X1 drc_bufs35540 ( .a(n_4530), .o(n_3201) );
NAND2_Z01 g58725 ( .a(n_2207), .b(GPR_22__6_), .o(n_2382) );
NOR2_Z1 g34696 ( .a(n_3570), .b(n_4400), .o(n_3869) );
BUF_X2 newInst_1649 ( .a(newNet_1648), .o(newNet_1649) );
AND4_X1 g59040 ( .a(n_4614), .b(n_4682), .c(n_1810), .d(n_4617), .o(n_2082) );
BUF_X2 newInst_1860 ( .a(newNet_1859), .o(newNet_1860) );
NOR3_Z1 g58939 ( .a(n_1754), .b(n_2096), .c(n_1798), .o(n_2168) );
INV_X1 g59019 ( .a(n_2089), .o(n_2088) );
NAND2_Z01 g58173 ( .a(n_873), .b(n_2834), .o(n_2852) );
XOR2_X1 g59451 ( .a(n_1628), .b(n_101), .o(n_1671) );
NAND2_Z01 g59652 ( .a(n_1268), .b(n_1396), .o(n_1473) );
NAND2_Z01 g34314 ( .a(n_4166), .b(n_4547), .o(n_4219) );
NAND4_Z1 g59662 ( .a(n_815), .b(n_946), .c(n_1361), .d(n_918), .o(n_1465) );
NAND2_Z01 g60511 ( .a(n_361), .b(GPR_5__7_), .o(n_635) );
BUF_X2 newInst_775 ( .a(newNet_774), .o(newNet_775) );
NAND2_Z01 g60713 ( .a(n_257), .b(n_4684), .o(n_425) );
BUF_X2 newInst_406 ( .a(newNet_405), .o(newNet_406) );
BUF_X2 newInst_377 ( .a(newNet_376), .o(newNet_377) );
NAND2_Z01 g60966 ( .a(n_55), .b(pmem_d_9), .o(n_154) );
BUF_X2 newInst_75 ( .a(newNet_70), .o(newNet_75) );
INV_X1 g61066 ( .a(PC_3_), .o(n_86) );
NAND2_Z01 g58809 ( .a(n_2197), .b(U_7_), .o(n_2291) );
fflopd GPR_reg_23__6_ ( .CK(newNet_1035), .D(n_3073), .Q(GPR_23__6_) );
BUF_X2 newInst_1207 ( .a(newNet_1206), .o(newNet_1207) );
BUF_X2 newInst_1704 ( .a(newNet_1703), .o(newNet_1704) );
BUF_X2 newInst_658 ( .a(newNet_657), .o(newNet_658) );
NAND2_Z01 g61017 ( .a(n_87), .b(n_44), .o(n_129) );
NAND4_Z1 g34124 ( .a(n_4251), .b(n_4275), .c(n_4309), .d(n_4116), .o(n_4382) );
NOR2_Z1 g34239 ( .a(n_4230), .b(n_3246), .o(n_4294) );
NAND2_Z01 g60253 ( .a(n_584), .b(GPR_18__7_), .o(n_893) );
NAND3_Z1 g58343 ( .a(n_2473), .b(n_2646), .c(n_2109), .o(n_2726) );
NOR2_Z1 g60839 ( .a(n_197), .b(n_248), .o(n_342) );
NAND2_Z01 g58171 ( .a(n_2795), .b(n_2220), .o(n_2839) );
BUF_X2 newInst_1460 ( .a(newNet_1459), .o(newNet_1460) );
INV_X1 g61094 ( .a(n_4628), .o(n_58) );
NAND2_Z01 g60204 ( .a(n_578), .b(GPR_19__3_), .o(n_941) );
NAND4_Z1 g60379 ( .a(n_430), .b(n_454), .c(n_429), .d(n_451), .o(n_766) );
BUF_X2 newInst_161 ( .a(newNet_160), .o(newNet_161) );
XOR2_X1 g34384 ( .a(n_4095), .b(pY_12_), .o(n_4154) );
AND2_X1 g58509 ( .a(n_2567), .b(n_2207), .o(n_2587) );
NAND2_Z01 g59143 ( .a(n_1894), .b(n_475), .o(n_1956) );
NOR2_Z1 g34357 ( .a(n_4149), .b(n_3661), .o(n_4174) );
NAND2_Z01 g60042 ( .a(n_856), .b(n_4605), .o(n_1088) );
fflopd GPR_reg_11__7_ ( .CK(newNet_1678), .D(n_3169), .Q(GPR_11__7_) );
BUF_X2 newInst_968 ( .a(newNet_967), .o(newNet_968) );
BUF_X2 newInst_602 ( .a(newNet_601), .o(newNet_602) );
NAND2_Z01 g34309 ( .a(n_4158), .b(n_4062), .o(n_4224) );
NAND2_Z01 g60191 ( .a(n_4556), .b(n_673), .o(n_954) );
NAND2_Z01 g58580 ( .a(n_2465), .b(pY_7_), .o(n_2518) );
XOR2_X1 final_adder_mux_R16_278_6_g397 ( .a(final_adder_mux_R16_278_6_n_50), .b(final_adder_mux_R16_278_6_n_38), .o(R16_3_) );
NAND4_Z1 g57657 ( .a(n_1913), .b(n_1925), .c(n_3173), .d(n_1430), .o(n_3185) );
AND2_X1 g58124 ( .a(n_2850), .b(n_2201), .o(n_2888) );
NAND2_Z01 g58741 ( .a(n_2205), .b(GPR_2__6_), .o(n_2366) );
BUF_X2 newInst_95 ( .a(newNet_94), .o(newNet_95) );
BUF_X2 newInst_1833 ( .a(newNet_1832), .o(newNet_1833) );
BUF_X2 newInst_1668 ( .a(newNet_236), .o(newNet_1668) );
NAND2_Z01 g34283 ( .a(n_4162), .b(pY_10_), .o(n_4250) );
BUF_X2 newInst_1343 ( .a(newNet_1342), .o(newNet_1343) );
NOR2_Z1 g60030 ( .a(n_840), .b(n_378), .o(n_1099) );
NOR2_Z1 g34172 ( .a(n_4324), .b(n_4644), .o(n_4421) );
NOR3_Z2 g60152 ( .a(n_568), .b(n_4556), .c(pmem_d_9), .o(n_1026) );
NOR2_Z1 g59760 ( .a(n_1218), .b(n_1288), .o(n_1388) );
AND2_X1 g58007 ( .a(n_2940), .b(n_2201), .o(n_2964) );
NOR2_Z1 g60096 ( .a(n_842), .b(pmem_d_7), .o(n_1023) );
NAND2_Z01 g57882 ( .a(n_3011), .b(n_2196), .o(n_3057) );
NAND2_Z01 g35159 ( .a(n_3198), .b(pmem_d_6), .o(n_3467) );
INV_X1 g60534 ( .a(n_599), .o(n_600) );
NAND2_Z01 g60292 ( .a(n_578), .b(GPR_19__5_), .o(n_832) );
NAND2_Z01 g60472 ( .a(n_380), .b(GPR_4__3_), .o(n_674) );
NAND2_Z01 g58737 ( .a(n_2205), .b(GPR_2__2_), .o(n_2370) );
NAND4_Z2 g35195 ( .a(n_3340), .b(n_3381), .c(n_3371), .d(n_3396), .o(n_4620) );
NOR2_Z1 g59947 ( .a(n_1112), .b(n_4525), .o(n_1205) );
BUF_X2 newInst_1180 ( .a(newNet_1179), .o(newNet_1180) );
NAND3_Z1 g60843 ( .a(pmem_d_4), .b(n_48), .c(pmem_d_6), .o(n_339) );
BUF_X2 newInst_491 ( .a(newNet_490), .o(newNet_491) );
INV_X2 newInst_469 ( .a(newNet_468), .o(newNet_469) );
NAND2_Z01 g58709 ( .a(n_2209), .b(GPR_20__6_), .o(n_2398) );
INV_X1 g35502 ( .a(pmem_d_5), .o(n_3225) );
NAND2_Z01 g59064 ( .a(n_1902), .b(n_4590), .o(n_2043) );
NAND2_Z01 g58796 ( .a(n_2197), .b(U_0_), .o(n_2304) );
BUF_X2 newInst_1545 ( .a(newNet_1544), .o(newNet_1545) );
NOR2_Z1 g34302 ( .a(n_4159), .b(n_4080), .o(n_4232) );
NOR2_Z1 g58563 ( .a(n_2485), .b(n_1619), .o(n_2535) );
NAND4_Z1 g59995 ( .a(n_935), .b(n_926), .c(n_939), .d(n_875), .o(n_1134) );
INV_X1 g59232 ( .a(n_1879), .o(n_1880) );
BUF_X1 mybuffer3 ( .o(io_a_3), .a(pmem_d_3) );
NAND2_Z01 g58674 ( .a(n_2213), .b(GPR_17__0_), .o(n_2432) );
NAND2_Z01 g60222 ( .a(n_580), .b(GPR_14__5_), .o(n_923) );
NAND2_Z01 g34672 ( .a(n_3607), .b(n_3608), .o(n_3893) );
fflopd GPR_reg_17__4_ ( .CK(newNet_1389), .D(n_2938), .Q(GPR_17__4_) );
INV_X1 drc_bufs35536 ( .a(n_4620), .o(n_3202) );
NOR2_Z1 g34288 ( .a(n_4163), .b(n_3254), .o(n_4245) );
BUF_X2 newInst_1792 ( .a(newNet_1791), .o(newNet_1792) );
BUF_X2 newInst_1576 ( .a(newNet_1575), .o(newNet_1576) );
NAND2_Z01 g34802 ( .a(n_3592), .b(GPR_23__3_), .o(n_3761) );
NAND3_Z1 g59894 ( .a(io_do_2), .b(n_1026), .c(n_56), .o(n_1235) );
NAND2_Z01 g34771 ( .a(n_3592), .b(GPR_23__4_), .o(n_3794) );
BUF_X2 newInst_1178 ( .a(newNet_1177), .o(newNet_1178) );
NAND4_Z2 g60658 ( .a(n_36), .b(n_71), .c(n_4658), .d(pmem_d_13), .o(n_568) );
NAND2_Z01 g58704 ( .a(n_2209), .b(GPR_20__1_), .o(n_2403) );
BUF_X2 newInst_467 ( .a(newNet_466), .o(newNet_467) );
BUF_X2 newInst_1246 ( .a(newNet_1245), .o(newNet_1246) );
BUF_X2 newInst_835 ( .a(newNet_834), .o(newNet_835) );
NAND2_Z01 g58351 ( .a(n_2649), .b(n_1735), .o(n_2720) );
NAND2_Z01 g35112 ( .a(n_3458), .b(n_3304), .o(n_3494) );
BUF_X2 newInst_1254 ( .a(newNet_1253), .o(newNet_1254) );
NOR2_Z1 g35415 ( .a(n_3233), .b(n_3248), .o(n_4668) );
BUF_X2 newInst_1301 ( .a(newNet_1300), .o(newNet_1301) );
AND2_X1 g58258 ( .a(n_2752), .b(n_2212), .o(n_2809) );
BUF_X2 newInst_1502 ( .a(newNet_1501), .o(newNet_1502) );
BUF_X2 newInst_147 ( .a(newNet_146), .o(newNet_147) );
AND2_X1 g59953 ( .a(n_177), .b(n_1049), .o(n_1200) );
NAND2_Z01 g59634 ( .a(n_1422), .b(SP_0_), .o(n_1495) );
INV_X2 newInst_1127 ( .a(newNet_1126), .o(newNet_1127) );
INV_X2 g61090 ( .a(pmem_d_0), .o(n_62) );
fflopd GPR_reg_22__2_ ( .CK(newNet_1102), .D(n_2760), .Q(GPR_22__2_) );
AND2_X1 g59935 ( .a(n_1043), .b(n_48), .o(n_1208) );
NAND2_Z01 g57825 ( .a(n_3051), .b(n_2239), .o(n_3088) );
NAND2_Z01 g58750 ( .a(n_2204), .b(GPR_3__2_), .o(n_2350) );
NAND2_Z01 g60523 ( .a(n_371), .b(GPR_23__4_), .o(n_623) );
NAND2_Z01 g58629 ( .a(n_2353), .b(n_2013), .o(n_2481) );
NAND2_Z01 g59097 ( .a(n_1902), .b(n_354), .o(n_2011) );
XOR2_X1 g34479 ( .a(n_4038), .b(pY_8_), .o(n_4063) );
NAND2_Z01 g34528 ( .a(n_3959), .b(pY_6_), .o(n_4026) );
AND3_X1 g60367 ( .a(n_311), .b(n_406), .c(n_4685), .o(n_774) );
XOR2_X1 g60009 ( .a(n_863), .b(pmem_d_1), .o(n_1156) );
NAND2_Z01 g59645 ( .a(io_do_2), .b(n_1418), .o(n_1476) );
BUF_X2 newInst_838 ( .a(newNet_339), .o(newNet_838) );
NOR2_Z1 g59914 ( .a(n_1100), .b(n_1099), .o(n_1198) );
INV_Y1 g35148 ( .a(n_3469), .o(Rd_0_) );
NAND2_Z01 g58887 ( .a(n_2140), .b(GPR_9__3_), .o(n_2220) );
AND2_X1 g58117 ( .a(n_2850), .b(n_2207), .o(n_2895) );
NAND2_Z01 g60502 ( .a(n_347), .b(GPR_9__7_), .o(n_644) );
NAND4_Z1 g60378 ( .a(n_437), .b(n_447), .c(n_422), .d(n_419), .o(n_767) );
AND2_X1 g58497 ( .a(n_2567), .b(n_2139), .o(n_2600) );
NAND2_Z01 g35152 ( .a(n_3446), .b(pmem_d_14), .o(n_3459) );
fflopd pZ_reg_1_ ( .CK(newNet_81), .D(n_2874), .Q(pZ_1_) );
NAND2_Z03 g34295 ( .a(n_4170), .b(n_4066), .o(io_do_5) );
NAND2_Z01 final_adder_mux_R16_278_6_g403 ( .a(final_adder_mux_R16_278_6_n_45), .b(final_adder_mux_R16_278_6_n_16), .o(final_adder_mux_R16_278_6_n_46) );
NAND2_Z01 g60914 ( .a(n_111), .b(pZ_7_), .o(n_227) );
NAND2_Z01 g58857 ( .a(n_2157), .b(GPR_13__5_), .o(n_2250) );
BUF_X2 newInst_736 ( .a(newNet_735), .o(newNet_736) );
BUF_X2 newInst_608 ( .a(newNet_607), .o(newNet_608) );
NAND2_Z01 g58705 ( .a(n_2209), .b(GPR_20__2_), .o(n_2402) );
NAND2_Z01 g34676 ( .a(n_3635), .b(GPR_14__7_), .o(n_3889) );
AND2_X1 g60993 ( .a(n_4446), .b(n_4430), .o(n_179) );
BUF_X2 newInst_1728 ( .a(newNet_1727), .o(newNet_1728) );
INV_X1 g59815 ( .a(n_1310), .o(n_1311) );
AND2_X1 g35238 ( .a(n_4631), .b(n_4483), .o(n_3430) );
NOR4_Z1 g58528 ( .a(n_4663), .b(n_1530), .c(n_2527), .d(state_0_), .o(n_2569) );
INV_X1 g61050 ( .a(pX_8_), .o(n_102) );
NAND2_Z01 g59078 ( .a(n_1875), .b(n_4569), .o(n_2029) );
AND2_X1 g35314 ( .a(n_3230), .b(n_3309), .o(n_3363) );
NAND4_Z1 g34577 ( .a(n_3804), .b(n_3803), .c(n_3681), .d(n_3802), .o(n_3983) );
NAND4_Z1 g58136 ( .a(n_1956), .b(n_2467), .c(n_2824), .d(n_2048), .o(n_2877) );
AND3_X1 g34497 ( .a(n_3968), .b(n_4004), .c(n_4015), .o(n_4047) );
XNOR2_X1 g60166 ( .a(n_616), .b(pZ_4_), .o(n_971) );
NAND4_Z1 g59254 ( .a(n_1428), .b(n_1525), .c(n_1750), .d(n_1258), .o(n_1858) );
XOR2_X1 g60670 ( .a(n_164), .b(n_118), .o(n_479) );
BUF_X2 newInst_1679 ( .a(newNet_1490), .o(newNet_1679) );
NAND4_Z1 g58016 ( .a(n_1941), .b(n_2466), .c(n_2914), .d(n_2044), .o(n_2956) );
fflopd U_reg_12_ ( .CK(newNet_424), .D(n_3023), .Q(U_12_) );
NAND2_Z01 g58743 ( .a(n_2205), .b(GPR_2__7_), .o(n_2364) );
BUF_X2 newInst_359 ( .a(newNet_358), .o(newNet_359) );
AND2_X1 g60598 ( .a(n_4556), .b(n_346), .o(n_601) );
NOR2_Z4 g58344 ( .a(n_2717), .b(n_1588), .o(n_2752) );
NOR4_Z1 g59966 ( .a(pmem_d_9), .b(n_36), .c(n_645), .d(pmem_d_11), .o(n_1153) );
NAND2_Z01 final_adder_mux_R16_278_6_g369 ( .a(final_adder_mux_R16_278_6_n_78), .b(final_adder_mux_R16_278_6_n_18), .o(final_adder_mux_R16_278_6_n_80) );
AND2_X1 g60972 ( .a(n_4558), .b(n_4637), .o(n_150) );
fflopd GPR_reg_12__2_ ( .CK(newNet_1656), .D(n_2782), .Q(GPR_12__2_) );
NAND2_Z01 g60498 ( .a(n_457), .b(GPR_16__3_), .o(n_648) );
NAND2_Z01 g34109 ( .a(n_4337), .b(n_4351), .o(n_4449) );
NAND2_Z01 g34793 ( .a(n_3597), .b(GPR_17__3_), .o(n_3772) );
AND2_X1 g59024 ( .a(n_1982), .b(pZ_8_), .o(n_2078) );
NAND2_Z01 g59158 ( .a(n_1902), .b(n_572), .o(n_1942) );
AND2_X1 g60818 ( .a(n_177), .b(n_4531), .o(n_308) );
BUF_X2 newInst_1112 ( .a(newNet_1111), .o(newNet_1112) );
INV_X1 g61071 ( .a(SP_11_), .o(n_81) );
NOR4_Z1 g58985 ( .a(n_1830), .b(n_1769), .c(n_1864), .d(n_1879), .o(n_2122) );
NAND2_Z01 g35237 ( .a(n_3352), .b(n_3252), .o(n_4639) );
AND2_X1 g60988 ( .a(n_4442), .b(n_4426), .o(n_184) );
AND2_X1 g57733 ( .a(n_3115), .b(n_2157), .o(n_3139) );
BUF_X2 newInst_374 ( .a(newNet_373), .o(newNet_374) );
BUF_X2 newInst_1155 ( .a(newNet_1154), .o(newNet_1155) );
NAND2_Z01 g57838 ( .a(n_3038), .b(n_2366), .o(n_3072) );
BUF_X2 newInst_1317 ( .a(newNet_1316), .o(newNet_1317) );
NAND2_Z01 g35032 ( .a(n_4515), .b(n_3253), .o(n_3547) );
NAND2_Z01 g34743 ( .a(n_3594), .b(GPR_7__3_), .o(n_3822) );
BUF_X2 newInst_909 ( .a(newNet_908), .o(newNet_909) );
BUF_X2 newInst_856 ( .a(newNet_855), .o(newNet_856) );
AND2_X1 g35439 ( .a(state_0_), .b(state_1_), .o(n_4637) );
AND2_X1 g60068 ( .a(n_845), .b(n_36), .o(n_1066) );
BUF_X2 newInst_574 ( .a(newNet_573), .o(newNet_574) );
NAND2_Z01 g35002 ( .a(n_3509), .b(n_3536), .o(n_3578) );
NAND2_Z01 g35081 ( .a(n_3494), .b(n_3282), .o(n_3504) );
NOR2_Z1 g60649 ( .a(n_327), .b(n_191), .o(n_492) );
NAND2_Z01 g58773 ( .a(n_2201), .b(GPR_6__1_), .o(n_2327) );
INV_X1 g35500 ( .a(state_1_), .o(n_3227) );
NAND2_Z01 g60262 ( .a(n_598), .b(GPR_15__6_), .o(n_884) );
NAND2_Z01 g58972 ( .a(n_31), .b(n_2062), .o(n_2134) );
NAND2_Z01 g60438 ( .a(n_347), .b(GPR_11__1_), .o(n_708) );
NAND2_Z01 g35371 ( .a(n_3284), .b(n_3303), .o(n_3319) );
NAND2_Z01 g34738 ( .a(n_3599), .b(GPR_5__5_), .o(n_3827) );
NAND2_Z01 g59746 ( .a(n_1232), .b(n_676), .o(n_1376) );
AND2_X1 g58266 ( .a(n_2752), .b(n_2204), .o(n_2801) );
BUF_X2 newInst_1279 ( .a(newNet_1278), .o(newNet_1279) );
NAND4_Z1 g60003 ( .a(n_893), .b(n_894), .c(n_934), .d(n_892), .o(n_1126) );
NOR2_Z1 g34509 ( .a(n_4027), .b(n_3215), .o(n_4037) );
BUF_X2 newInst_65 ( .a(newNet_64), .o(newNet_65) );
INV_X1 g35231 ( .a(n_4485), .o(n_3423) );
NAND4_Z1 g58924 ( .a(n_1727), .b(n_2024), .c(n_2105), .d(n_1092), .o(n_2179) );
NAND3_Z1 g34069 ( .a(n_4393), .b(n_4386), .c(n_4238), .o(dmem_do_7) );
BUF_X2 newInst_1386 ( .a(newNet_1385), .o(newNet_1386) );
NOR2_Z1 g59710 ( .a(n_1346), .b(io_do_0), .o(n_1412) );
NAND2_Z01 g59162 ( .a(n_1898), .b(n_192), .o(n_1938) );
BUF_X2 newInst_1632 ( .a(newNet_1631), .o(newNet_1632) );
XOR2_X1 g35078 ( .a(n_3495), .b(pmem_d_10), .o(n_3513) );
NAND2_Z01 g60650 ( .a(n_322), .b(n_193), .o(n_491) );
NAND2_Z02 g58918 ( .a(n_2152), .b(n_1202), .o(n_2204) );
BUF_X2 newInst_715 ( .a(newNet_714), .o(newNet_715) );
BUF_X2 newInst_226 ( .a(newNet_56), .o(newNet_226) );
BUF_X2 newInst_1167 ( .a(newNet_1083), .o(newNet_1167) );
AND2_X1 g58971 ( .a(n_2063), .b(n_587), .o(n_2135) );
NOR2_Z2 g34377 ( .a(n_4643), .b(n_4645), .o(n_4164) );
BUF_X2 newInst_232 ( .a(newNet_231), .o(newNet_232) );
NOR2_Z1 g34246 ( .a(n_4181), .b(n_4178), .o(n_4287) );
AND2_X1 g57893 ( .a(n_3009), .b(n_2212), .o(n_3045) );
BUF_X2 newInst_1025 ( .a(newNet_1024), .o(newNet_1025) );
NAND2_Z01 g60231 ( .a(n_597), .b(pX_15_), .o(n_914) );
INV_X1 g35509 ( .a(pY_12_), .o(n_3219) );
NAND2_Z01 g34294 ( .a(n_4164), .b(pmem_d_0), .o(n_4239) );
BUF_X2 newInst_1702 ( .a(newNet_1701), .o(newNet_1702) );
NOR2_Z1 g35452 ( .a(pX_1_), .b(pX_0_), .o(n_3277) );
BUF_X2 newInst_830 ( .a(newNet_829), .o(newNet_830) );
NOR2_Z1 g60801 ( .a(n_276), .b(n_260), .o(n_366) );
NOR2_Z1 g34922 ( .a(n_3560), .b(n_3280), .o(n_3643) );
BUF_X2 newInst_1101 ( .a(newNet_1100), .o(newNet_1101) );
BUF_X2 newInst_1820 ( .a(newNet_1819), .o(newNet_1820) );
BUF_X2 newInst_1239 ( .a(newNet_1238), .o(newNet_1239) );
fflopd PC_reg_4_ ( .CK(newNet_624), .D(n_1), .Q(PC_4_) );
NAND2_Z01 g58059 ( .a(n_2885), .b(n_2192), .o(n_2923) );
NAND2_Z01 g34850 ( .a(n_3579), .b(GPR_12__0_), .o(n_3713) );
BUF_X2 newInst_29 ( .a(newNet_28), .o(newNet_29) );
NOR2_Z1 g60601 ( .a(n_330), .b(n_168), .o(n_518) );
NAND2_Z01 g59614 ( .a(n_1413), .b(io_sp_1_), .o(n_1513) );
NAND4_Z1 g58653 ( .a(n_1770), .b(n_1876), .c(n_2122), .d(n_2087), .o(n_2449) );
NOR2_Z1 g35220 ( .a(n_4660), .b(n_3217), .o(n_3435) );
NAND2_Z01 g59298 ( .a(n_1769), .b(n_1037), .o(n_1814) );
NOR3_Z1 g34564 ( .a(n_3683), .b(n_3958), .c(n_3659), .o(n_3996) );
NAND2_Z01 g58535 ( .a(n_2531), .b(pX_15_), .o(n_2562) );
INV_X1 drc_bufs35559 ( .a(n_3309), .o(n_3199) );
fflopd GPR_reg_13__7_ ( .CK(newNet_1589), .D(n_3166), .Q(GPR_13__7_) );
BUF_X2 newInst_735 ( .a(newNet_734), .o(newNet_735) );
AND2_X1 g57907 ( .a(n_3009), .b(n_2140), .o(n_3031) );
NAND2_Z01 g60025 ( .a(n_967), .b(n_966), .o(n_1118) );
NAND2_Z01 g34537 ( .a(n_3931), .b(n_3538), .o(n_4599) );
NAND2_Z01 g34804 ( .a(n_3579), .b(GPR_12__2_), .o(n_3759) );
BUF_X2 newInst_1160 ( .a(newNet_1159), .o(newNet_1160) );
INV_X1 g59527 ( .a(n_1601), .o(n_1602) );
fflopd GPR_reg_6__5_ ( .CK(newNet_805), .D(n_2999), .Q(GPR_6__5_) );
BUF_X2 newInst_1169 ( .a(newNet_1168), .o(newNet_1169) );
AND2_X1 g59970 ( .a(n_1034), .b(n_205), .o(n_1168) );
NAND2_Z01 g34133 ( .a(n_4325), .b(n_4644), .o(n_4375) );
NAND4_Z1 g34589 ( .a(n_3731), .b(n_3733), .c(n_3730), .d(n_3732), .o(n_3971) );
NAND2_Z01 g34971 ( .a(n_3551), .b(n_3491), .o(n_3626) );
NAND2_Z01 g60553 ( .a(n_400), .b(n_401), .o(n_553) );
BUF_X2 newInst_1736 ( .a(newNet_1735), .o(newNet_1736) );
NAND2_Z01 g60591 ( .a(n_330), .b(n_168), .o(n_523) );
AND2_X1 g58499 ( .a(n_2567), .b(n_2157), .o(n_2598) );
XOR2_X1 g60853 ( .a(n_83), .b(pmem_d_9), .o(n_289) );
NOR2_Z2 g35428 ( .a(n_3225), .b(pmem_d_4), .o(n_3289) );
NAND2_Z01 final_adder_mux_R16_278_6_g435 ( .a(n_4446), .b(n_4430), .o(final_adder_mux_R16_278_6_n_14) );
NAND2_Z02 g58912 ( .a(n_2152), .b(n_1204), .o(n_2210) );
BUF_X1 drc_bufs61249 ( .a(n_2169), .o(n_2) );
NAND2_Z01 g60399 ( .a(n_236), .b(n_425), .o(n_747) );
NOR2_Z1 g34345 ( .a(n_16064_BAR), .b(n_3345), .o(n_4189) );
BUF_X2 newInst_1650 ( .a(newNet_1649), .o(newNet_1650) );
NOR2_Z1 g60615 ( .a(n_8), .b(pmem_d_3), .o(n_509) );
NOR2_Z1 g34469 ( .a(n_4647), .b(n_4025), .o(n_4071) );
NOR2_Z1 g59582 ( .a(n_1491), .b(n_461), .o(n_1549) );
INV_X1 drc_bufs61246 ( .a(n_1700), .o(n_3) );
BUF_X2 newInst_1367 ( .a(newNet_1366), .o(newNet_1367) );
AND2_X1 g58955 ( .a(n_2091), .b(pZ_15_), .o(n_2145) );
AND2_X1 g58104 ( .a(n_2850), .b(n_2159), .o(n_2909) );
AND2_X1 g35086 ( .a(n_3479), .b(n_3430), .o(n_3502) );
BUF_X2 newInst_630 ( .a(newNet_629), .o(newNet_630) );
AND2_X1 g58512 ( .a(n_2567), .b(n_2204), .o(n_2584) );
NAND2_Z01 g34102 ( .a(n_4359), .b(n_4358), .o(n_4444) );
NAND2_Z01 g34081 ( .a(n_4164), .b(GPR_Rd_r_3_), .o(n_4392) );
BUF_X2 newInst_1106 ( .a(newNet_283), .o(newNet_1106) );
AND2_X1 g34444 ( .a(n_4074), .b(n_3235), .o(n_4095) );
BUF_X2 newInst_1272 ( .a(newNet_1271), .o(newNet_1272) );
AND2_X1 g58406 ( .a(n_2656), .b(n_2199), .o(n_2662) );
BUF_X2 newInst_1077 ( .a(newNet_614), .o(newNet_1077) );
NAND2_Z01 g60500 ( .a(n_457), .b(GPR_16__7_), .o(n_646) );
INV_X1 g59961 ( .a(n_1167), .o(n_1166) );
NAND2_Z01 g60727 ( .a(n_200), .b(GPR_13__4_), .o(n_411) );
NAND2_Z01 g58711 ( .a(n_2208), .b(GPR_21__0_), .o(n_2396) );
AND3_X1 g34477 ( .a(n_4560), .b(n_4035), .c(n_3280), .o(n_4065) );
BUF_X2 newInst_727 ( .a(newNet_726), .o(newNet_727) );
NOR2_Z1 g60626 ( .a(n_328), .b(n_190), .o(n_504) );
NAND2_Z01 g57699 ( .a(n_3117), .b(n_2287), .o(n_3170) );
BUF_X2 newInst_432 ( .a(newNet_431), .o(newNet_432) );
BUF_X2 newInst_157 ( .a(newNet_156), .o(newNet_157) );
NAND2_Z01 g60084 ( .a(n_851), .b(n_122), .o(n_1106) );
fflopd GPR_reg_3__1_ ( .CK(newNet_966), .D(n_2748), .Q(GPR_3__1_) );
fflopd GPR_reg_15__1_ ( .CK(newNet_1514), .D(n_2776), .Q(GPR_15__1_) );
NAND2_Z01 g59318 ( .a(n_1699), .b(dmem_di_2), .o(n_1795) );
NAND2_Z01 g59314 ( .a(n_1723), .b(n_1090), .o(n_1799) );
AND2_X1 g58367 ( .a(n_2656), .b(n_2155), .o(n_2704) );
BUF_X2 newInst_1646 ( .a(newNet_1295), .o(newNet_1646) );
BUF_X2 newInst_1375 ( .a(newNet_1374), .o(newNet_1375) );
NAND3_Z1 g59488 ( .a(n_1243), .b(n_1558), .c(n_1094), .o(n_1650) );
BUF_X2 newInst_1016 ( .a(newNet_1015), .o(newNet_1016) );
NAND2_Z01 g60575 ( .a(n_372), .b(pX_12_), .o(n_536) );
NAND2_Z01 g34099 ( .a(n_4365), .b(n_4364), .o(n_4441) );
fflopd GPR_reg_8__5_ ( .CK(newNet_699), .D(n_2997), .Q(GPR_8__5_) );
NOR2_Z1 g59937 ( .a(n_1108), .b(n_44), .o(n_1187) );
XOR2_X1 g35101 ( .a(n_3463), .b(pX_5_), .o(n_4569) );
BUF_X2 newInst_1466 ( .a(newNet_1465), .o(newNet_1466) );
BUF_X2 newInst_109 ( .a(newNet_108), .o(newNet_109) );
NAND2_Z01 g60442 ( .a(n_358), .b(GPR_2__1_), .o(n_704) );
BUF_X2 newInst_336 ( .a(newNet_11), .o(newNet_336) );
NAND2_Z01 g59141 ( .a(n_1894), .b(n_51), .o(n_1958) );
AND2_X1 g34514 ( .a(n_3975), .b(n_3974), .o(n_4031) );
NAND2_Z01 g58459 ( .a(n_2599), .b(n_2183), .o(n_2637) );
AND2_X1 g57738 ( .a(n_3115), .b(n_2213), .o(n_3134) );
BUF_X2 newInst_408 ( .a(newNet_407), .o(newNet_408) );
NAND2_Z01 g60205 ( .a(n_578), .b(GPR_19__7_), .o(n_940) );
NAND2_Z01 g58726 ( .a(n_2207), .b(GPR_22__7_), .o(n_2381) );
NOR2_Z1 g34924 ( .a(n_3559), .b(n_3473), .o(n_3641) );
NAND2_Z01 g58598 ( .a(n_2458), .b(pX_9_), .o(n_2497) );
XOR2_X1 g59734 ( .a(n_1309), .b(n_90), .o(n_1396) );
NAND2_Z01 g59930 ( .a(n_1079), .b(n_212), .o(n_1216) );
NOR2_Z1 g59520 ( .a(n_1551), .b(n_367), .o(n_1621) );
BUF_X2 newInst_243 ( .a(newNet_242), .o(newNet_243) );
NOR2_Z2 g60352 ( .a(n_565), .b(rst), .o(n_856) );
BUF_X2 newInst_902 ( .a(newNet_901), .o(newNet_902) );
AND2_X1 g34505 ( .a(n_4013), .b(state_0_), .o(n_4036) );
NAND2_Z01 g59647 ( .a(io_do_7), .b(n_1418), .o(n_1474) );
BUF_X2 newInst_1471 ( .a(newNet_1470), .o(newNet_1471) );
NAND2_Z01 g60567 ( .a(n_341), .b(pY_2_), .o(n_542) );
BUF_X2 newInst_1473 ( .a(newNet_1472), .o(newNet_1473) );
NAND2_Z01 g57980 ( .a(n_2942), .b(n_2217), .o(n_2992) );
NAND2_Z01 g60470 ( .a(n_472), .b(n_255), .o(n_676) );
NOR2_Z1 g60347 ( .a(n_515), .b(n_525), .o(n_784) );
NOR2_Z1 g60811 ( .a(n_182), .b(n_160), .o(n_358) );
NAND2_Z01 g57944 ( .a(n_2963), .b(n_2314), .o(n_2998) );
BUF_X2 newInst_1242 ( .a(newNet_1241), .o(newNet_1242) );
NAND2_Z01 g59368 ( .a(n_1038), .b(n_1732), .o(n_1746) );
NAND2_Z01 g59008 ( .a(n_1922), .b(io_do_6), .o(n_2100) );
NAND2_Z01 g60303 ( .a(n_570), .b(pZ_7_), .o(n_821) );
NAND2_Z01 g60190 ( .a(n_644), .b(n_742), .o(n_955) );
fflopd SP_reg_15_ ( .CK(newNet_534), .D(n_2075), .Q(SP_15_) );
AND4_X1 g34127 ( .a(n_4263), .b(n_4303), .c(n_4304), .d(n_4111), .o(dmem_a_3) );
BUF_X2 newInst_490 ( .a(newNet_420), .o(newNet_490) );
AND2_X1 g60978 ( .a(n_4450), .b(n_4434), .o(n_190) );
fflopd pZ_reg_4_ ( .CK(newNet_76), .D(n_3025), .Q(pZ_4_) );
BUF_X2 newInst_323 ( .a(newNet_259), .o(newNet_323) );
NAND4_Z1 g58064 ( .a(n_1584), .b(n_2793), .c(n_2488), .d(n_2072), .o(n_2920) );
INV_X1 g61049 ( .a(pY_5_), .o(n_103) );
NOR2_Z1 g61022 ( .a(pmem_d_9), .b(pmem_d_1), .o(n_163) );
NAND2_Z01 g57843 ( .a(n_3033), .b(n_2313), .o(n_3067) );
NOR4_Z1 g58657 ( .a(n_1305), .b(n_2178), .c(n_1464), .d(n_1187), .o(n_2445) );
NAND2_Z01 g59839 ( .a(n_1135), .b(n_227), .o(n_1287) );
NAND2_Z01 g59923 ( .a(n_1027), .b(n_4649), .o(n_1218) );
NAND2_Z01 g59706 ( .a(io_do_7), .b(n_1353), .o(n_1424) );
NAND2_Z01 g34780 ( .a(n_3582), .b(GPR_0__3_), .o(n_3785) );
AND2_X1 g57996 ( .a(n_2940), .b(n_2212), .o(n_2975) );
AND2_X1 g60981 ( .a(PC_7_), .b(pmem_d_7), .o(n_187) );
NAND2_Z01 g57924 ( .a(n_2983), .b(n_2268), .o(n_3021) );
NAND2_Z01 g57932 ( .a(n_2975), .b(n_2425), .o(n_3013) );
fflopd GPR_reg_23__0_ ( .CK(newNet_1063), .D(n_2626), .Q(GPR_23__0_) );
INV_X1 drc_bufs35573 ( .a(n_3196), .o(n_3197) );
BUF_X2 newInst_397 ( .a(newNet_396), .o(newNet_397) );
BUF_X2 newInst_1140 ( .a(newNet_1139), .o(newNet_1140) );
NAND3_Z1 g60103 ( .a(n_682), .b(n_693), .c(n_634), .o(n_1017) );
fflopd GPR_reg_7__6_ ( .CK(newNet_748), .D(n_3067), .Q(GPR_7__6_) );
NAND2_Z01 g58884 ( .a(n_2140), .b(GPR_9__0_), .o(n_2223) );
NAND2_Z01 g35434 ( .a(n_3231), .b(pmem_d_0), .o(n_3286) );
BUF_X2 newInst_1582 ( .a(newNet_1581), .o(newNet_1582) );
INV_X1 g61053 ( .a(pX_14_), .o(n_99) );
NAND4_Z1 g59982 ( .a(n_491), .b(n_784), .c(n_762), .d(n_488), .o(n_1146) );
BUF_X2 newInst_1436 ( .a(newNet_1435), .o(newNet_1436) );
fflopd GPR_reg_22__0_ ( .CK(newNet_1108), .D(n_2627), .Q(GPR_22__0_) );
AND2_X1 g58501 ( .a(n_2567), .b(n_2156), .o(n_2596) );
NAND4_Z1 g57913 ( .a(n_2066), .b(n_2547), .c(n_2992), .d(n_2036), .o(n_3026) );
BUF_X2 newInst_676 ( .a(newNet_5), .o(newNet_676) );
NAND2_Z01 g60793 ( .a(n_194), .b(n_267), .o(n_316) );
BUF_X2 newInst_1760 ( .a(newNet_1759), .o(newNet_1760) );
AND2_X1 g58108 ( .a(n_2850), .b(n_2155), .o(n_2904) );
NAND2_Z01 g57717 ( .a(n_3123), .b(n_2337), .o(n_3150) );
fflopd GPR_reg_14__7_ ( .CK(newNet_1535), .D(n_3165), .Q(GPR_14__7_) );
NAND2_Z01 g34851 ( .a(n_3572), .b(GPR_4__0_), .o(n_3712) );
XOR2_X1 g60829 ( .a(PC_1_), .b(pmem_d_1), .o(n_302) );
fflopd U_reg_4_ ( .CK(newNet_377), .D(n_3022), .Q(U_4_) );
AND2_X1 g58252 ( .a(n_2752), .b(n_2158), .o(n_2815) );
NAND2_Z01 g34712 ( .a(n_3599), .b(GPR_5__6_), .o(n_3853) );
BUF_X2 newInst_254 ( .a(newNet_253), .o(newNet_254) );
BUF_X2 newInst_1001 ( .a(newNet_1000), .o(newNet_1001) );
BUF_X2 newInst_1806 ( .a(newNet_1805), .o(newNet_1806) );
BUF_X2 newInst_1249 ( .a(newNet_1248), .o(newNet_1249) );
BUF_X2 newInst_1529 ( .a(newNet_1528), .o(newNet_1529) );
fflopd pY_reg_2_ ( .CK(newNet_157), .D(n_2877), .Q(pY_2_) );
BUF_X2 newInst_950 ( .a(newNet_949), .o(newNet_950) );
BUF_X2 newInst_800 ( .a(newNet_799), .o(newNet_800) );
NAND2_Z01 g58869 ( .a(n_2139), .b(GPR_11__3_), .o(n_2238) );
BUF_X2 newInst_1790 ( .a(newNet_1789), .o(newNet_1790) );
NAND2_Z01 g60693 ( .a(U_9_), .b(n_249), .o(n_445) );
NAND2_Z01 g59107 ( .a(n_1875), .b(pX_14_), .o(n_2002) );
NAND2_Z01 g34789 ( .a(n_3629), .b(GPR_3__3_), .o(n_3776) );
NAND2_Z01 g60651 ( .a(n_334), .b(n_184), .o(n_490) );
NAND2_Z01 g60105 ( .a(n_847), .b(n_98), .o(n_1047) );
INV_X2 g59861 ( .a(n_1269), .o(n_1268) );
fflopd GPR_reg_3__3_ ( .CK(newNet_953), .D(n_2845), .Q(GPR_3__3_) );
NAND2_Z01 g59609 ( .a(n_1392), .b(n_4664), .o(n_1529) );
NAND2_Z02 g34362 ( .a(n_3209), .b(n_4075), .o(n_4178) );
BUF_X2 newInst_354 ( .a(newNet_167), .o(newNet_354) );
BUF_X2 newInst_533 ( .a(newNet_532), .o(newNet_533) );
NOR2_Z1 g34326 ( .a(n_16064_BAR), .b(n_3475), .o(n_4208) );
NAND2_Z01 g35418 ( .a(pZ_0_), .b(pmem_d_0), .o(n_3300) );
NAND2_Z01 g35208 ( .a(n_3412), .b(state_2_), .o(n_3440) );
AND2_X1 g35446 ( .a(state_3_), .b(state_0_), .o(n_4560) );
INV_X1 g60876 ( .a(n_248), .o(n_247) );
NAND2_Z01 g34986 ( .a(n_3549), .b(n_3461), .o(n_3596) );
NAND4_Z1 g34071 ( .a(n_4204), .b(n_4391), .c(n_4385), .d(n_4205), .o(dmem_do_1) );
BUF_X2 newInst_1047 ( .a(newNet_1046), .o(newNet_1047) );
NAND2_Z01 g59626 ( .a(n_1414), .b(io_di_6), .o(n_1501) );
NAND2_Z01 g58815 ( .a(n_2219), .b(n_1774), .o(n_2286) );
INV_X1 g60533 ( .a(n_602), .o(n_603) );
NAND2_Z01 g57831 ( .a(n_3045), .b(n_2424), .o(n_3082) );
AND2_X1 final_adder_mux_R16_278_6_g446 ( .a(n_4442), .b(n_4426), .o(final_adder_mux_R16_278_6_n_3) );
BUF_X2 newInst_1626 ( .a(newNet_1625), .o(newNet_1626) );
NAND2_Z01 g58848 ( .a(n_2158), .b(GPR_12__1_), .o(n_2259) );
NAND2_Z01 g60509 ( .a(Rd_4_), .b(n_345), .o(n_637) );
NOR2_Z1 g59761 ( .a(n_1268), .b(n_178), .o(n_1364) );
BUF_X2 newInst_1596 ( .a(newNet_1595), .o(newNet_1596) );
BUF_X2 newInst_1210 ( .a(newNet_440), .o(newNet_1210) );
BUF_X2 newInst_386 ( .a(newNet_385), .o(newNet_386) );
NAND2_Z01 g59875 ( .a(n_1164), .b(n_64), .o(n_1252) );
XOR2_X1 g35196 ( .a(n_3349), .b(n_3212), .o(n_4594) );
NAND2_Z01 g60841 ( .a(n_174), .b(n_273), .o(n_295) );
BUF_X2 newInst_1332 ( .a(newNet_1331), .o(newNet_1332) );
BUF_X2 newInst_525 ( .a(newNet_246), .o(newNet_525) );
BUF_X2 newInst_1743 ( .a(newNet_1406), .o(newNet_1743) );
BUF_X2 newInst_266 ( .a(newNet_265), .o(newNet_266) );
NAND2_Z01 g59161 ( .a(n_852), .b(n_1878), .o(n_1939) );
INV_Z1 g16801 ( .a(n_4467), .o(n_4413) );
fflopd GPR_reg_16__7_ ( .CK(newNet_1423), .D(n_3163), .Q(GPR_16__7_) );
BUF_X2 newInst_515 ( .a(newNet_437), .o(newNet_515) );
NOR2_Z1 g59872 ( .a(n_1219), .b(n_365), .o(n_1255) );
NAND2_Z01 g59853 ( .a(n_1016), .b(n_1173), .o(n_1275) );
NAND3_Z1 g59197 ( .a(n_1762), .b(n_1891), .c(n_1645), .o(n_1912) );
BUF_X2 newInst_916 ( .a(newNet_915), .o(newNet_916) );
BUF_X2 newInst_773 ( .a(newNet_772), .o(newNet_773) );
NAND2_Z01 g60319 ( .a(n_577), .b(pZ_8_), .o(n_807) );
BUF_X2 newInst_112 ( .a(newNet_22), .o(newNet_112) );
BUF_X2 newInst_1218 ( .a(newNet_1217), .o(newNet_1218) );
XOR2_X1 g35052 ( .a(n_3512), .b(PC_7_), .o(n_4541) );
BUF_X2 newInst_884 ( .a(newNet_883), .o(newNet_884) );
NAND2_Z01 g60422 ( .a(n_380), .b(GPR_6__4_), .o(n_724) );
fflopd GPR_reg_6__1_ ( .CK(newNet_824), .D(n_2742), .Q(GPR_6__1_) );
BUF_X2 newInst_730 ( .a(newNet_312), .o(newNet_730) );
XOR2_X1 g60863 ( .a(n_4449), .b(n_4433), .o(n_327) );
NAND2_Z01 g58895 ( .a(n_2139), .b(GPR_11__1_), .o(n_2187) );
XOR2_X1 g59810 ( .a(n_1199), .b(io_do_7), .o(n_1345) );
NAND2_Z01 g35122 ( .a(n_3469), .b(n_3461), .o(n_3490) );
INV_Z1 g16806 ( .a(GPR_21__1_), .o(n_4401) );
BUF_X2 newInst_240 ( .a(newNet_239), .o(newNet_240) );
NOR2_Z1 g34757 ( .a(n_3576), .b(n_4405), .o(n_3808) );
BUF_X2 newInst_1098 ( .a(newNet_1097), .o(newNet_1098) );
BUF_X2 newInst_819 ( .a(newNet_818), .o(newNet_819) );
NAND2_Z01 g58781 ( .a(n_2200), .b(GPR_7__1_), .o(n_2319) );
NAND2_Z01 g34834 ( .a(n_3587), .b(GPR_2__1_), .o(n_3729) );
BUF_X2 newInst_416 ( .a(newNet_31), .o(newNet_416) );
BUF_X2 newInst_22 ( .a(newNet_21), .o(newNet_22) );
NAND2_Z01 g35296 ( .a(n_3299), .b(pX_1_), .o(n_3379) );
NAND3_Z1 g35069 ( .a(n_3447), .b(n_3487), .c(n_3357), .o(n_3518) );
NAND2_Z01 g58834 ( .a(n_2159), .b(GPR_10__0_), .o(n_2273) );
NOR3_Z1 g59727 ( .a(n_1224), .b(n_161), .c(io_sel_0_), .o(n_1415) );
BUF_X2 newInst_1765 ( .a(newNet_1764), .o(newNet_1765) );
NAND2_Z01 g58147 ( .a(n_2819), .b(n_2289), .o(n_2866) );
BUF_X2 newInst_455 ( .a(newNet_37), .o(newNet_455) );
NAND4_Z1 g57814 ( .a(n_1927), .b(n_2520), .c(n_3054), .d(n_1928), .o(n_3093) );
NAND2_Z01 g58846 ( .a(n_2155), .b(GPR_14__0_), .o(n_2261) );
NAND2_Z01 g59010 ( .a(n_1993), .b(n_1593), .o(n_2098) );
NAND2_Z01 g59324 ( .a(n_1700), .b(n_4543), .o(n_1789) );
NAND2_Z01 g60925 ( .a(pmem_d_11), .b(pmem_d_10), .o(n_260) );
NAND2_Z01 g34192 ( .a(n_4325), .b(n_4468), .o(n_4331) );
NOR4_Z1 g58522 ( .a(n_2474), .b(n_2535), .c(n_2102), .d(n_1693), .o(n_2575) );
fflopd H_reg ( .CK(newNet_665), .D(n_0), .Q(H) );
NAND2_Z01 g35043 ( .a(n_4520), .b(n_4519), .o(n_3538) );
NAND2_Z02 g58956 ( .a(n_2088), .b(n_1215), .o(n_2159) );
NAND2_Z01 g58306 ( .a(n_2691), .b(n_2402), .o(n_2764) );
AND2_X1 g59288 ( .a(n_853), .b(n_1804), .o(n_1821) );
NAND2_Z01 g58641 ( .a(n_2358), .b(pZ_4_), .o(n_2455) );
BUF_X2 newInst_119 ( .a(newNet_118), .o(newNet_119) );
BUF_X2 newInst_672 ( .a(newNet_671), .o(newNet_672) );
XNOR2_X1 g59046 ( .a(n_1899), .b(n_1768), .o(n_2063) );
NAND2_Z01 g60245 ( .a(n_591), .b(GPR_22__0_), .o(n_900) );
AND2_X1 g59287 ( .a(n_1039), .b(n_1800), .o(n_1822) );
NAND2_Z01 g59067 ( .a(n_1896), .b(n_4514), .o(n_2040) );
NOR2_Z1 g35060 ( .a(n_3508), .b(pZ_7_), .o(n_4520) );
NAND2_Z01 g57722 ( .a(n_3118), .b(n_2189), .o(n_3145) );
BUF_X2 newInst_446 ( .a(newNet_445), .o(newNet_446) );
NOR2_Z1 g34418 ( .a(n_4043), .b(n_4088), .o(n_4119) );
INV_X1 g59126 ( .a(n_1973), .o(n_1974) );
NOR2_Z1 g34602 ( .a(n_3790), .b(n_3789), .o(n_3957) );
INV_X1 g35490 ( .a(pY_11_), .o(n_3235) );
BUF_X2 newInst_349 ( .a(newNet_10), .o(newNet_349) );
INV_X2 newInst_46 ( .a(newNet_45), .o(newNet_46) );
NAND2_Z01 g60401 ( .a(n_403), .b(n_418), .o(n_745) );
BUF_X2 newInst_1396 ( .a(newNet_1395), .o(newNet_1396) );
AND3_X1 g59204 ( .a(n_607), .b(n_1874), .c(pX_14_), .o(n_1968) );
NAND4_Z1 g34196 ( .a(n_4226), .b(n_4224), .c(n_4306), .d(n_4122), .o(n_4327) );
BUF_X2 newInst_219 ( .a(newNet_218), .o(newNet_219) );
INV_Z1 g16808 ( .a(GPR_12__1_), .o(n_4406) );
AND2_X1 g60333 ( .a(n_589), .b(n_36), .o(n_796) );
INV_X1 g35497 ( .a(pZ_1_), .o(n_3230) );
BUF_X2 newInst_126 ( .a(newNet_125), .o(newNet_126) );
NAND2_Z01 g60320 ( .a(n_614), .b(pX_4_), .o(n_864) );
AND2_X1 g58508 ( .a(n_2567), .b(n_2208), .o(n_2589) );
NAND2_Z01 g34333 ( .a(n_4158), .b(n_3556), .o(n_4201) );
BUF_X2 newInst_1565 ( .a(newNet_1153), .o(newNet_1565) );
BUF_X2 newInst_820 ( .a(newNet_449), .o(newNet_820) );
AND2_X1 g58965 ( .a(n_2086), .b(n_1212), .o(n_2141) );
NAND2_Z01 g60043 ( .a(n_4601), .b(n_856), .o(n_1087) );
NOR2_Z1 g59574 ( .a(n_1484), .b(SP_11_), .o(n_1568) );
NAND2_Z01 g34545 ( .a(n_3919), .b(n_3914), .o(pmem_a_7) );
BUF_X2 newInst_1788 ( .a(newNet_1787), .o(newNet_1788) );
BUF_X2 newInst_1310 ( .a(newNet_893), .o(newNet_1310) );
XOR2_X1 g59380 ( .a(n_1629), .b(pmem_d_6), .o(n_1738) );
fflopd GPR_reg_10__4_ ( .CK(newNet_1737), .D(n_2949), .Q(GPR_10__4_) );
AND2_X1 g59423 ( .a(n_1668), .b(n_1040), .o(n_1701) );
BUF_X2 newInst_130 ( .a(newNet_129), .o(newNet_130) );
AND2_X1 g60058 ( .a(n_845), .b(n_32), .o(n_1076) );
fflopd pX_reg_4_ ( .CK(newNet_225), .D(n_3029), .Q(pX_4_) );
BUF_X2 newInst_1346 ( .a(newNet_712), .o(newNet_1346) );
NAND2_Z01 g34689 ( .a(n_3631), .b(GPR_11__3_), .o(n_3876) );
BUF_X2 newInst_1062 ( .a(newNet_1061), .o(newNet_1062) );
BUF_X2 newInst_174 ( .a(newNet_173), .o(newNet_174) );
INV_X1 g34936 ( .a(n_3624), .o(n_3625) );
INV_X1 g59577 ( .a(n_1550), .o(n_1551) );
XOR2_X1 g35367 ( .a(pZ_1_), .b(pmem_d_1), .o(n_3322) );
BUF_X2 newInst_271 ( .a(newNet_270), .o(newNet_271) );
BUF_X2 newInst_1188 ( .a(newNet_466), .o(newNet_1188) );
NAND2_Z01 g60295 ( .a(n_746), .b(n_201), .o(n_829) );
BUF_X2 newInst_284 ( .a(newNet_283), .o(newNet_284) );
fflopd GPR_reg_2__4_ ( .CK(newNet_992), .D(n_2930), .Q(GPR_2__4_) );
NOR2_Z1 g35360 ( .a(n_3311), .b(n_3302), .o(n_4658) );
INV_X1 g35473 ( .a(pmem_d_6), .o(n_3251) );
NAND4_Z1 g58140 ( .a(n_1934), .b(n_2456), .c(n_2833), .d(n_2021), .o(n_2873) );
BUF_X2 newInst_882 ( .a(newNet_881), .o(newNet_882) );
NAND2_Z01 g34947 ( .a(n_3551), .b(GPR_13__6_), .o(n_3615) );
NAND2_Z01 g58879 ( .a(n_2153), .b(GPR_8__5_), .o(n_2228) );
NAND2_Z01 g34606 ( .a(n_3735), .b(n_3734), .o(n_3954) );
NAND3_Z1 g59446 ( .a(n_1609), .b(n_1417), .c(n_313), .o(n_1676) );
NOR2_Z1 g59826 ( .a(n_1194), .b(n_4472), .o(n_1298) );
fflopd PC_reg_1_ ( .CK(newNet_649), .D(n_2173), .Q(PC_1_) );
BUF_X2 newInst_1695 ( .a(newNet_1694), .o(newNet_1695) );
NOR2_Z1 g59007 ( .a(n_1970), .b(n_121), .o(n_2101) );
BUF_X2 newInst_407 ( .a(newNet_406), .o(newNet_407) );
BUF_X2 newInst_1487 ( .a(newNet_1469), .o(newNet_1487) );
INV_X1 g60953 ( .a(n_183), .o(n_182) );
NAND2_X2 g58931 ( .a(n_2128), .b(n_2083), .o(n_2194) );
NAND2_Z01 g60514 ( .a(n_370), .b(GPR_20__6_), .o(n_632) );
NAND4_Z1 g34594 ( .a(n_3705), .b(n_3706), .c(n_3708), .d(n_3707), .o(n_3966) );
NAND2_Z01 g35289 ( .a(n_3299), .b(pX_4_), .o(n_3386) );
NAND2_Z01 g59463 ( .a(n_1041), .b(n_1615), .o(n_1658) );
NAND2_Z01 g59915 ( .a(n_1068), .b(n_961), .o(n_1197) );
NOR2_Z1 g60684 ( .a(n_33), .b(n_256), .o(n_470) );
NAND2_Z01 g34263 ( .a(n_4176), .b(pX_1_), .o(n_4270) );
NAND2_Z01 g60244 ( .a(n_598), .b(GPR_15__3_), .o(n_901) );
NAND2_Z01 g34953 ( .a(n_3551), .b(GPR_7__4_), .o(n_3609) );
NOR3_Z1 g60128 ( .a(n_44), .b(n_601), .c(pmem_d_3), .o(n_1033) );
NAND2_Z01 g34701 ( .a(n_3575), .b(GPR_8__6_), .o(n_3864) );
NAND2_Z01 g58673 ( .a(n_2214), .b(GPR_16__7_), .o(n_2433) );
INV_X2 newInst_187 ( .a(newNet_158), .o(newNet_187) );
INV_X1 g60279 ( .a(n_864), .o(n_865) );
NAND2_Z01 g59783 ( .a(n_1268), .b(n_479), .o(n_1341) );
BUF_X2 newInst_876 ( .a(newNet_875), .o(newNet_876) );
BUF_X2 newInst_536 ( .a(newNet_535), .o(newNet_536) );
NAND2_Z01 g58162 ( .a(n_2804), .b(n_2385), .o(n_2848) );
NAND4_Z1 g34074 ( .a(n_4276), .b(n_4300), .c(n_4381), .d(n_4140), .o(dmem_a_6) );
BUF_X2 newInst_85 ( .a(newNet_84), .o(newNet_85) );
INV_X1 g35108 ( .a(n_3492), .o(n_3491) );
NAND2_Z01 g35429 ( .a(n_3248), .b(pmem_d_10), .o(n_4633) );
BUF_X2 newInst_1554 ( .a(newNet_1553), .o(newNet_1554) );
NOR2_Z1 g58175 ( .a(n_2792), .b(n_587), .o(n_2837) );
fflopd GPR_reg_17__3_ ( .CK(newNet_1398), .D(n_2858), .Q(GPR_17__3_) );
NOR2_Z1 g35331 ( .a(n_3218), .b(n_3309), .o(n_3338) );
BUF_X2 newInst_1815 ( .a(newNet_1814), .o(newNet_1815) );
AND2_X1 g58396 ( .a(n_2656), .b(n_2202), .o(n_2672) );
NOR2_Z1 g59114 ( .a(n_1874), .b(n_106), .o(n_1995) );
BUF_X2 newInst_1181 ( .a(newNet_1180), .o(newNet_1181) );
NOR3_Z1 g59187 ( .a(n_1446), .b(n_1893), .c(n_77), .o(n_1920) );
NAND4_Z1 g34579 ( .a(n_3794), .b(n_3797), .c(n_3796), .d(n_3795), .o(n_3981) );
NAND2_Z01 g59142 ( .a(n_1894), .b(n_1455), .o(n_1957) );
NAND2_Z01 g58738 ( .a(n_2205), .b(GPR_2__3_), .o(n_2369) );
BUF_X2 newInst_1255 ( .a(newNet_1254), .o(newNet_1255) );
BUF_X2 newInst_718 ( .a(newNet_717), .o(newNet_718) );
BUF_X2 newInst_1388 ( .a(newNet_1387), .o(newNet_1388) );
BUF_X2 newInst_1714 ( .a(newNet_1713), .o(newNet_1714) );
BUF_X2 newInst_1407 ( .a(newNet_1406), .o(newNet_1407) );
BUF_X2 newInst_1115 ( .a(newNet_1114), .o(newNet_1115) );
NAND2_Z01 g58298 ( .a(n_2699), .b(n_2310), .o(n_2772) );
NAND2_Z01 g59687 ( .a(n_1389), .b(n_156), .o(n_1440) );
BUF_X2 newInst_472 ( .a(newNet_471), .o(newNet_472) );
NAND2_Z01 g60484 ( .a(n_20), .b(Rd_r_1_), .o(n_662) );
BUF_X2 newInst_1771 ( .a(newNet_1770), .o(newNet_1771) );
BUF_X2 newInst_320 ( .a(newNet_319), .o(newNet_320) );
NAND2_Z01 g59695 ( .a(io_do_1), .b(n_1384), .o(n_1435) );
NAND2_Z01 g34253 ( .a(n_4179), .b(SP_8_), .o(n_4280) );
NAND2_Z01 final_adder_mux_R16_278_6_g427 ( .a(n_4442), .b(n_4426), .o(final_adder_mux_R16_278_6_n_21) );
AND3_X1 g59594 ( .a(n_1041), .b(n_1450), .c(pmem_d_12), .o(n_1535) );
INV_X1 drc_bufs35591 ( .a(n_4125), .o(n_3209) );
INV_X1 g60949 ( .a(n_200), .o(n_199) );
NAND2_Z01 g60942 ( .a(io_do_2), .b(n_44), .o(n_209) );
NAND3_Z1 g34552 ( .a(n_3791), .b(n_3793), .c(n_3792), .o(n_4007) );
BUF_X2 newInst_592 ( .a(newNet_591), .o(newNet_592) );
BUF_X2 newInst_1719 ( .a(newNet_1718), .o(newNet_1719) );
BUF_X2 newInst_278 ( .a(newNet_277), .o(newNet_278) );
BUF_X2 newInst_1777 ( .a(newNet_1776), .o(newNet_1777) );
NAND2_Z01 g59558 ( .a(n_1516), .b(n_229), .o(n_1574) );
AND2_X1 final_adder_mux_R16_278_6_g447 ( .a(n_4443), .b(n_4427), .o(final_adder_mux_R16_278_6_n_2) );
NAND2_Z01 g57700 ( .a(n_3142), .b(n_2260), .o(n_3169) );
NOR3_Z1 g59805 ( .a(n_850), .b(n_1156), .c(io_do_1), .o(n_1323) );
NAND2_Z01 final_adder_mux_R16_278_6_g371 ( .a(final_adder_mux_R16_278_6_n_77), .b(final_adder_mux_R16_278_6_n_1), .o(final_adder_mux_R16_278_6_n_78) );
BUF_X2 newInst_910 ( .a(newNet_909), .o(newNet_910) );
BUF_X2 newInst_146 ( .a(newNet_145), .o(newNet_146) );
NAND2_Z01 g57709 ( .a(n_3132), .b(n_2414), .o(n_3160) );
NAND2_Z01 g58575 ( .a(n_2459), .b(n_2040), .o(n_2521) );
BUF_X2 newInst_784 ( .a(newNet_783), .o(newNet_784) );
BUF_X2 newInst_437 ( .a(newNet_436), .o(newNet_437) );
NAND2_Z01 g59137 ( .a(n_1872), .b(n_1318), .o(n_1961) );
NAND2_Z01 g60618 ( .a(n_66), .b(n_470), .o(n_589) );
NAND2_Z01 g35330 ( .a(pZ_9_), .b(n_3199), .o(n_3339) );
NAND2_Z01 g34629 ( .a(n_3645), .b(pZ_11_), .o(n_3931) );
NAND2_Z01 g60708 ( .a(U_13_), .b(n_249), .o(n_430) );
NAND2_Z01 g35255 ( .a(n_3328), .b(n_3220), .o(n_4485) );
INV_X1 g35516 ( .a(pY_3_), .o(n_3212) );
BUF_X2 newInst_1605 ( .a(newNet_1604), .o(newNet_1605) );
NAND4_Z1 g34457 ( .a(n_3882), .b(n_4001), .c(n_4053), .d(n_3888), .o(n_4085) );
BUF_X2 newInst_1316 ( .a(newNet_1315), .o(newNet_1316) );
NOR2_Z1 g60971 ( .a(n_4440), .b(n_4424), .o(n_151) );
AND2_X1 g60763 ( .a(n_160), .b(n_35), .o(n_460) );
AND2_X1 g59404 ( .a(n_39), .b(n_1664), .o(n_1712) );
INV_X1 drc_bufs61162 ( .a(n_571), .o(n_24) );
BUF_X2 newInst_848 ( .a(newNet_316), .o(newNet_848) );
NAND2_Z01 g59941 ( .a(n_1033), .b(pmem_d_1), .o(n_1207) );
NAND2_Z01 g58631 ( .a(n_2359), .b(n_2009), .o(n_2478) );
AND2_X1 g58123 ( .a(n_2850), .b(n_2202), .o(n_2889) );
AND2_X1 g35242 ( .a(n_4683), .b(pmem_d_13), .o(n_3418) );
NOR4_Z1 g59901 ( .a(n_998), .b(n_980), .c(n_993), .d(n_982), .o(n_1229) );
NAND4_Z1 g59552 ( .a(n_1473), .b(n_1437), .c(n_1493), .d(n_1050), .o(n_1576) );
BUF_X2 newInst_995 ( .a(newNet_994), .o(newNet_995) );
XOR2_X1 final_adder_mux_R16_278_6_g408 ( .a(n_4445), .b(n_4429), .o(final_adder_mux_R16_278_6_n_41) );
XOR2_X1 g60856 ( .a(PC_10_), .b(pmem_d_10), .o(n_288) );
AND2_X1 g35297 ( .a(n_3228), .b(n_3298), .o(n_3378) );
BUF_X2 newInst_1179 ( .a(newNet_571), .o(newNet_1179) );
AND3_X1 g59192 ( .a(n_611), .b(n_1870), .c(pZ_14_), .o(n_1973) );
XOR2_X1 g59675 ( .a(n_1348), .b(n_76), .o(n_1454) );
NAND2_Z01 g60199 ( .a(n_749), .b(n_22), .o(n_946) );
NAND3_Z1 g59447 ( .a(n_849), .b(n_1600), .c(n_64), .o(n_1675) );
NAND2_Z01 g59263 ( .a(n_1807), .b(n_194), .o(n_1847) );
NAND2_Z01 g35281 ( .a(U_15_), .b(n_3275), .o(n_3394) );
NAND2_Z01 g58241 ( .a(n_2756), .b(n_2215), .o(n_2826) );
AND2_X1 g61021 ( .a(SP_0_), .b(SP_1_), .o(n_164) );
AND2_X1 g60635 ( .a(n_369), .b(SP_2_), .o(n_499) );
NAND2_Z01 g60992 ( .a(n_71), .b(n_62), .o(n_142) );
NAND2_Z01 g58697 ( .a(n_2210), .b(GPR_1__4_), .o(n_2409) );
NAND2_Z01 g34471 ( .a(n_4647), .b(n_4025), .o(n_4072) );
NAND2_Z01 g60451 ( .a(n_370), .b(GPR_22__1_), .o(n_695) );
NAND2_Z01 g59320 ( .a(n_4), .b(n_4551), .o(n_1793) );
NAND2_Z01 g58329 ( .a(n_2664), .b(n_2221), .o(n_2736) );
NAND2_Z01 g35406 ( .a(pY_2_), .b(pmem_d_2), .o(n_3304) );
AND2_X1 g58263 ( .a(n_2752), .b(n_2207), .o(n_2804) );
NAND2_Z01 g59637 ( .a(n_1402), .b(io_do_1), .o(n_1492) );
NAND2_Z01 g59100 ( .a(n_1885), .b(n_1713), .o(n_2060) );
BUF_X2 newInst_757 ( .a(newNet_659), .o(newNet_757) );
BUF_X2 newInst_1093 ( .a(newNet_1092), .o(newNet_1093) );
NOR2_Z1 g34390 ( .a(n_4083), .b(n_3469), .o(n_4148) );
BUF_X2 newInst_1331 ( .a(newNet_1330), .o(newNet_1331) );
NAND2_Z01 g35308 ( .a(n_3289), .b(pY_1_), .o(n_3368) );
NAND2_Z01 g34768 ( .a(n_3625), .b(GPR_1__4_), .o(n_3797) );
INV_X1 g35321 ( .a(n_3351), .o(n_3350) );
BUF_X2 newInst_1265 ( .a(newNet_1264), .o(newNet_1265) );
NAND2_Z01 g59056 ( .a(n_1894), .b(n_4524), .o(n_2051) );
XOR2_X1 g34662 ( .a(n_3555), .b(pZ_4_), .o(n_3903) );
BUF_X2 newInst_324 ( .a(newNet_323), .o(newNet_324) );
NAND2_Z01 g60526 ( .a(n_368), .b(GPR_13__5_), .o(n_620) );
NAND2_Z01 g57828 ( .a(n_3048), .b(n_2241), .o(n_3085) );
NAND2_Z01 g59096 ( .a(n_1897), .b(n_262), .o(n_2012) );
NAND2_Z01 g58324 ( .a(n_2670), .b(n_2326), .o(n_2741) );
XNOR2_X1 g60868 ( .a(n_4445), .b(n_4429), .o(n_326) );
BUF_X2 newInst_1787 ( .a(newNet_1786), .o(newNet_1787) );
NAND2_Z01 g59829 ( .a(n_1142), .b(pmem_d_15), .o(n_1295) );
NAND2_Z01 g58292 ( .a(n_2704), .b(n_2234), .o(n_2778) );
NAND2_Z01 g34488 ( .a(n_4037), .b(n_3305), .o(n_4058) );
NAND2_Z01 g34727 ( .a(n_3599), .b(GPR_4__5_), .o(n_3838) );
NOR2_Z1 g35170 ( .a(n_3427), .b(pY_4_), .o(n_3462) );
fflopd U_reg_6_ ( .CK(newNet_366), .D(n_3110), .Q(U_6_) );
BUF_X2 newInst_1573 ( .a(newNet_1011), .o(newNet_1573) );
NAND2_Z01 g60747 ( .a(SP_9_), .b(n_180), .o(n_395) );
BUF_X2 newInst_1480 ( .a(newNet_271), .o(newNet_1480) );
NAND2_Z01 g60998 ( .a(n_119), .b(n_104), .o(n_175) );
NAND2_Z01 g59629 ( .a(n_1414), .b(io_di_7), .o(n_1498) );
fflopd GPR_reg_22__3_ ( .CK(newNet_1096), .D(n_2848), .Q(GPR_22__3_) );
BUF_X2 newInst_825 ( .a(newNet_753), .o(newNet_825) );
XOR2_X1 g60870 ( .a(n_4447), .b(n_4431), .o(n_323) );
BUF_X2 newInst_1640 ( .a(newNet_1639), .o(newNet_1640) );
NOR2_Z1 g60806 ( .a(n_134), .b(pmem_d_1), .o(n_312) );
NOR4_Z1 g59902 ( .a(n_990), .b(n_985), .c(n_1002), .d(n_997), .o(n_1228) );
NOR2_Z1 g59885 ( .a(n_1219), .b(n_459), .o(n_1242) );
NAND2_Z01 g59754 ( .a(n_1312), .b(io_do_2), .o(n_1370) );
NOR2_Z1 g34963 ( .a(n_3511), .b(n_3553), .o(n_3636) );
NAND2_Z01 g58551 ( .a(n_2496), .b(pY_10_), .o(n_2546) );
NAND2_Z01 g61007 ( .a(n_35), .b(n_62), .o(n_172) );
BUF_X2 newInst_1079 ( .a(newNet_1078), .o(newNet_1079) );
BUF_X2 newInst_963 ( .a(newNet_962), .o(newNet_963) );
XOR2_X1 g35145 ( .a(n_3451), .b(n_3325), .o(n_3472) );
NAND2_Z01 g58443 ( .a(n_2622), .b(n_2216), .o(n_2650) );
BUF_X2 newInst_1440 ( .a(newNet_1439), .o(newNet_1440) );
NAND2_Z01 g58234 ( .a(n_2754), .b(n_2218), .o(n_2833) );
NOR2_Z1 g34910 ( .a(n_3632), .b(n_3218), .o(n_3653) );
BUF_X2 newInst_162 ( .a(newNet_161), .o(newNet_162) );
NOR2_Z1 g59936 ( .a(n_1108), .b(n_62), .o(n_1188) );
BUF_X2 newInst_705 ( .a(newNet_704), .o(newNet_705) );
AND2_X1 g58357 ( .a(n_2656), .b(n_2159), .o(n_2714) );
BUF_X2 newInst_1526 ( .a(newNet_1525), .o(newNet_1526) );
BUF_X2 newInst_1416 ( .a(newNet_1415), .o(newNet_1416) );
NOR2_Z1 g34361 ( .a(n_4139), .b(n_3656), .o(n_4171) );
NAND2_Z01 g59916 ( .a(n_1039), .b(n_961), .o(n_1223) );
AND2_X1 g58604 ( .a(n_2444), .b(n_587), .o(n_2491) );
NAND4_Z1 g59666 ( .a(n_1155), .b(n_1265), .c(n_1419), .d(n_1024), .o(n_1462) );
NAND2_Z01 g58095 ( .a(n_2852), .b(n_2217), .o(n_2918) );
BUF_X2 newInst_936 ( .a(newNet_935), .o(newNet_936) );
BUF_X2 newInst_836 ( .a(newNet_835), .o(newNet_836) );
NAND2_Z01 g60963 ( .a(n_68), .b(pmem_d_3), .o(n_156) );
NAND2_Z01 g58303 ( .a(n_2694), .b(n_2412), .o(n_2767) );
NAND2_Z01 g34882 ( .a(n_3564), .b(pX_4_), .o(n_3681) );
AND2_X1 g58385 ( .a(n_2656), .b(n_2207), .o(n_2683) );
NAND2_Z01 g34892 ( .a(n_3633), .b(pZ_12_), .o(n_3671) );
BUF_X2 newInst_765 ( .a(newNet_764), .o(newNet_765) );
fflopd GPR_reg_5__5_ ( .CK(newNet_847), .D(n_3000), .Q(GPR_5__5_) );
AND2_X1 g59217 ( .a(n_1844), .b(SP_15_), .o(n_1888) );
NAND2_Z01 g58165 ( .a(n_2801), .b(n_2349), .o(n_2845) );
NAND2_Z01 g57986 ( .a(n_2941), .b(n_2198), .o(n_2986) );
fflopd GPR_reg_11__3_ ( .CK(newNet_1696), .D(n_2864), .Q(GPR_11__3_) );
NAND4_Z1 g34565 ( .a(n_3866), .b(n_3867), .c(n_3868), .d(n_3865), .o(n_3995) );
NAND2_Z01 g58687 ( .a(n_2211), .b(GPR_19__3_), .o(n_2419) );
BUF_X2 newInst_289 ( .a(newNet_288), .o(newNet_289) );
BUF_X2 newInst_580 ( .a(newNet_579), .o(newNet_580) );
NAND2_Z01 g58883 ( .a(n_2153), .b(GPR_8__7_), .o(n_2224) );
NOR2_Z1 g34300 ( .a(n_4155), .b(n_4159), .o(n_4234) );
INV_X1 g59237 ( .a(n_1869), .o(n_1868) );
BUF_X2 newInst_1046 ( .a(newNet_1004), .o(newNet_1046) );
NOR2_Z1 g35443 ( .a(pmem_d_11), .b(pmem_d_10), .o(n_4659) );
BUF_X2 newInst_1621 ( .a(newNet_1620), .o(newNet_1621) );
BUF_X2 newInst_694 ( .a(newNet_693), .o(newNet_694) );
NAND2_Z01 g61001 ( .a(n_122), .b(n_65), .o(n_138) );
NOR2_Z1 g60113 ( .a(n_855), .b(n_4609), .o(n_1013) );
NAND2_Z01 g34205 ( .a(io_do_2), .b(n_4177), .o(n_4321) );
AND2_X1 g57997 ( .a(n_2940), .b(n_2211), .o(n_2974) );
NAND2_Z01 g35274 ( .a(n_3289), .b(pY_14_), .o(n_3401) );
NAND2_Z01 g35218 ( .a(n_4559), .b(state_2_), .o(n_3448) );
NAND2_Z01 g60031 ( .a(n_846), .b(pmem_d_14), .o(n_1098) );
XOR2_X1 g34481 ( .a(n_4040), .b(SP_1_), .o(n_4061) );
BUF_X2 newInst_659 ( .a(newNet_658), .o(newNet_659) );
BUF_X2 newInst_420 ( .a(newNet_419), .o(newNet_420) );
BUF_X2 newInst_208 ( .a(newNet_25), .o(newNet_208) );
BUF_X2 newInst_52 ( .a(newNet_51), .o(newNet_52) );
BUF_X2 newInst_1417 ( .a(newNet_1416), .o(newNet_1417) );
AND2_X1 g58272 ( .a(n_2752), .b(n_2140), .o(n_2795) );
BUF_X2 newInst_895 ( .a(newNet_894), .o(newNet_895) );
BUF_X2 newInst_1442 ( .a(newNet_544), .o(newNet_1442) );
BUF_X2 newInst_575 ( .a(newNet_496), .o(newNet_575) );
NAND4_Z1 g34584 ( .a(n_3757), .b(n_3758), .c(n_3759), .d(n_3760), .o(n_3976) );
NAND2_Z01 g60340 ( .a(n_487), .b(pmem_d_3), .o(n_790) );
BUF_X2 newInst_927 ( .a(newNet_926), .o(newNet_927) );
BUF_X2 newInst_367 ( .a(newNet_325), .o(newNet_367) );
NOR2_Z1 g61000 ( .a(PC_1_), .b(pmem_d_4), .o(n_173) );
NOR2_Z1 g60647 ( .a(n_324), .b(n_188), .o(n_493) );
NOR2_Z1 g60614 ( .a(n_469), .b(n_260), .o(n_510) );
NAND2_Z01 g34872 ( .a(n_3575), .b(GPR_8__7_), .o(n_3691) );
NAND2_Z01 g59705 ( .a(io_do_6), .b(n_1384), .o(n_1425) );
NOR2_Z1 g34447 ( .a(n_4069), .b(n_3930), .o(n_4093) );
BUF_X2 newInst_1513 ( .a(newNet_1512), .o(newNet_1513) );
fflopd state_reg_1_ ( .CK(newNet_26), .D(n_2910), .Q(state_1_) );
NOR4_Z1 g34213 ( .a(n_3979), .b(n_3980), .c(n_4289), .d(n_3956), .o(n_4313) );
NAND2_Z01 g60969 ( .a(n_38), .b(pmem_d_1), .o(n_196) );
INV_X2 g61093 ( .a(pmem_d_9), .o(n_59) );
NOR2_Z1 g60744 ( .a(n_279), .b(n_115), .o(n_466) );
AND2_X1 g58006 ( .a(n_2940), .b(n_2202), .o(n_2965) );
BUF_X2 newInst_76 ( .a(newNet_75), .o(newNet_76) );
BUF_X2 newInst_1758 ( .a(newNet_1757), .o(newNet_1758) );
AND2_X1 g57906 ( .a(n_3009), .b(n_2153), .o(n_3032) );
NAND2_Z01 g34177 ( .a(n_4325), .b(n_4472), .o(n_4339) );
NAND2_Z01 g34282 ( .a(n_4162), .b(pY_5_), .o(n_4251) );
NAND2_Z01 g60473 ( .a(n_4530), .b(n_340), .o(n_673) );
BUF_X2 newInst_1232 ( .a(newNet_1231), .o(newNet_1232) );
NAND2_Z01 g60087 ( .a(n_857), .b(n_90), .o(n_1050) );
BUF_X2 newInst_45 ( .a(newNet_44), .o(newNet_45) );
NAND2_Z01 g58049 ( .a(n_2896), .b(n_2392), .o(n_2933) );
INV_X2 newInst_1456 ( .a(newNet_1455), .o(newNet_1456) );
BUF_X2 newInst_646 ( .a(newNet_645), .o(newNet_646) );
NOR2_Z1 g58564 ( .a(n_2484), .b(n_579), .o(n_2534) );
NAND2_Z01 g35113 ( .a(n_3470), .b(PC_5_), .o(n_3493) );
NAND2_Z01 g34821 ( .a(n_3625), .b(GPR_1__2_), .o(n_3742) );
NOR2_Z1 g59971 ( .a(n_1042), .b(n_252), .o(n_1167) );
NAND2_Z01 g58628 ( .a(n_2286), .b(n_1778), .o(n_2482) );
NAND4_Z1 g34125 ( .a(n_4105), .b(n_4186), .c(n_4328), .d(n_4133), .o(dmem_a_0) );
NOR2_Z1 g35211 ( .a(n_3365), .b(n_3343), .o(n_3439) );
BUF_X2 newInst_335 ( .a(newNet_149), .o(newNet_335) );
BUF_X2 newInst_920 ( .a(newNet_795), .o(newNet_920) );
NOR2_Z1 g59770 ( .a(n_1307), .b(pmem_d_6), .o(n_1358) );
AND2_X1 g58118 ( .a(n_2850), .b(n_2206), .o(n_2894) );
fflopd GPR_reg_4__6_ ( .CK(newNet_899), .D(n_3070), .Q(GPR_4__6_) );
BUF_X2 newInst_978 ( .a(newNet_892), .o(newNet_978) );
NOR2_Z1 g59948 ( .a(n_1117), .b(n_969), .o(n_1204) );
NAND2_Z01 g59065 ( .a(n_1902), .b(n_4588), .o(n_2042) );
NAND2_Z01 g60408 ( .a(n_349), .b(U_7_), .o(n_738) );
NOR2_Z1 g34301 ( .a(n_4081), .b(n_4159), .o(n_4233) );
fflopd GPR_reg_12__7_ ( .CK(newNet_1619), .D(n_3167), .Q(GPR_12__7_) );
NAND2_Z01 g34972 ( .a(n_3552), .b(n_3461), .o(n_3624) );
BUF_X2 newInst_302 ( .a(newNet_301), .o(newNet_302) );
NAND2_Z01 g34747 ( .a(n_3629), .b(GPR_3__5_), .o(n_3818) );
BUF_X2 newInst_865 ( .a(newNet_864), .o(newNet_865) );
NAND2_Z01 g58334 ( .a(n_2689), .b(n_835), .o(n_2755) );
NAND2_Z01 g58795 ( .a(n_2199), .b(GPR_0__5_), .o(n_2305) );
NAND2_Z01 g60936 ( .a(pmem_d_1), .b(pmem_d_0), .o(n_252) );
INV_X1 g59233 ( .a(n_1878), .o(n_1877) );
BUF_X2 newInst_603 ( .a(newNet_230), .o(newNet_603) );
BUF_X2 newInst_56 ( .a(newNet_55), .o(newNet_56) );
INV_X1 g35319 ( .a(n_3353), .o(n_3354) );
NAND2_Z01 g60238 ( .a(n_584), .b(GPR_18__2_), .o(n_907) );
BUF_X2 newInst_1795 ( .a(newNet_1794), .o(newNet_1795) );
NAND2_Z01 g60563 ( .a(n_349), .b(pX_4_), .o(n_545) );
NAND2_Z01 g59840 ( .a(n_1138), .b(n_226), .o(n_1286) );
AND2_X1 g58257 ( .a(n_2752), .b(n_2213), .o(n_2810) );
NOR2_Z1 g60097 ( .a(n_4556), .b(n_860), .o(n_1022) );
INV_X1 g35151 ( .a(n_4641), .o(n_3460) );
NAND2_Z01 g58722 ( .a(n_2207), .b(GPR_22__3_), .o(n_2385) );
AND2_X1 g57885 ( .a(n_3009), .b(n_2159), .o(n_3053) );
INV_X1 g60287 ( .a(n_767), .o(n_838) );
NAND2_Z01 g60913 ( .a(PC_1_), .b(pmem_d_1), .o(n_228) );
NAND2_Z01 g35154 ( .a(n_3451), .b(n_3283), .o(n_3458) );
BUF_X2 newInst_609 ( .a(newNet_422), .o(newNet_609) );
INV_X1 drc_bufs61226 ( .a(n_1661), .o(n_29) );
fflopd pX_reg_14_ ( .CK(newNet_256), .D(n_3116), .Q(pX_14_) );
BUF_X2 newInst_1224 ( .a(newNet_1223), .o(newNet_1224) );
NAND2_Z01 g58056 ( .a(n_2888), .b(n_2324), .o(n_2926) );
NAND3_Z1 g59895 ( .a(io_do_4), .b(n_1026), .c(n_365), .o(n_1234) );
NAND2_Z01 g59393 ( .a(n_1648), .b(dmem_di_4), .o(n_1722) );
NAND2_Z01 g57824 ( .a(n_3052), .b(n_2262), .o(n_3089) );
NAND2_Z01 g34673 ( .a(n_3605), .b(n_3606), .o(n_3892) );
BUF_X2 newInst_814 ( .a(newNet_388), .o(newNet_814) );
AND2_X1 g58954 ( .a(n_2081), .b(pY_15_), .o(n_2146) );
BUF_X2 newInst_1834 ( .a(newNet_1833), .o(newNet_1834) );
XOR2_X1 g60669 ( .a(n_162), .b(io_do_2), .o(n_563) );
NAND2_Z01 g58858 ( .a(n_2157), .b(GPR_13__6_), .o(n_2249) );
XOR2_X1 g35102 ( .a(n_4624), .b(n_3231), .o(n_4468) );
BUF_X2 newInst_664 ( .a(newNet_1), .o(newNet_664) );
NAND2_Z01 g60471 ( .a(n_342), .b(GPR_17__3_), .o(n_675) );
fflopd GPR_reg_4__7_ ( .CK(newNet_888), .D(n_3150), .Q(GPR_4__7_) );
BUF_X2 newInst_796 ( .a(newNet_795), .o(newNet_796) );
BUF_X2 newInst_1206 ( .a(newNet_1205), .o(newNet_1206) );
BUF_X2 newInst_639 ( .a(newNet_638), .o(newNet_639) );
NAND2_Z01 g60826 ( .a(n_178), .b(n_93), .o(n_303) );
NAND2_Z01 g60276 ( .a(n_591), .b(GPR_22__5_), .o(n_870) );
INV_X1 g60677 ( .a(n_466), .o(n_465) );
BUF_X2 newInst_1692 ( .a(newNet_1691), .o(newNet_1692) );
BUF_X2 newInst_807 ( .a(newNet_806), .o(newNet_807) );
BUF_X2 newInst_1054 ( .a(newNet_1053), .o(newNet_1054) );
BUF_X2 newInst_1171 ( .a(newNet_780), .o(newNet_1171) );
BUF_X2 newInst_1669 ( .a(newNet_1668), .o(newNet_1669) );
NAND2_Z01 g59072 ( .a(n_1902), .b(n_4589), .o(n_2035) );
INV_X1 g35465 ( .a(pmem_d_8), .o(n_3259) );
NAND2_Z01 g34677 ( .a(n_3633), .b(pZ_15_), .o(n_3888) );
INV_X1 g35501 ( .a(pZ_12_), .o(n_3226) );
XOR2_X1 g34436 ( .a(n_4074), .b(pY_11_), .o(n_4103) );
NAND2_Z01 g34811 ( .a(n_3587), .b(GPR_2__2_), .o(n_3752) );
NAND2_Z01 g34762 ( .a(n_3572), .b(GPR_4__4_), .o(n_3803) );
NAND2_Z01 g60904 ( .a(PC_8_), .b(pmem_d_8), .o(n_267) );
NAND3_Z1 g60368 ( .a(n_4533), .b(n_608), .c(n_97), .o(n_773) );
NAND2_Z01 g58560 ( .a(n_2502), .b(pX_14_), .o(n_2538) );
fflopd GPR_reg_10__3_ ( .CK(newNet_1742), .D(n_2865), .Q(GPR_10__3_) );
BUF_X2 newInst_1533 ( .a(newNet_1532), .o(newNet_1533) );
NOR2_Z1 g60212 ( .a(n_581), .b(n_79), .o(n_933) );
fflopd GPR_reg_13__5_ ( .CK(newNet_1594), .D(n_3018), .Q(GPR_13__5_) );
NAND2_Z01 g59693 ( .a(io_do_0), .b(n_1353), .o(n_1437) );
NAND2_Z01 g34258 ( .a(n_4176), .b(pX_5_), .o(n_4275) );
AND2_X1 g59959 ( .a(n_1029), .b(pmem_d_7), .o(n_1173) );
NAND3_Z1 g59533 ( .a(n_1423), .b(n_1481), .c(n_1495), .o(n_1594) );
NOR2_Z1 g61018 ( .a(n_4557), .b(state_2_), .o(n_128) );
NOR2_Z1 g59952 ( .a(n_1001), .b(n_1053), .o(n_1178) );
AND2_X1 final_adder_mux_R16_278_6_g440 ( .a(n_4448), .b(n_4432), .o(final_adder_mux_R16_278_6_n_9) );
AND3_X1 g60377 ( .a(pmem_d_3), .b(n_346), .c(pmem_d_2), .o(n_839) );
AND2_X1 g58360 ( .a(n_2656), .b(n_2139), .o(n_2711) );
fflopd GPR_reg_20__5_ ( .CK(newNet_1187), .D(n_3007), .Q(GPR_20__5_) );
NAND2_Z01 g34138 ( .a(n_4317), .b(n_4617), .o(n_4370) );
INV_X2 newInst_1503 ( .a(newNet_300), .o(newNet_1503) );
BUF_X2 newInst_1157 ( .a(newNet_1156), .o(newNet_1157) );
NAND2_Z01 g60510 ( .a(n_360), .b(GPR_1__6_), .o(n_636) );
BUF_X2 newInst_1425 ( .a(newNet_1424), .o(newNet_1425) );
NOR3_Z1 g60660 ( .a(n_116), .b(n_253), .c(pZ_0_), .o(n_485) );
NOR2_Z1 g60585 ( .a(n_471), .b(n_71), .o(n_527) );
NAND2_Z01 g34744 ( .a(n_3591), .b(U_13_), .o(n_3821) );
NAND2_Z01 g58874 ( .a(n_2153), .b(GPR_8__0_), .o(n_2233) );
AND2_X1 g58451 ( .a(n_2604), .b(n_587), .o(n_2643) );
NAND2_Z01 g34901 ( .a(n_3590), .b(pY_9_), .o(n_3662) );
NAND2_Z01 g60572 ( .a(n_341), .b(pZ_4_), .o(n_539) );
NAND2_Z01 g60431 ( .a(n_457), .b(GPR_18__4_), .o(n_715) );
AND2_X1 g60059 ( .a(n_844), .b(n_52), .o(n_1075) );
NAND2_Z03 g34173 ( .a(n_4314), .b(n_3951), .o(io_do_7) );
BUF_X2 newInst_319 ( .a(newNet_318), .o(newNet_319) );
BUF_X2 newInst_461 ( .a(newNet_460), .o(newNet_461) );
NAND2_Z01 g59430 ( .a(n_1647), .b(n_763), .o(n_1689) );
NOR2_Z1 g59433 ( .a(n_1646), .b(n_1107), .o(n_1686) );
NAND2_Z01 g58472 ( .a(n_2363), .b(n_2584), .o(n_2624) );
NAND2_Z01 g59085 ( .a(n_1857), .b(SP_15_), .o(n_2022) );
NAND2_Z01 g58758 ( .a(n_2203), .b(GPR_4__2_), .o(n_2342) );
NOR3_Z1 g35372 ( .a(n_3249), .b(n_3231), .c(n_3233), .o(n_3318) );
NAND2_Z01 g59755 ( .a(n_1312), .b(io_do_4), .o(n_1369) );
BUF_X2 newInst_127 ( .a(newNet_6), .o(newNet_127) );
XOR2_X1 g59450 ( .a(n_1622), .b(SP_13_), .o(n_1672) );
NAND2_Z01 g58749 ( .a(n_2204), .b(GPR_3__1_), .o(n_2351) );
BUF_X2 newInst_41 ( .a(newNet_40), .o(newNet_41) );
NAND2_Z01 g60184 ( .a(n_686), .b(n_685), .o(n_956) );
NAND2_Z01 g61011 ( .a(n_36), .b(n_43), .o(n_170) );
NOR2_Z1 g60642 ( .a(n_460), .b(n_182), .o(n_575) );
NAND2_Z01 g34307 ( .a(n_4161), .b(n_4566), .o(n_4226) );
NAND2_Z01 g34693 ( .a(n_3635), .b(GPR_14__6_), .o(n_3872) );
NAND2_Z01 g35301 ( .a(n_3289), .b(pY_2_), .o(n_3374) );
NAND3_Z1 g59249 ( .a(n_1745), .b(n_1365), .c(n_1279), .o(n_1863) );
NAND4_Z1 g57910 ( .a(n_1964), .b(n_2507), .c(n_2990), .d(n_2027), .o(n_3029) );
NOR4_Z1 g34232 ( .a(n_4222), .b(n_4223), .c(n_4246), .d(n_4121), .o(n_4299) );
BUF_X2 newInst_1520 ( .a(newNet_1519), .o(newNet_1520) );
BUF_X2 newInst_1322 ( .a(newNet_1321), .o(newNet_1322) );
BUF_X2 newInst_1300 ( .a(newNet_479), .o(newNet_1300) );
XOR2_X1 final_adder_mux_R16_278_6_g420 ( .a(n_4441), .b(n_4425), .o(final_adder_mux_R16_278_6_n_29) );
NOR4_Z1 g59030 ( .a(n_1780), .b(n_1461), .c(n_1251), .d(n_1816), .o(n_2074) );
fflopd GPR_reg_17__5_ ( .CK(newNet_1384), .D(n_3014), .Q(GPR_17__5_) );
NAND2_Z02 g34381 ( .a(n_3209), .b(n_4070), .o(n_4159) );
NOR2_Z1 g34343 ( .a(n_4159), .b(n_3454), .o(n_4191) );
NAND2_Z01 g60250 ( .a(n_596), .b(GPR_3__7_), .o(n_895) );
NAND2_Z01 g60738 ( .a(SP_11_), .b(n_180), .o(n_401) );
NAND2_Z01 g34640 ( .a(n_3769), .b(pZ_10_), .o(n_3920) );
NAND2_Z01 g60712 ( .a(GPR_4__4_), .b(n_183), .o(n_426) );
BUF_X2 newInst_982 ( .a(newNet_981), .o(newNet_982) );
NOR2_Z1 g60830 ( .a(n_216), .b(n_4668), .o(n_301) );
INV_X1 g60778 ( .a(n_337), .o(n_336) );
BUF_X2 newInst_31 ( .a(newNet_30), .o(newNet_31) );
NAND2_Z01 g35035 ( .a(n_4517), .b(n_3255), .o(n_3545) );
AND2_X1 g59470 ( .a(n_1628), .b(n_101), .o(n_1654) );
NAND2_Z01 g58152 ( .a(n_2813), .b(n_2242), .o(n_2861) );
NAND2_Z02 g60359 ( .a(n_66), .b(n_573), .o(n_850) );
INV_X1 g35488 ( .a(pZ_10_), .o(n_3237) );
NAND2_Z01 g58763 ( .a(n_2203), .b(GPR_4__7_), .o(n_2337) );
fflopd GPR_reg_7__1_ ( .CK(newNet_779), .D(n_2740), .Q(GPR_7__1_) );
BUF_X2 newInst_917 ( .a(newNet_400), .o(newNet_917) );
NAND4_Z1 g60135 ( .a(n_713), .b(n_716), .c(n_714), .d(n_717), .o(n_997) );
BUF_X2 newInst_489 ( .a(newNet_488), .o(newNet_489) );
NAND4_Z1 g59989 ( .a(n_871), .b(n_833), .c(n_937), .d(n_886), .o(n_1140) );
NOR2_Z1 g59483 ( .a(n_1619), .b(n_972), .o(n_1642) );
NAND2_Z01 g34866 ( .a(n_3585), .b(GPR_13__0_), .o(n_3697) );
NAND2_Z01 g60491 ( .a(n_372), .b(U_10_), .o(n_655) );
NAND2_Z01 g57693 ( .a(n_3158), .b(n_1771), .o(n_3173) );
BUF_X2 newInst_1383 ( .a(newNet_1382), .o(newNet_1383) );
NAND2_Z01 g58995 ( .a(n_2023), .b(n_265), .o(n_2111) );
NAND2_Z01 g57929 ( .a(n_2978), .b(n_2237), .o(n_3016) );
fflopd GPR_reg_4__0_ ( .CK(newNet_929), .D(n_2623), .Q(GPR_4__0_) );
NOR2_Z1 g60933 ( .a(n_104), .b(rst), .o(n_255) );
BUF_X2 newInst_1379 ( .a(newNet_1370), .o(newNet_1379) );
NOR2_Z1 g60782 ( .a(io_do_0), .b(n_261), .o(n_381) );
NOR2_Z1 g59790 ( .a(n_1248), .b(n_1023), .o(n_1334) );
NAND2_Z01 g60214 ( .a(n_577), .b(pZ_10_), .o(n_931) );
AND4_X1 g58938 ( .a(n_1820), .b(n_1862), .c(n_2093), .d(n_1687), .o(n_2169) );
NAND2_Z01 g58331 ( .a(n_2662), .b(n_2308), .o(n_2734) );
BUF_X2 newInst_66 ( .a(newNet_65), .o(newNet_66) );
BUF_X2 newInst_614 ( .a(newNet_613), .o(newNet_614) );
BUF_X2 newInst_1861 ( .a(newNet_1860), .o(newNet_1861) );
NOR2_Z1 g59793 ( .a(n_1265), .b(n_1166), .o(n_1331) );
INV_Z1 g16805 ( .a(GPR_8__3_), .o(n_4404) );
BUF_X2 newInst_1752 ( .a(newNet_54), .o(newNet_1752) );
NAND2_Z01 g59059 ( .a(n_1902), .b(n_4595), .o(n_2048) );
NAND2_Z01 g58808 ( .a(n_2197), .b(U_6_), .o(n_2292) );
BUF_X2 newInst_776 ( .a(newNet_775), .o(newNet_776) );
NAND2_Z01 g60547 ( .a(n_370), .b(GPR_20__2_), .o(n_559) );
NAND4_Z1 g57725 ( .a(n_2953), .b(n_3009), .c(n_3115), .d(n_24), .o(n_3144) );
NAND2_Z01 g34628 ( .a(n_3769), .b(pZ_11_), .o(n_3932) );
BUF_X2 newInst_78 ( .a(newNet_46), .o(newNet_78) );
NAND2_Z01 g58172 ( .a(n_2794), .b(n_2307), .o(n_2838) );
NAND2_Z01 g59224 ( .a(n_1824), .b(n_1804), .o(n_1899) );
XOR2_X1 final_adder_mux_R16_278_6_g385 ( .a(final_adder_mux_R16_278_6_n_62), .b(final_adder_mux_R16_278_6_n_42), .o(R16_7_) );
NAND2_Z01 g34147 ( .a(n_4325), .b(n_4614), .o(n_4361) );
BUF_X2 newInst_9 ( .a(newNet_8), .o(newNet_9) );
BUF_X2 newInst_1819 ( .a(newNet_1818), .o(newNet_1819) );
INV_X1 g61042 ( .a(pZ_12_), .o(n_110) );
NOR4_Z1 g60161 ( .a(n_484), .b(n_312), .c(n_4480), .d(n_4642), .o(n_975) );
NAND2_Z01 g34520 ( .a(n_3870), .b(n_3948), .o(n_4023) );
NAND2_Z01 g58588 ( .a(n_2482), .b(n_1705), .o(n_2510) );
fflopd GPR_reg_22__1_ ( .CK(newNet_1105), .D(n_2761), .Q(GPR_22__1_) );
NAND2_Z01 g34697 ( .a(n_3567), .b(GPR_6__6_), .o(n_3868) );
NAND2_Z01 g58898 ( .a(n_2157), .b(GPR_13__4_), .o(n_2184) );
NOR2_Z1 g34399 ( .a(n_4086), .b(n_3469), .o(n_4139) );
NAND2_Z01 g60731 ( .a(n_200), .b(GPR_9__1_), .o(n_408) );
NOR2_Z2 g35419 ( .a(n_3244), .b(pmem_d_5), .o(n_3299) );
XNOR2_X1 g58833 ( .a(n_2136), .b(PC_10_), .o(n_2274) );
BUF_X2 newInst_417 ( .a(newNet_416), .o(newNet_417) );
NOR2_Z1 g34339 ( .a(n_4612), .b(n_3421), .o(n_4195) );
XOR2_X1 g59811 ( .a(n_1217), .b(pX_7_), .o(n_1318) );
INV_X1 g35023 ( .a(n_3551), .o(n_3550) );
BUF_X2 newInst_1061 ( .a(newNet_1060), .o(newNet_1061) );
NOR2_Z1 g60931 ( .a(n_4560), .b(n_104), .o(n_215) );
NAND2_Z01 g60739 ( .a(n_203), .b(SP_3_), .o(n_400) );
NAND2_Z01 g60699 ( .a(GPR_4__1_), .b(n_183), .o(n_439) );
NAND2_Z01 g57686 ( .a(n_3157), .b(n_2218), .o(n_3180) );
BUF_X2 newInst_707 ( .a(newNet_706), .o(newNet_707) );
BUF_X2 newInst_445 ( .a(newNet_444), .o(newNet_445) );
NOR2_Z1 g60590 ( .a(n_369), .b(n_4536), .o(n_608) );
AND2_X1 g34332 ( .a(n_4178), .b(n_4101), .o(n_4202) );
BUF_X2 newInst_456 ( .a(newNet_455), .o(newNet_456) );
XNOR2_X1 g34932 ( .a(n_3539), .b(pX_12_), .o(n_4562) );
BUF_X2 newInst_1131 ( .a(newNet_1130), .o(newNet_1131) );
XOR2_X1 g60007 ( .a(n_859), .b(n_55), .o(n_1157) );
NAND2_Z01 g59696 ( .a(io_do_3), .b(n_1353), .o(n_1434) );
NAND4_Z1 g59591 ( .a(n_1383), .b(n_842), .c(n_66), .d(n_860), .o(n_1537) );
BUF_X2 newInst_440 ( .a(newNet_439), .o(newNet_440) );
XOR2_X1 g60864 ( .a(n_4443), .b(n_4427), .o(n_284) );
AND2_X1 g60062 ( .a(n_844), .b(n_47), .o(n_1072) );
NAND3_Z1 g34553 ( .a(n_3761), .b(n_3770), .c(n_3771), .o(n_4006) );
BUF_X2 newInst_885 ( .a(newNet_884), .o(newNet_885) );
NAND2_Z01 g58301 ( .a(n_2695), .b(n_2421), .o(n_2769) );
NAND2_Z01 g34601 ( .a(n_3814), .b(n_3303), .o(n_3960) );
fflopd U_reg_2_ ( .CK(newNet_384), .D(n_2867), .Q(U_2_) );
NAND2_Z01 g59333 ( .a(n_1223), .b(n_15), .o(n_1781) );
BUF_X2 newInst_1261 ( .a(newNet_188), .o(newNet_1261) );
BUF_X2 newInst_914 ( .a(newNet_913), .o(newNet_914) );
XOR2_X1 g35256 ( .a(n_3285), .b(pZ_2_), .o(n_4608) );
AND2_X1 g57904 ( .a(n_3009), .b(n_2201), .o(n_3034) );
NOR2_Z1 g60361 ( .a(n_592), .b(SP_4_), .o(n_847) );
NAND2_Z01 g59150 ( .a(n_1896), .b(n_752), .o(n_1949) );
NAND2_Z01 g34363 ( .a(n_3209), .b(n_4039), .o(n_4177) );
NAND2_Z01 g58353 ( .a(n_2647), .b(n_2290), .o(n_2718) );
BUF_X2 newInst_546 ( .a(newNet_545), .o(newNet_546) );
NAND4_Z1 g58141 ( .a(n_2126), .b(n_2542), .c(n_2831), .d(n_2033), .o(n_2872) );
NAND2_Z01 g60430 ( .a(n_457), .b(GPR_16__2_), .o(n_716) );
AND2_X1 g58105 ( .a(n_2850), .b(n_2139), .o(n_2907) );
NOR2_Z1 g34313 ( .a(n_4612), .b(n_3520), .o(n_4220) );
BUF_X2 newInst_1826 ( .a(newNet_1825), .o(newNet_1826) );
BUF_X2 newInst_1076 ( .a(newNet_1075), .o(newNet_1076) );
NAND2_Z01 g59615 ( .a(n_1414), .b(io_di_2), .o(n_1512) );
BUF_X2 newInst_930 ( .a(newNet_363), .o(newNet_930) );
BUF_X2 newInst_388 ( .a(newNet_387), .o(newNet_388) );
NAND2_Z01 g59571 ( .a(n_1469), .b(n_222), .o(n_1557) );
AND2_X1 g34445 ( .a(n_4073), .b(n_3218), .o(n_4094) );
fflopd GPR_reg_8__6_ ( .CK(newNet_698), .D(n_3066), .Q(GPR_8__6_) );
BUF_X2 newInst_593 ( .a(newNet_592), .o(newNet_593) );
NAND2_Z01 g59608 ( .a(n_1413), .b(io_sp_0_), .o(n_1518) );
NOR4_Z1 g34195 ( .a(n_4185), .b(n_4259), .c(n_4301), .d(n_4104), .o(n_4328) );
NAND2_Z01 g34831 ( .a(n_3571), .b(GPR_20__1_), .o(n_3732) );
NAND2_Z01 g58812 ( .a(n_2199), .b(GPR_0__6_), .o(n_2288) );
BUF_X2 newInst_1199 ( .a(newNet_114), .o(newNet_1199) );
BUF_X2 newInst_760 ( .a(newNet_759), .o(newNet_760) );
NAND2_Z01 g34536 ( .a(n_3907), .b(n_3933), .o(pmem_a_0) );
NOR2_Z1 g59286 ( .a(n_1760), .b(n_1548), .o(n_1834) );
NAND2_Z01 g34758 ( .a(n_3636), .b(GPR_10__4_), .o(n_3807) );
BUF_X2 newInst_1676 ( .a(newNet_1675), .o(newNet_1676) );
BUF_X2 newInst_1422 ( .a(newNet_1421), .o(newNet_1422) );
BUF_X2 newInst_1619 ( .a(newNet_1618), .o(newNet_1619) );
BUF_X2 newInst_562 ( .a(newNet_561), .o(newNet_562) );
BUF_X2 newInst_333 ( .a(newNet_332), .o(newNet_333) );
BUF_X2 newInst_1562 ( .a(newNet_1561), .o(newNet_1562) );
NOR2_Z1 g34993 ( .a(n_3531), .b(state_3_), .o(n_3560) );
NAND2_Z01 g35134 ( .a(Rd_3_), .b(n_3225), .o(n_3484) );
NAND2_Z01 g59140 ( .a(n_1894), .b(n_46), .o(n_1959) );
NAND2_Z01 g58710 ( .a(n_2209), .b(GPR_20__7_), .o(n_2397) );
XOR2_X1 g35199 ( .a(n_3415), .b(PC_3_), .o(n_4549) );
NOR2_Z1 g60742 ( .a(n_278), .b(n_107), .o(n_467) );
NAND2_Z01 g58843 ( .a(n_2139), .b(GPR_11__2_), .o(n_2264) );
NAND2_Z01 g57724 ( .a(n_3131), .b(n_915), .o(n_3157) );
NAND4_Z1 g59305 ( .a(n_1604), .b(n_1434), .c(n_1715), .d(n_1007), .o(n_1809) );
NAND2_Z01 g58786 ( .a(n_2200), .b(GPR_7__5_), .o(n_2314) );
NAND2_Z01 g35044 ( .a(n_4517), .b(n_4518), .o(n_3537) );
NAND2_Z01 g60445 ( .a(n_457), .b(GPR_18__1_), .o(n_701) );
NAND2_Z01 g34191 ( .a(n_4325), .b(n_4467), .o(n_4332) );
INV_X1 g58992 ( .a(n_2116), .o(n_2115) );
XOR2_X1 g59207 ( .a(n_1851), .b(n_320), .o(n_1904) );
NAND2_Z01 g59973 ( .a(n_973), .b(n_849), .o(n_1151) );
AND2_X1 g59277 ( .a(n_1739), .b(n_1269), .o(n_1837) );
NOR2_Z1 g35125 ( .a(n_4656), .b(n_3297), .o(n_4655) );
NOR2_Z1 g34808 ( .a(n_3598), .b(n_4402), .o(n_3755) );
INV_X1 drc_bufs35519 ( .a(n_3208), .o(n_4611) );
BUF_X2 newInst_1791 ( .a(newNet_953), .o(newNet_1791) );
BUF_X2 newInst_1737 ( .a(newNet_1736), .o(newNet_1737) );
NAND2_Z01 g35287 ( .a(U_2_), .b(n_3275), .o(n_3388) );
NAND2_Z01 g60926 ( .a(io_do_0), .b(io_do_1), .o(n_259) );
NAND2_Z01 g60321 ( .a(n_600), .b(pX_3_), .o(n_806) );
NAND3_Z1 g59767 ( .a(n_494), .b(n_1175), .c(n_242), .o(n_1385) );
NAND2_Z01 g59129 ( .a(n_1872), .b(n_1557), .o(n_1967) );
NOR2_Z1 g59490 ( .a(n_1565), .b(n_1602), .o(n_1648) );
fflopd GPR_reg_15__5_ ( .CK(newNet_1491), .D(n_3016), .Q(GPR_15__5_) );
BUF_X2 newInst_673 ( .a(newNet_672), .o(newNet_673) );
NAND4_Z1 g59985 ( .a(n_731), .b(n_505), .c(n_755), .d(n_240), .o(n_1143) );
INV_X1 g34978 ( .a(n_3578), .o(n_3577) );
BUF_X2 newInst_1193 ( .a(newNet_1192), .o(newNet_1193) );
BUF_X2 newInst_1126 ( .a(newNet_546), .o(newNet_1126) );
BUF_X2 newInst_316 ( .a(newNet_114), .o(newNet_316) );
BUF_X2 newInst_88 ( .a(newNet_0), .o(newNet_88) );
NAND2_Z01 g58319 ( .a(n_2676), .b(n_2343), .o(n_2746) );
INV_X1 g59576 ( .a(n_1552), .o(n_1553) );
NAND2_Z01 g59360 ( .a(n_1038), .b(n_1729), .o(n_1753) );
NAND2_Z01 g58952 ( .a(n_2114), .b(n_1835), .o(n_2148) );
BUF_X2 newInst_17 ( .a(newNet_1), .o(newNet_17) );
BUF_X2 newInst_21 ( .a(newNet_20), .o(newNet_21) );
AND2_X1 g58507 ( .a(n_2567), .b(n_2209), .o(n_2590) );
BUF_X2 newInst_1543 ( .a(newNet_1542), .o(newNet_1543) );
BUF_X2 newInst_1004 ( .a(newNet_1003), .o(newNet_1004) );
NAND2_Z01 g58305 ( .a(n_2692), .b(n_2403), .o(n_2765) );
NAND2_Z01 g35399 ( .a(pmem_d_5), .b(pmem_d_4), .o(n_3309) );
NAND2_Z01 g57943 ( .a(n_2964), .b(n_2323), .o(n_2999) );
NAND2_Z01 g59601 ( .a(n_1451), .b(SP_13_), .o(n_1525) );
BUF_X2 newInst_242 ( .a(newNet_241), .o(newNet_242) );
NOR2_Z1 g60577 ( .a(n_301), .b(n_32), .o(n_534) );
NAND2_Z01 g58878 ( .a(n_2153), .b(GPR_8__4_), .o(n_2229) );
NAND4_Z1 g59253 ( .a(n_1638), .b(n_1431), .c(n_1779), .d(n_1008), .o(n_1859) );
BUF_X2 newInst_214 ( .a(newNet_211), .o(newNet_214) );
BUF_X2 newInst_1248 ( .a(newNet_1247), .o(newNet_1248) );
NAND2_Z01 g61025 ( .a(n_44), .b(n_62), .o(n_160) );
BUF_X2 newInst_385 ( .a(newNet_65), .o(newNet_385) );
NOR3_Z2 g59424 ( .a(n_1040), .b(n_1489), .c(n_1602), .o(n_1700) );
BUF_X2 newInst_1625 ( .a(newNet_1624), .o(newNet_1625) );
BUF_X2 newInst_1393 ( .a(newNet_1392), .o(newNet_1393) );
NAND2_Z01 g60202 ( .a(n_577), .b(pZ_11_), .o(n_943) );
NOR2_Z1 g34861 ( .a(n_3596), .b(n_4409), .o(n_3702) );
NAND2_Z01 g60490 ( .a(n_368), .b(GPR_15__1_), .o(n_656) );
BUF_X2 newInst_165 ( .a(newNet_164), .o(newNet_165) );
NAND2_Z01 g58446 ( .a(n_2621), .b(n_2196), .o(n_2647) );
NAND2_Z03 g34169 ( .a(n_4316), .b(n_3955), .o(io_do_1) );
NAND2_Z01 g34962 ( .a(n_3536), .b(pY_11_), .o(n_3600) );
INV_X1 g35472 ( .a(state_2_), .o(n_3252) );
INV_X1 g59210 ( .a(n_1896), .o(n_1895) );
INV_X1 g59909 ( .a(n_1214), .o(n_1215) );
NAND2_Z01 g58742 ( .a(n_2213), .b(GPR_17__3_), .o(n_2365) );
BUF_X2 newInst_1599 ( .a(newNet_1099), .o(newNet_1599) );
BUF_X2 newInst_1538 ( .a(newNet_1364), .o(newNet_1538) );
INV_Z1 g16797 ( .a(n_4466), .o(n_4415) );
BUF_X2 newInst_787 ( .a(newNet_786), .o(newNet_787) );
NOR2_Z1 g60261 ( .a(n_581), .b(n_75), .o(n_885) );
NAND2_Z01 g58526 ( .a(n_2563), .b(n_1817), .o(n_2571) );
fflopd pX_reg_12_ ( .CK(newNet_264), .D(n_3024), .Q(pX_12_) );
BUF_X2 newInst_210 ( .a(newNet_209), .o(newNet_210) );
INV_X1 drc_bufs35574 ( .a(n_3592), .o(n_3196) );
BUF_X2 newInst_821 ( .a(newNet_820), .o(newNet_821) );
NOR2_Z1 g59841 ( .a(n_1032), .b(n_1170), .o(n_1285) );
NAND2_Z01 g59238 ( .a(n_1850), .b(n_1852), .o(n_1879) );
NOR3_Z1 g35098 ( .a(n_4484), .b(n_3479), .c(n_4638), .o(n_3496) );
NAND2_Z01 g34359 ( .a(n_4152), .b(SP_5_), .o(n_4172) );
INV_X1 g35038 ( .a(n_4567), .o(n_3534) );
NAND2_Z01 g58707 ( .a(n_2209), .b(GPR_20__4_), .o(n_2400) );
AND2_X1 g60599 ( .a(n_381), .b(pmem_d_0), .o(n_519) );
BUF_X2 newInst_255 ( .a(newNet_254), .o(newNet_255) );
NAND2_Z01 g60410 ( .a(n_353), .b(GPR_8__5_), .o(n_736) );
NAND2_Z01 g34687 ( .a(n_3584), .b(GPR_21__7_), .o(n_3878) );
NAND2_Z01 g34714 ( .a(n_3584), .b(GPR_21__6_), .o(n_3851) );
NAND2_Z01 g34794 ( .a(n_3586), .b(GPR_9__3_), .o(n_3771) );
INV_X1 g35498 ( .a(pX_6_), .o(n_3229) );
NAND2_Z01 g35267 ( .a(n_3299), .b(pX_14_), .o(n_3406) );
NAND4_Z1 g58018 ( .a(n_1949), .b(n_2454), .c(n_2917), .d(n_2047), .o(n_2954) );
BUF_X2 newInst_1217 ( .a(newNet_1216), .o(newNet_1217) );
NAND2_Z01 g57803 ( .a(n_3079), .b(n_2194), .o(n_3104) );
BUF_X2 newInst_1401 ( .a(newNet_113), .o(newNet_1401) );
BUF_X2 newInst_360 ( .a(newNet_359), .o(newNet_360) );
INV_X1 g35325 ( .a(n_3344), .o(n_4573) );
BUF_X2 newInst_33 ( .a(newNet_32), .o(newNet_33) );
NAND2_Z01 g59336 ( .a(io_do_0), .b(n_1695), .o(n_1804) );
NOR2_Z1 g34327 ( .a(n_4159), .b(n_3903), .o(n_4207) );
NOR3_Z1 g34496 ( .a(n_4005), .b(n_3972), .c(n_4016), .o(n_4048) );
NAND2_Z01 g59053 ( .a(n_1875), .b(n_4568), .o(n_2054) );
BUF_X2 newInst_1187 ( .a(newNet_1186), .o(newNet_1187) );
NAND2_Z01 g34080 ( .a(n_4164), .b(GPR_Rd_r_7_), .o(n_4393) );
NAND2_Z01 g60694 ( .a(n_198), .b(GPR_17__1_), .o(n_444) );
NOR2_Z1 g34270 ( .a(n_4613), .b(n_3212), .o(n_4263) );
BUF_X2 newInst_747 ( .a(newNet_746), .o(newNet_747) );
NAND2_Z01 g34966 ( .a(n_3536), .b(n_3491), .o(n_3632) );
INV_X1 g61110 ( .a(pmem_d_15), .o(n_42) );
NAND2_Z01 g59701 ( .a(io_do_2), .b(n_1353), .o(n_1429) );
AND4_X1 g34067 ( .a(n_4236), .b(n_4245), .c(n_4396), .d(n_4135), .o(dmem_a_10) );
NAND2_Z01 g60248 ( .a(n_590), .b(GPR_6__7_), .o(n_897) );
AND2_X1 g59348 ( .a(io_do_3), .b(n_30), .o(n_1772) );
NAND2_Z01 g59267 ( .a(n_1782), .b(n_206), .o(n_1854) );
BUF_X2 newInst_1813 ( .a(newNet_1317), .o(newNet_1813) );
BUF_X2 newInst_780 ( .a(newNet_484), .o(newNet_780) );
BUF_X2 newInst_1517 ( .a(newNet_1516), .o(newNet_1517) );
NOR3_Z1 g60844 ( .a(n_71), .b(n_4651), .c(n_44), .o(n_294) );
BUF_X2 newInst_532 ( .a(newNet_531), .o(newNet_532) );
BUF_X2 newInst_1844 ( .a(newNet_1843), .o(newNet_1844) );
NAND2_Z01 g60306 ( .a(n_597), .b(pX_11_), .o(n_818) );
BUF_X2 newInst_1276 ( .a(newNet_1275), .o(newNet_1276) );
NAND4_Z1 g58988 ( .a(n_1936), .b(n_1261), .c(n_1843), .d(n_1262), .o(n_2119) );
BUF_X2 newInst_125 ( .a(newNet_124), .o(newNet_125) );
NAND4_Z1 g59546 ( .a(n_796), .b(n_1297), .c(n_1501), .d(n_1075), .o(n_1582) );
NAND2_Z01 g34526 ( .a(n_3822), .b(n_3943), .o(n_4018) );
NAND2_Z01 g35453 ( .a(n_3245), .b(n_3254), .o(n_3268) );
INV_Z1 g16802 ( .a(n_4468), .o(n_4416) );
BUF_X2 newInst_1483 ( .a(newNet_1482), .o(newNet_1483) );
NAND2_Z01 g34852 ( .a(n_3571), .b(GPR_20__0_), .o(n_3711) );
NAND2_Z01 g60421 ( .a(n_342), .b(GPR_19__4_), .o(n_725) );
NOR2_Z1 g58925 ( .a(n_2118), .b(n_579), .o(n_2178) );
XOR2_X1 final_adder_mux_R16_278_6_g405 ( .a(n_4442), .b(n_4426), .o(final_adder_mux_R16_278_6_n_44) );
NAND2_Z01 g60767 ( .a(n_178), .b(n_90), .o(n_382) );
BUF_X2 newInst_353 ( .a(newNet_352), .o(newNet_353) );
INV_X1 g61044 ( .a(C), .o(n_108) );
INV_X2 newInst_328 ( .a(newNet_327), .o(newNet_328) );
BUF_X2 newInst_1561 ( .a(newNet_1560), .o(newNet_1561) );
NOR2_Z1 g34417 ( .a(n_4096), .b(n_3982), .o(n_4120) );
BUF_X2 newInst_288 ( .a(newNet_287), .o(newNet_288) );
AND2_X1 g59856 ( .a(n_1219), .b(n_165), .o(n_1273) );
XOR2_X1 g60857 ( .a(n_4561), .b(n_119), .o(n_287) );
XOR2_X1 g60389 ( .a(n_290), .b(n_136), .o(n_757) );
NAND2_Z01 g59131 ( .a(n_1900), .b(n_1892), .o(n_1984) );
BUF_X2 newInst_1087 ( .a(newNet_1086), .o(newNet_1087) );
fflopd GPR_reg_1__6_ ( .CK(newNet_1222), .D(n_3077), .Q(GPR_1__6_) );
BUF_X2 newInst_979 ( .a(newNet_978), .o(newNet_979) );
NAND2_Z01 g60419 ( .a(n_342), .b(GPR_17__2_), .o(n_727) );
AND2_X1 g58500 ( .a(n_2567), .b(n_2155), .o(n_2597) );
NAND2_Z01 g59612 ( .a(n_1415), .b(Z), .o(n_1515) );
NOR4_Z1 g58654 ( .a(n_1438), .b(n_2127), .c(n_2064), .d(n_1412), .o(n_2448) );
NAND2_Z01 g60701 ( .a(pY_9_), .b(n_249), .o(n_437) );
BUF_X2 newInst_81 ( .a(newNet_80), .o(newNet_81) );
NAND2_Z01 g34635 ( .a(n_3769), .b(pZ_7_), .o(n_3925) );
fflopd GPR_reg_2__1_ ( .CK(newNet_1018), .D(n_2750), .Q(GPR_2__1_) );
NAND2_Z01 g35295 ( .a(n_3299), .b(pX_2_), .o(n_3380) );
AND2_X1 g58337 ( .a(n_2688), .b(n_587), .o(n_2732) );
NAND4_Z1 g57813 ( .a(n_1948), .b(n_2453), .c(n_3061), .d(n_2028), .o(n_3094) );
NAND4_Z1 g57735 ( .a(n_2073), .b(n_2539), .c(n_3107), .d(n_1973), .o(n_3137) );
NAND2_Z01 g60983 ( .a(n_122), .b(n_48), .o(n_146) );
BUF_X2 newInst_1100 ( .a(newNet_1099), .o(newNet_1100) );
BUF_X2 newInst_567 ( .a(newNet_566), .o(newNet_567) );
NAND2_Z01 g58538 ( .a(n_2541), .b(n_1988), .o(n_2563) );
fflopd GPR_reg_15__4_ ( .CK(newNet_1502), .D(n_2944), .Q(GPR_15__4_) );
BUF_X2 newInst_670 ( .a(newNet_533), .o(newNet_670) );
BUF_X2 newInst_405 ( .a(newNet_301), .o(newNet_405) );
NAND4_Z1 g60132 ( .a(n_681), .b(n_555), .c(n_653), .d(n_626), .o(n_1000) );
INV_X2 newInst_1362 ( .a(newNet_1361), .o(newNet_1362) );
NAND2_Z01 g34619 ( .a(n_3893), .b(n_3461), .o(n_3941) );
NAND2_Z01 g60265 ( .a(n_578), .b(GPR_19__6_), .o(n_881) );
NAND2_Z01 g60956 ( .a(n_35), .b(pmem_d_0), .o(n_205) );
NAND2_Z01 g59329 ( .a(n_1699), .b(dmem_di_1), .o(n_1784) );
NAND4_Z1 g60155 ( .a(n_540), .b(n_632), .c(n_633), .d(n_631), .o(n_980) );
NOR2_Z1 g34923 ( .a(n_3569), .b(n_3348), .o(n_3642) );
NAND2_Z01 final_adder_mux_R16_278_6_g430 ( .a(n_4444), .b(n_4428), .o(final_adder_mux_R16_278_6_n_19) );
AND2_X1 g57892 ( .a(n_3009), .b(n_2213), .o(n_3046) );
NOR2_Z1 g58967 ( .a(n_2089), .b(n_965), .o(n_2152) );
NAND2_Z01 g57701 ( .a(n_3143), .b(n_2266), .o(n_3168) );
NOR3_Z1 g34925 ( .a(n_3530), .b(n_3525), .c(pmem_d_1), .o(n_3640) );
fflopd N_reg ( .CK(newNet_663), .D(n_3185), .Q(N) );
NAND2_Z01 g60221 ( .a(n_582), .b(GPR_11__2_), .o(n_924) );
NAND2_Z01 g34508 ( .a(n_4010), .b(n_3932), .o(pmem_a_10) );
BUF_X2 newInst_1610 ( .a(newNet_2), .o(newNet_1610) );
NAND3_Z1 g59585 ( .a(n_1374), .b(n_1488), .c(n_409), .o(n_1543) );
NAND2_Z01 g34105 ( .a(n_4336), .b(n_4355), .o(n_4451) );
AND2_X1 g57741 ( .a(n_3115), .b(n_2210), .o(n_3130) );
NAND2_Z01 g58624 ( .a(n_2354), .b(pX_0_), .o(n_2473) );
XOR2_X1 g35106 ( .a(n_3470), .b(PC_5_), .o(n_4545) );
AND2_X1 g58647 ( .a(n_2354), .b(n_1963), .o(n_2460) );
BUF_X2 newInst_1366 ( .a(newNet_1365), .o(newNet_1366) );
AND3_X1 g59492 ( .a(n_1312), .b(n_1539), .c(n_1038), .o(n_1635) );
NAND2_Z01 g34683 ( .a(n_3627), .b(GPR_15__7_), .o(n_3882) );
BUF_X2 newInst_1374 ( .a(newNet_1373), .o(newNet_1374) );
BUF_X2 newInst_1288 ( .a(newNet_1287), .o(newNet_1288) );
NAND2_Z01 g60714 ( .a(n_200), .b(GPR_8__1_), .o(n_424) );
AND2_X1 g58125 ( .a(n_2850), .b(n_2200), .o(n_2887) );
NAND2_Z01 g58053 ( .a(n_2891), .b(n_2348), .o(n_2929) );
NAND3_Z1 g35185 ( .a(n_3376), .b(n_3437), .c(n_3393), .o(n_4623) );
fflopd io_sp_reg_2_ ( .CK(newNet_329), .D(n_550), .Q(io_sp_2_) );
BUF_X2 newInst_818 ( .a(newNet_817), .o(newNet_818) );
AND2_X1 g58001 ( .a(n_2940), .b(n_2207), .o(n_2970) );
NAND4_Z1 g57756 ( .a(n_2080), .b(n_2538), .c(n_3105), .d(n_1968), .o(n_3116) );
NAND2_Z01 g59512 ( .a(n_1541), .b(SP_9_), .o(n_1610) );
BUF_X2 newInst_721 ( .a(newNet_720), .o(newNet_721) );
AND2_X1 g58403 ( .a(n_2657), .b(n_2140), .o(n_2665) );
NAND2_Z01 g34504 ( .a(n_4002), .b(SP_0_), .o(n_4040) );
BUF_X2 newInst_1707 ( .a(newNet_1706), .o(newNet_1707) );
AND2_X1 g34468 ( .a(n_4057), .b(n_3222), .o(n_4074) );
NOR2_Z1 g60652 ( .a(n_364), .b(n_152), .o(n_489) );
NAND2_Z01 g35223 ( .a(n_4658), .b(pmem_d_13), .o(n_3446) );
INV_X1 g61056 ( .a(pY_2_), .o(n_96) );
AND3_X1 g59189 ( .a(n_465), .b(n_1873), .c(pX_3_), .o(n_1918) );
NAND2_Z01 g58979 ( .a(n_2084), .b(n_1215), .o(n_2128) );
BUF_X2 newInst_1647 ( .a(newNet_1646), .o(newNet_1647) );
NOR3_Z1 g59184 ( .a(n_1666), .b(n_1873), .c(n_99), .o(n_1923) );
BUF_X2 newInst_1467 ( .a(newNet_1466), .o(newNet_1467) );
fflopd GPR_reg_2__0_ ( .CK(newNet_1019), .D(n_2625), .Q(GPR_2__0_) );
NAND2_Z01 g60311 ( .a(n_600), .b(pX_2_), .o(n_815) );
NAND2_Z01 g34130 ( .a(n_4164), .b(GPR_Rd_r_6_), .o(n_4378) );
NAND2_Z01 g60889 ( .a(n_58), .b(n_4479), .o(n_238) );
NAND2_Z01 g59088 ( .a(n_1875), .b(n_4564), .o(n_2019) );
INV_X1 g34372 ( .a(n_16064_BAR), .o(n_4160) );
fflopd pZ_reg_15_ ( .CK(newNet_87), .D(n_3190), .Q(pZ_15_) );
NAND2_Z01 g60044 ( .a(n_856), .b(n_4604), .o(n_1086) );
AND2_X1 g60636 ( .a(n_292), .b(n_4529), .o(n_498) );
NAND2_Z01 g59505 ( .a(n_1537), .b(n_954), .o(n_1615) );
NAND3_Z1 g58453 ( .a(n_356), .b(n_2611), .c(n_41), .o(n_2642) );
NAND2_Z01 g59648 ( .a(n_1420), .b(n_1387), .o(n_1491) );
NOR2_Z4 g57760 ( .a(n_3108), .b(n_1579), .o(n_3115) );
fflopd pX_reg_7_ ( .CK(newNet_207), .D(n_3188), .Q(pX_7_) );
BUF_X2 newInst_1837 ( .a(newNet_1836), .o(newNet_1837) );
BUF_X2 newInst_1722 ( .a(newNet_477), .o(newNet_1722) );
BUF_X2 newInst_1585 ( .a(newNet_1584), .o(newNet_1585) );
NAND2_Z01 g60728 ( .a(n_257), .b(n_4486), .o(n_469) );
AND2_X1 g35224 ( .a(n_3357), .b(n_3231), .o(n_3445) );
XOR2_X1 g34354 ( .a(n_4151), .b(SP_5_), .o(n_4181) );
NAND2_Z01 g35402 ( .a(pY_4_), .b(pmem_d_11), .o(n_3307) );
NAND2_Z01 g57940 ( .a(n_2967), .b(n_2347), .o(n_3002) );
NAND2_Z01 g59159 ( .a(n_1894), .b(n_759), .o(n_1941) );
NAND2_Z01 g34805 ( .a(n_3575), .b(GPR_8__2_), .o(n_3758) );
BUF_X2 newInst_1658 ( .a(newNet_1657), .o(newNet_1658) );
NAND2_Z01 g34262 ( .a(n_4176), .b(pX_2_), .o(n_4271) );
BUF_X2 newInst_677 ( .a(newNet_676), .o(newNet_677) );
BUF_X2 newInst_1727 ( .a(newNet_1726), .o(newNet_1727) );
BUF_X2 newInst_1635 ( .a(newNet_1634), .o(newNet_1635) );
fflopd GPR_reg_23__3_ ( .CK(newNet_1045), .D(n_2847), .Q(GPR_23__3_) );
AND2_X1 g59016 ( .a(n_1984), .b(n_43), .o(n_2092) );
fflopd GPR_reg_6__2_ ( .CK(newNet_819), .D(n_2741), .Q(GPR_6__2_) );
NAND2_Z01 g58011 ( .a(n_2939), .b(n_24), .o(n_2985) );
NAND2_Z01 g59827 ( .a(n_1171), .b(dmem_di_6), .o(n_1297) );
NAND4_Z1 g57639 ( .a(n_1910), .b(n_1924), .c(n_3189), .d(n_1426), .o(n_3194) );
NOR2_Z1 g35085 ( .a(n_3484), .b(Rd_0_), .o(n_3509) );
NAND2_Z01 g34952 ( .a(n_3552), .b(GPR_3__4_), .o(n_3610) );
NAND2_Z01 g58999 ( .a(n_2015), .b(n_1892), .o(n_2108) );
BUF_X2 newInst_256 ( .a(newNet_255), .o(newNet_256) );
AND4_X1 g60127 ( .a(n_44), .b(n_250), .c(n_471), .d(n_36), .o(n_1035) );
NAND2_Z01 final_adder_mux_R16_278_6_g375 ( .a(final_adder_mux_R16_278_6_n_72), .b(final_adder_mux_R16_278_6_n_27), .o(final_adder_mux_R16_278_6_n_74) );
INV_X1 g35460 ( .a(SP_11_), .o(n_3264) );
BUF_X2 newInst_586 ( .a(newNet_315), .o(newNet_586) );
fflopd GPR_reg_9__7_ ( .CK(newNet_666), .D(n_3145), .Q(GPR_9__7_) );
XOR2_X1 g34461 ( .a(n_4058), .b(pZ_10_), .o(n_4081) );
XOR2_X1 final_adder_mux_R16_278_6_g370 ( .a(final_adder_mux_R16_278_6_n_77), .b(final_adder_mux_R16_278_6_n_31), .o(R16_12_) );
AND2_X1 g59475 ( .a(n_1622), .b(SP_13_), .o(n_1662) );
NAND2_Z01 g35278 ( .a(U_7_), .b(n_3275), .o(n_3397) );
BUF_X2 newInst_1494 ( .a(newNet_1493), .o(newNet_1494) );
NAND3_Z1 g60083 ( .a(n_539), .b(n_621), .c(n_699), .o(n_1053) );
INV_X2 newInst_1268 ( .a(newNet_291), .o(newNet_1268) );
NAND2_Z01 g59178 ( .a(n_1872), .b(n_1651), .o(n_1929) );
NAND2_Z01 g34174 ( .a(n_4325), .b(n_4470), .o(n_4341) );
NOR2_Z1 g60688 ( .a(n_197), .b(n_74), .o(n_450) );
fflopd GPR_reg_15__0_ ( .CK(newNet_1524), .D(n_2634), .Q(GPR_15__0_) );
BUF_X2 newInst_1022 ( .a(newNet_1021), .o(newNet_1022) );
BUF_X2 newInst_607 ( .a(newNet_606), .o(newNet_607) );
NAND2_Z01 g60446 ( .a(n_349), .b(pX_1_), .o(n_700) );
fflopd GPR_reg_16__3_ ( .CK(newNet_1461), .D(n_2859), .Q(GPR_16__3_) );
AND2_X1 g35163 ( .a(n_3442), .b(pZ_4_), .o(n_3466) );
BUF_X2 newInst_195 ( .a(newNet_194), .o(newNet_195) );
NAND2_Z01 g60879 ( .a(n_4683), .b(pmem_d_13), .o(n_245) );
NAND2_Z01 g60225 ( .a(n_600), .b(pX_0_), .o(n_920) );
NOR2_Z1 g59292 ( .a(n_853), .b(n_1765), .o(n_1818) );
NOR2_Z1 g59837 ( .a(n_1162), .b(n_62), .o(n_1288) );
NOR4_Z1 g35063 ( .a(n_3238), .b(n_3287), .c(n_4630), .d(pmem_d_0), .o(n_3523) );
BUF_X2 newInst_1608 ( .a(newNet_183), .o(newNet_1608) );
NOR2_Z1 g59682 ( .a(n_1329), .b(pmem_d_1), .o(n_1443) );
NAND2_Z01 g34820 ( .a(n_3586), .b(GPR_9__2_), .o(n_3743) );
BUF_X2 newInst_1448 ( .a(newNet_1447), .o(newNet_1448) );
BUF_X2 newInst_1380 ( .a(newNet_1379), .o(newNet_1380) );
NAND2_Z01 g58297 ( .a(n_2706), .b(n_2438), .o(n_2773) );
BUF_X2 newInst_429 ( .a(newNet_428), .o(newNet_429) );
XNOR2_X1 g59735 ( .a(n_1313), .b(pX_8_), .o(n_1395) );
fflopd U_reg_15_ ( .CK(newNet_397), .D(n_3184), .Q(U_15_) );
BUF_X2 newInst_1476 ( .a(newNet_1475), .o(newNet_1476) );
NAND2_Z01 g34106 ( .a(io_do_3), .b(n_4177), .o(n_4387) );
BUF_X2 newInst_1220 ( .a(newNet_1219), .o(newNet_1220) );
NAND2_Z01 g35263 ( .a(U_4_), .b(n_3275), .o(n_3409) );
BUF_X2 newInst_1245 ( .a(newNet_378), .o(newNet_1245) );
INV_X1 g61070 ( .a(pX_3_), .o(n_82) );
NAND2_Z01 g60917 ( .a(PC_2_), .b(pmem_d_2), .o(n_225) );
NAND4_Z1 g34571 ( .a(n_3832), .b(n_3829), .c(n_3831), .d(n_3830), .o(n_3989) );
NAND2_Z01 g34783 ( .a(n_3581), .b(GPR_16__3_), .o(n_3782) );
BUF_X2 newInst_479 ( .a(newNet_478), .o(newNet_479) );
AND3_X1 g58609 ( .a(n_1947), .b(n_2481), .c(n_1995), .o(n_2502) );
NAND2_Z01 g58061 ( .a(n_874), .b(n_2908), .o(n_2942) );
AND2_X1 g58516 ( .a(n_2567), .b(n_2200), .o(n_2580) );
NAND2_Z01 g58477 ( .a(n_2316), .b(n_2577), .o(n_2617) );
NAND2_Z01 g57933 ( .a(n_2974), .b(n_2417), .o(n_3012) );
BUF_X2 newInst_699 ( .a(newNet_166), .o(newNet_699) );
NAND2_Z01 g34767 ( .a(n_3586), .b(GPR_9__4_), .o(n_3798) );
INV_X1 g60091 ( .a(n_1036), .o(n_1037) );
BUF_X2 newInst_1680 ( .a(newNet_1679), .o(newNet_1680) );
BUF_X2 newInst_100 ( .a(newNet_14), .o(newNet_100) );
NOR2_Z2 g59245 ( .a(n_1829), .b(n_4610), .o(n_1871) );
NAND2_Z01 g34694 ( .a(n_3581), .b(GPR_16__6_), .o(n_3871) );
BUF_X2 newInst_523 ( .a(newNet_522), .o(newNet_523) );
AND2_X1 g59363 ( .a(n_1672), .b(n_1269), .o(n_1750) );
NAND2_Z01 g60453 ( .a(n_374), .b(GPR_12__0_), .o(n_693) );
NAND4_Z1 g58132 ( .a(n_1966), .b(n_2470), .c(n_2828), .d(n_2056), .o(n_2881) );
BUF_X2 newInst_683 ( .a(newNet_682), .o(newNet_683) );
fflopd GPR_reg_20__1_ ( .CK(newNet_1202), .D(n_2765), .Q(GPR_20__1_) );
NAND2_Z01 g34611 ( .a(n_3901), .b(n_3483), .o(n_3949) );
fflopd PC_reg_3_ ( .CK(newNet_630), .D(n_2172), .Q(PC_3_) );
BUF_X2 newInst_235 ( .a(newNet_191), .o(newNet_235) );
NAND2_Z01 g60117 ( .a(n_854), .b(n_352), .o(n_1040) );
BUF_X2 newInst_600 ( .a(newNet_599), .o(newNet_600) );
BUF_X2 newInst_1800 ( .a(newNet_1799), .o(newNet_1800) );
NAND2_Z01 g59562 ( .a(n_1528), .b(n_453), .o(n_1573) );
NAND2_Z01 g58793 ( .a(n_2199), .b(GPR_0__3_), .o(n_2307) );
NOR4_Z1 g59299 ( .a(n_1125), .b(n_1139), .c(n_1706), .d(n_1104), .o(n_1813) );
NAND2_Z01 g60497 ( .a(n_370), .b(GPR_20__3_), .o(n_649) );
INV_X1 drc_bufs61138 ( .a(n_1696), .o(n_30) );
NAND2_Z01 g60880 ( .a(pX_0_), .b(pX_1_), .o(n_279) );
NAND2_Z01 g59788 ( .a(n_1268), .b(n_1047), .o(n_1336) );
AND2_X1 g58372 ( .a(n_2657), .b(n_2213), .o(n_2699) );
INV_X1 g35234 ( .a(n_3420), .o(n_4595) );
NAND2_Z01 g57844 ( .a(n_3032), .b(n_2225), .o(n_3066) );
NOR2_Z1 g35243 ( .a(n_4660), .b(pmem_d_3), .o(n_3417) );
BUF_X2 newInst_118 ( .a(newNet_117), .o(newNet_118) );
NAND2_Z01 g60278 ( .a(R16_4_), .b(n_571), .o(n_868) );
XNOR2_X1 g34663 ( .a(n_3637), .b(pmem_d_13), .o(n_3902) );
fflopd io_sp_reg_4_ ( .CK(newNet_315), .D(n_548), .Q(io_sp_4_) );
NAND2_Z01 g59711 ( .a(n_1388), .b(n_41), .o(n_1421) );
AND2_X1 g60110 ( .a(n_4556), .b(n_839), .o(n_1042) );
NAND2_Z01 g58696 ( .a(n_2210), .b(GPR_1__3_), .o(n_2410) );
BUF_X2 newInst_279 ( .a(newNet_278), .o(newNet_279) );
BUF_X2 newInst_1665 ( .a(newNet_1664), .o(newNet_1665) );
INV_X2 g61081 ( .a(pmem_d_3), .o(n_71) );
NAND2_Z02 g58917 ( .a(n_2152), .b(n_1203), .o(n_2205) );
NOR2_Z1 g35214 ( .a(n_3334), .b(n_3331), .o(n_3436) );
NAND3_Z1 g58277 ( .a(n_1234), .b(n_2659), .c(n_1078), .o(n_2791) );
BUF_X2 newInst_1095 ( .a(newNet_1094), .o(newNet_1095) );
NOR2_Z1 g59432 ( .a(n_1630), .b(n_1619), .o(n_1687) );
NAND2_Z01 g60338 ( .a(n_25), .b(n_261), .o(n_792) );
NAND2_Z01 g34647 ( .a(n_3768), .b(n_4543), .o(n_3913) );
BUF_X2 newInst_1121 ( .a(newNet_1120), .o(newNet_1121) );
XNOR2_X1 g58454 ( .a(n_2603), .b(n_1769), .o(n_2655) );
BUF_X2 newInst_941 ( .a(newNet_940), .o(newNet_941) );
BUF_X1 mybuffer2 ( .o(io_a_2), .a(pmem_d_2) );
INV_X1 g61032 ( .a(pY_8_), .o(n_120) );
AND2_X1 g58957 ( .a(n_2086), .b(n_1210), .o(n_2144) );
NAND2_Z01 g34749 ( .a(n_3628), .b(GPR_19__5_), .o(n_3816) );
NAND2_Z01 g34898 ( .a(n_3633), .b(pZ_5_), .o(n_3665) );
INV_Z1 g16809 ( .a(GPR_12__7_), .o(n_4407) );
NAND2_Z01 g60312 ( .a(n_570), .b(pZ_0_), .o(n_814) );
NAND2_Z01 g34259 ( .a(n_4176), .b(pX_4_), .o(n_4274) );
NAND2_Z01 g34148 ( .a(n_4317), .b(n_4627), .o(n_4360) );
BUF_X2 newInst_1252 ( .a(newNet_1251), .o(newNet_1252) );
NAND4_Z1 g60372 ( .a(n_420), .b(n_421), .c(n_432), .d(n_435), .o(n_771) );
INV_X1 g35131 ( .a(n_3475), .o(n_4593) );
AND3_X1 g60845 ( .a(n_35), .b(T), .c(n_44), .o(n_293) );
BUF_X2 newInst_1475 ( .a(newNet_1474), .o(newNet_1475) );
NAND2_Z01 g60833 ( .a(n_167), .b(n_269), .o(n_298) );
BUF_X2 newInst_1732 ( .a(newNet_1731), .o(newNet_1732) );
BUF_X2 newInst_428 ( .a(newNet_427), .o(newNet_428) );
BUF_X2 newInst_1313 ( .a(newNet_1312), .o(newNet_1313) );
AND2_X1 g60107 ( .a(n_968), .b(n_966), .o(n_1044) );
NAND2_Z01 g58863 ( .a(n_2156), .b(GPR_15__2_), .o(n_2244) );
BUF_X2 newInst_1641 ( .a(newNet_1340), .o(newNet_1641) );
BUF_X2 newInst_1012 ( .a(newNet_1011), .o(newNet_1012) );
NAND2_Z01 g34777 ( .a(n_3579), .b(GPR_12__3_), .o(n_3788) );
BUF_X2 newInst_79 ( .a(newNet_10), .o(newNet_79) );
NAND2_Z01 g60437 ( .a(Rd_3_), .b(n_345), .o(n_709) );
BUF_X2 newInst_1491 ( .a(newNet_908), .o(newNet_1491) );
BUF_X2 newInst_1856 ( .a(newNet_1855), .o(newNet_1856) );
NOR2_Z1 g59021 ( .a(n_1972), .b(n_1920), .o(n_2081) );
BUF_X2 newInst_1508 ( .a(newNet_1507), .o(newNet_1508) );
NAND2_Z01 g57690 ( .a(n_3158), .b(n_2217), .o(n_3176) );
NAND2_Z01 g34698 ( .a(n_3566), .b(GPR_18__6_), .o(n_3867) );
BUF_X2 newInst_1378 ( .a(newNet_1377), .o(newNet_1378) );
INV_X1 g61055 ( .a(SP_7_), .o(n_97) );
BUF_X2 newInst_1045 ( .a(newNet_1044), .o(newNet_1045) );
NOR2_Z1 g61008 ( .a(n_4622), .b(pmem_d_2), .o(n_132) );
fflopd SP_reg_9_ ( .CK(newNet_465), .D(n_1636), .Q(SP_9_) );
BUF_X2 newInst_60 ( .a(newNet_59), .o(newNet_60) );
NAND2_Z01 g59480 ( .a(n_27), .b(n_71), .o(n_1645) );
NAND2_Z01 g58285 ( .a(n_2711), .b(n_2264), .o(n_2785) );
INV_X1 g60770 ( .a(n_376), .o(n_375) );
fflopd PC_reg_0_ ( .CK(newNet_660), .D(n_2179), .Q(PC_0_) );
NOR2_Z1 g60807 ( .a(n_170), .b(pmem_d_14), .o(n_311) );
NAND4_Z1 g59669 ( .a(n_1058), .b(n_1292), .c(n_1371), .d(n_1063), .o(n_1459) );
BUF_X2 newInst_1572 ( .a(newNet_1571), .o(newNet_1572) );
NAND2_Z01 final_adder_mux_R16_278_6_g366 ( .a(final_adder_mux_R16_278_6_n_81), .b(final_adder_mux_R16_278_6_n_15), .o(final_adder_mux_R16_278_6_n_83) );
NAND2_Z01 g58780 ( .a(n_2200), .b(GPR_7__0_), .o(n_2320) );
NAND2_Z01 g34297 ( .a(n_4102), .b(n_4158), .o(n_4237) );
NAND4_Z1 g34599 ( .a(n_3684), .b(n_3685), .c(n_3686), .d(n_3862), .o(n_3961) );
BUF_X2 newInst_1750 ( .a(newNet_1749), .o(newNet_1750) );
INV_X1 g61105 ( .a(pmem_d_4), .o(n_47) );
NAND2_Z01 g60185 ( .a(n_668), .b(n_667), .o(n_969) );
NAND2_Z01 g58686 ( .a(n_2211), .b(GPR_19__2_), .o(n_2420) );
NAND2_Z01 g34306 ( .a(n_4160), .b(n_4589), .o(n_4227) );
NOR2_Z1 g34298 ( .a(n_16064_BAR), .b(n_3929), .o(n_4236) );
NOR3_Z1 g60661 ( .a(n_275), .b(n_39083_BAR), .c(n_4536), .o(n_567) );
NOR2_Z1 g59650 ( .a(n_1416), .b(n_1410), .o(n_1488) );
NAND2_Z01 g58158 ( .a(n_2807), .b(n_2410), .o(n_2855) );
NAND2_Z01 g34916 ( .a(n_3633), .b(pZ_8_), .o(n_3647) );
NAND2_Z01 g58340 ( .a(n_2661), .b(n_2660), .o(n_2729) );
NAND2_Z01 g58597 ( .a(n_2458), .b(pX_10_), .o(n_2498) );
NAND2_Z01 g35310 ( .a(n_3289), .b(pY_9_), .o(n_3366) );
NAND2_Z01 g58872 ( .a(n_2158), .b(GPR_12__4_), .o(n_2235) );
NAND2_Z01 g60294 ( .a(R16_15_), .b(n_14), .o(n_830) );
BUF_X2 newInst_1818 ( .a(newNet_1817), .o(newNet_1818) );
BUF_X2 newInst_619 ( .a(newNet_618), .o(newNet_619) );
BUF_X2 newInst_16 ( .a(newNet_15), .o(newNet_16) );
NAND2_Z01 g58886 ( .a(n_2140), .b(GPR_9__2_), .o(n_2221) );
INV_X1 g60779 ( .a(n_327), .o(n_328) );
NAND2_Z01 g59922 ( .a(n_1026), .b(T), .o(n_1219) );
NAND2_Z01 g34709 ( .a(n_3628), .b(GPR_19__6_), .o(n_3856) );
NAND2_Z01 g58782 ( .a(n_2200), .b(GPR_7__2_), .o(n_2318) );
NAND2_Z01 g60546 ( .a(n_368), .b(GPR_13__7_), .o(n_560) );
NOR4_Z1 g60162 ( .a(n_502), .b(n_526), .c(n_506), .d(n_317), .o(n_974) );
AND2_X1 g58251 ( .a(n_2752), .b(n_2139), .o(n_2816) );
NAND2_Z01 g58164 ( .a(n_2802), .b(n_2369), .o(n_2846) );
NOR3_Z1 g34491 ( .a(n_4011), .b(n_3997), .c(n_4024), .o(n_4053) );
BUF_X2 newInst_37 ( .a(newNet_11), .o(newNet_37) );
NOR2_Z1 g58341 ( .a(n_2688), .b(n_1732), .o(n_2728) );
NAND2_Z01 g60478 ( .a(Rd_3_), .b(n_340), .o(n_668) );
BUF_X2 newInst_1330 ( .a(newNet_1329), .o(newNet_1330) );
NAND2_Z01 g58700 ( .a(n_2213), .b(GPR_17__4_), .o(n_2406) );
NAND2_Z01 g58048 ( .a(n_2897), .b(n_2400), .o(n_2934) );
NAND2_Z01 g57845 ( .a(n_3031), .b(n_2190), .o(n_3065) );
BUF_X2 newInst_613 ( .a(newNet_612), .o(newNet_613) );
NOR2_Z1 g34281 ( .a(n_4613), .b(n_3223), .o(n_4252) );
NAND2_Z01 g59623 ( .a(n_1414), .b(io_di_5), .o(n_1504) );
NOR2_Z1 g60815 ( .a(n_177), .b(n_4533), .o(n_309) );
INV_X1 drc_bufs61207 ( .a(n_462), .o(n_22) );
fflopd SP_reg_5_ ( .CK(newNet_489), .D(n_1740), .Q(SP_5_) );
INV_X1 g61064 ( .a(pY_12_), .o(n_88) );
fflopd GPR_reg_18__1_ ( .CK(newNet_1362), .D(n_2770), .Q(GPR_18__1_) );
BUF_X2 newInst_207 ( .a(newNet_206), .o(newNet_207) );
NOR2_Z1 g60327 ( .a(n_521), .b(n_116), .o(n_801) );
NAND2_Z01 g58332 ( .a(n_2663), .b(n_2309), .o(n_2733) );
NAND2_Z01 g58794 ( .a(n_2199), .b(GPR_0__4_), .o(n_2306) );
NAND2_Z01 g60781 ( .a(n_178), .b(n_118), .o(n_321) );
AND2_X1 g58110 ( .a(n_2850), .b(n_2214), .o(n_2902) );
BUF_X2 newInst_1681 ( .a(newNet_1680), .o(newNet_1681) );
NOR2_Z1 g34316 ( .a(n_4159), .b(n_4029), .o(n_4217) );
fflopd GPR_reg_12__3_ ( .CK(newNet_1645), .D(n_2863), .Q(GPR_12__3_) );
BUF_X2 newInst_459 ( .a(newNet_458), .o(newNet_459) );
NAND2_Z01 g59340 ( .a(n_1692), .b(pmem_d_9), .o(n_1801) );
BUF_X2 newInst_649 ( .a(newNet_648), .o(newNet_649) );
NAND2_Z01 g60715 ( .a(GPR_7__7_), .b(n_183), .o(n_423) );
NAND2_Z01 g35351 ( .a(n_3281), .b(n_3307), .o(n_3329) );
AND2_X1 g60982 ( .a(n_4620), .b(pmem_d_3), .o(n_186) );
NAND2_Z02 g58916 ( .a(n_2160), .b(n_1202), .o(n_2206) );
BUF_X2 newInst_1339 ( .a(newNet_1251), .o(newNet_1339) );
BUF_X2 newInst_864 ( .a(newNet_863), .o(newNet_864) );
BUF_X2 newInst_1371 ( .a(newNet_849), .o(newNet_1371) );
AND2_X1 g58362 ( .a(n_2656), .b(n_2158), .o(n_2709) );
BUF_X2 newInst_1145 ( .a(newNet_1144), .o(newNet_1145) );
BUF_X2 newInst_955 ( .a(newNet_954), .o(newNet_955) );
NAND2_Z01 g60341 ( .a(n_11), .b(pmem_d_9), .o(n_789) );
NAND2_Z01 g60564 ( .a(n_341), .b(pY_3_), .o(n_544) );
NOR2_Z2 g59227 ( .a(n_1829), .b(n_4613), .o(n_1894) );
NOR4_Z1 g34456 ( .a(n_3777), .b(n_3978), .c(n_4049), .d(n_3653), .o(n_4086) );
NAND2_Z01 g59462 ( .a(n_1613), .b(n_1425), .o(n_1659) );
fflopd GPR_reg_16__5_ ( .CK(newNet_1441), .D(n_3015), .Q(GPR_16__5_) );
BUF_X2 newInst_520 ( .a(newNet_519), .o(newNet_520) );
NAND2_Z01 g58859 ( .a(n_2156), .b(GPR_15__1_), .o(n_2248) );
BUF_X2 newInst_1662 ( .a(newNet_1661), .o(newNet_1662) );
AND2_X1 g58126 ( .a(n_2850), .b(n_2153), .o(n_2886) );
NOR2_Z1 g35339 ( .a(n_4514), .b(n_3237), .o(n_4526) );
BUF_X2 newInst_1435 ( .a(newNet_1434), .o(newNet_1435) );
NAND2_Z01 g58244 ( .a(n_2753), .b(n_2215), .o(n_2823) );
INV_X1 g34518 ( .a(n_4646), .o(n_4025) );
AND2_X1 g34286 ( .a(n_4613), .b(n_4597), .o(n_4247) );
INV_X1 g59308 ( .a(n_1805), .o(n_1806) );
NAND4_Z1 g59664 ( .a(n_808), .b(n_916), .c(n_1360), .d(n_925), .o(n_1463) );
BUF_X2 newInst_404 ( .a(newNet_403), .o(newNet_404) );
fflopd pX_reg_9_ ( .CK(newNet_200), .D(n_2880), .Q(pX_9_) );
BUF_X2 newInst_966 ( .a(newNet_965), .o(newNet_966) );
XOR2_X1 g60388 ( .a(n_302), .b(n_270), .o(n_758) );
NAND4_Z1 g57812 ( .a(n_1950), .b(n_2517), .c(n_3062), .d(n_1952), .o(n_3095) );
NAND2_Z01 g58892 ( .a(n_2140), .b(GPR_9__6_), .o(n_2190) );
NAND2_Z03 g34170 ( .a(n_4315), .b(n_3953), .o(io_do_0) );
BUF_X2 newInst_1661 ( .a(newNet_1660), .o(newNet_1661) );
NAND2_Z01 final_adder_mux_R16_278_6_g431 ( .a(n_4439), .b(n_4423), .o(final_adder_mux_R16_278_6_n_18) );
INV_X1 g60532 ( .a(n_604), .o(n_605) );
INV_X1 g35504 ( .a(pY_6_), .o(n_3223) );
INV_X1 g61096 ( .a(n_4652), .o(n_56) );
NAND2_Z01 g60961 ( .a(n_62), .b(pmem_d_2), .o(n_202) );
NAND2_Z01 g57716 ( .a(n_3126), .b(n_2374), .o(n_3151) );
NAND2_Z01 g58853 ( .a(n_2157), .b(GPR_13__0_), .o(n_2254) );
INV_X1 g61092 ( .a(dmem_di_1), .o(n_60) );
NAND2_Z01 g34985 ( .a(n_3551), .b(n_3461), .o(n_3598) );
NAND2_Z01 g35401 ( .a(pY_3_), .b(pmem_d_10), .o(n_3308) );
BUF_X2 newInst_48 ( .a(newNet_12), .o(newNet_48) );
NAND2_Z01 g59229 ( .a(n_1834), .b(n_1823), .o(n_1891) );
BUF_X2 newInst_817 ( .a(newNet_816), .o(newNet_817) );
NAND3_Z1 g58568 ( .a(n_1976), .b(n_2506), .c(n_2001), .o(n_2530) );
NAND3_Z1 g60792 ( .a(n_4516), .b(n_4515), .c(n_78), .o(n_373) );
NAND2_Z01 g59315 ( .a(n_1720), .b(n_1088), .o(n_1798) );
NAND4_Z1 g57655 ( .a(n_1986), .b(n_2518), .c(n_3178), .d(n_2043), .o(n_3187) );
AND2_X1 final_adder_mux_R16_278_6_g448 ( .a(n_4439), .b(n_4423), .o(final_adder_mux_R16_278_6_n_1) );
NOR2_Z1 g60628 ( .a(n_458), .b(n_199), .o(n_582) );
BUF_X2 newInst_301 ( .a(newNet_300), .o(newNet_301) );
BUF_X2 newInst_55 ( .a(newNet_54), .o(newNet_55) );
NAND2_Z01 g60344 ( .a(n_11), .b(pmem_d_1), .o(n_787) );
BUF_X2 newInst_6 ( .a(newNet_3), .o(newNet_6) );
AND3_X1 g59200 ( .a(n_1806), .b(n_1826), .c(pmem_d_7), .o(n_1910) );
BUF_X2 newInst_623 ( .a(newNet_622), .o(newNet_623) );
NOR2_Z1 g35268 ( .a(n_3312), .b(n_3257), .o(n_3415) );
NAND2_Z01 g35410 ( .a(pZ_4_), .b(pmem_d_11), .o(n_3294) );
NOR4_Z1 g58930 ( .a(n_1887), .b(n_1460), .c(n_1331), .d(n_1932), .o(n_2175) );
BUF_X2 newInst_734 ( .a(newNet_733), .o(newNet_734) );
NAND2_Z01 g34331 ( .a(n_4160), .b(n_4594), .o(n_4203) );
BUF_X2 newInst_267 ( .a(newNet_266), .o(newNet_267) );
BUF_X2 newInst_606 ( .a(newNet_605), .o(newNet_606) );
XOR2_X1 g60382 ( .a(n_362), .b(n_86), .o(n_763) );
BUF_X2 newInst_1772 ( .a(newNet_397), .o(newNet_1772) );
BUF_X2 newInst_1584 ( .a(newNet_1583), .o(newNet_1584) );
NAND2_Z01 g60504 ( .a(n_21), .b(Rd_r_0_), .o(n_642) );
BUF_X2 newInst_1755 ( .a(newNet_1754), .o(newNet_1755) );
BUF_X2 newInst_1282 ( .a(newNet_1281), .o(newNet_1282) );
NOR2_Z1 g35153 ( .a(n_3452), .b(n_3211), .o(n_3470) );
NOR2_Z1 g59955 ( .a(n_979), .b(n_1051), .o(n_1176) );
AND2_X1 g59167 ( .a(n_1867), .b(n_4640), .o(n_1979) );
NAND2_Z01 g35417 ( .a(pY_0_), .b(pmem_d_0), .o(n_3301) );
AND3_X1 g59534 ( .a(n_850), .b(n_1483), .c(io_do_3), .o(n_1593) );
NAND2_Z01 g34678 ( .a(n_3631), .b(GPR_11__7_), .o(n_3887) );
INV_X2 newInst_93 ( .a(newNet_92), .o(newNet_93) );
AND3_X1 g60369 ( .a(n_118), .b(n_369), .c(SP_3_), .o(n_772) );
BUF_X2 newInst_347 ( .a(newNet_346), .o(newNet_347) );
NAND2_Z01 g34726 ( .a(n_3586), .b(GPR_8__5_), .o(n_3839) );
NAND2_Z01 g60557 ( .a(n_393), .b(n_395), .o(n_549) );
NOR2_Z1 g35062 ( .a(n_3506), .b(pY_7_), .o(n_4517) );
BUF_X2 newInst_1831 ( .a(newNet_1830), .o(newNet_1831) );
NAND2_Z01 g58672 ( .a(n_2214), .b(GPR_16__6_), .o(n_2434) );
NAND2_Z01 g60892 ( .a(n_4667), .b(n_32), .o(n_236) );
NAND2_Z01 g59062 ( .a(n_1902), .b(n_4592), .o(n_2045) );
AND2_X1 g58009 ( .a(n_2940), .b(n_2153), .o(n_2962) );
AND2_X1 g58949 ( .a(n_2103), .b(pX_15_), .o(n_2149) );
NAND4_Z1 g58020 ( .a(n_1907), .b(n_2525), .c(n_2911), .d(n_2018), .o(n_2952) );
BUF_X2 newInst_1794 ( .a(newNet_464), .o(newNet_1794) );
NAND3_Z1 g58348 ( .a(n_1277), .b(n_2642), .c(n_522), .o(n_2722) );
NAND2_Z01 g58803 ( .a(n_2197), .b(U_1_), .o(n_2297) );
NAND2_Z01 g34826 ( .a(n_3625), .b(GPR_1__1_), .o(n_3737) );
BUF_X2 newInst_1325 ( .a(newNet_1324), .o(newNet_1325) );
AND4_X1 g34062 ( .a(n_4147), .b(n_4234), .c(n_4399), .d(n_4132), .o(dmem_a_12) );
INV_X1 g60286 ( .a(n_769), .o(n_840) );
NAND3_Z1 g59896 ( .a(io_do_5), .b(n_1026), .c(n_344), .o(n_1233) );
NAND2_Z01 g34674 ( .a(n_3603), .b(n_3604), .o(n_3891) );
NAND2_Z01 g60098 ( .a(n_774), .b(n_32), .o(n_1021) );
INV_X1 g59709 ( .a(n_1416), .o(n_1417) );
fflopd pY_reg_8_ ( .CK(newNet_126), .D(n_2724), .Q(pY_8_) );
NAND2_Z01 g34942 ( .a(n_3551), .b(GPR_4__6_), .o(n_3620) );
BUF_X2 newInst_1030 ( .a(newNet_1029), .o(newNet_1030) );
fflopd SP_reg_1_ ( .CK(newNet_524), .D(n_1578), .Q(SP_1_) );
NAND2_Z01 g61019 ( .a(n_86), .b(n_71), .o(n_127) );
BUF_X2 newInst_1579 ( .a(newNet_577), .o(newNet_1579) );
NOR4_Z1 g34233 ( .a(n_4195), .b(n_4199), .c(n_4241), .d(n_4109), .o(n_4298) );
BUF_X2 newInst_435 ( .a(newNet_434), .o(newNet_435) );
BUF_X2 newInst_465 ( .a(newNet_464), .o(newNet_465) );
BUF_X2 newInst_70 ( .a(newNet_69), .o(newNet_70) );
NAND2_Z01 g34139 ( .a(n_4325), .b(n_4621), .o(n_4369) );
NAND2_Z01 g58752 ( .a(n_2204), .b(GPR_3__4_), .o(n_2348) );
NOR3_Z1 g60850 ( .a(n_4686), .b(n_276), .c(n_4659), .o(n_335) );
INV_X1 g59234 ( .a(n_1875), .o(n_1874) );
fflopd GPR_Rd_r_reg_5_ ( .CK(newNet_1844), .D(io_do_5), .Q(GPR_Rd_r_5_) );
AND2_X1 final_adder_mux_R16_278_6_g443 ( .a(n_4437), .b(n_4421), .o(final_adder_mux_R16_278_6_n_6) );
INV_X1 g58889 ( .a(n_2196), .o(n_2195) );
fflopd GPR_reg_19__0_ ( .CK(newNet_1325), .D(n_2631), .Q(GPR_19__0_) );
NAND4_Z1 g34581 ( .a(n_3780), .b(n_3781), .c(n_3783), .d(n_3782), .o(n_3979) );
AND2_X1 g60759 ( .a(n_259), .b(n_63), .o(n_463) );
NOR2_Z1 g60999 ( .a(io_do_7), .b(pmem_d_11), .o(n_139) );
AND2_X1 g34489 ( .a(n_4038), .b(n_3306), .o(n_4057) );
fflopd GPR_reg_5__2_ ( .CK(newNet_862), .D(n_2743), .Q(GPR_5__2_) );
NAND2_Z01 g58050 ( .a(n_2895), .b(n_2384), .o(n_2932) );
NAND2_Z01 g59099 ( .a(n_1894), .b(n_1220), .o(n_2009) );
NOR2_Z1 g34391 ( .a(n_4089), .b(n_3226), .o(n_4147) );
NAND2_Z01 g34665 ( .a(n_3620), .b(n_3621), .o(n_3900) );
NOR2_Z1 g58561 ( .a(n_2486), .b(n_2277), .o(n_2537) );
NAND3_Z1 g59801 ( .a(n_1169), .b(n_1152), .c(n_794), .o(n_1326) );
INV_X1 g59676 ( .a(n_1448), .o(n_1449) );
NAND4_Z1 g34250 ( .a(n_3890), .b(n_3938), .c(n_4150), .d(n_3889), .o(n_4283) );
NAND2_Z01 g60026 ( .a(n_4602), .b(n_856), .o(n_1103) );
BUF_X2 newInst_1402 ( .a(newNet_1401), .o(newNet_1402) );
BUF_X2 newInst_1273 ( .a(newNet_1272), .o(newNet_1273) );
NOR2_Z1 g60648 ( .a(n_354), .b(pY_13_), .o(n_572) );
BUF_X2 newInst_712 ( .a(newNet_711), .o(newNet_712) );
NAND4_Z1 g58545 ( .a(n_1598), .b(n_2452), .c(n_2509), .d(n_1432), .o(n_2553) );
NAND2_Z01 g59753 ( .a(n_1312), .b(io_do_3), .o(n_1371) );
NAND2_Z01 g60305 ( .a(n_597), .b(pX_8_), .o(n_819) );
NOR2_Z1 g59781 ( .a(n_1309), .b(SP_8_), .o(n_1351) );
NAND2_Z01 g60760 ( .a(n_251), .b(pmem_d_2), .o(n_462) );
AND2_X1 g61012 ( .a(n_4447), .b(n_4431), .o(n_169) );
NOR2_Z1 g35173 ( .a(n_3419), .b(n_3220), .o(n_4664) );
AND2_X1 g59444 ( .a(n_1637), .b(n_1133), .o(n_1695) );
NOR4_Z1 g58411 ( .a(n_2534), .b(n_2606), .c(n_2065), .d(n_1255), .o(n_2659) );
NAND2_Z01 g58035 ( .a(n_2912), .b(n_2295), .o(n_2950) );
NAND2_Z01 g60243 ( .a(n_574), .b(GPR_10__5_), .o(n_902) );
NOR2_Z1 g60116 ( .a(n_4651), .b(n_775), .o(n_1010) );
fflopd GPR_reg_16__4_ ( .CK(newNet_1451), .D(n_2943), .Q(GPR_16__4_) );
BUF_X2 newInst_970 ( .a(newNet_969), .o(newNet_970) );
NAND2_Z01 g34155 ( .a(n_4317), .b(n_4620), .o(n_4353) );
fflopd SP_reg_2_ ( .CK(newNet_514), .D(n_1632), .Q(SP_2_) );
NAND2_Z01 g60527 ( .a(n_21), .b(Rd_r_4_), .o(n_619) );
BUF_X2 newInst_1357 ( .a(newNet_1356), .o(newNet_1357) );
BUF_X2 newInst_1569 ( .a(newNet_1568), .o(newNet_1569) );
BUF_X2 newInst_1786 ( .a(newNet_1785), .o(newNet_1786) );
NAND2_Z01 g59095 ( .a(n_1875), .b(n_373), .o(n_2013) );
XOR2_X1 g35198 ( .a(n_3355), .b(n_3245), .o(n_4607) );
NOR2_Z1 g34186 ( .a(n_4324), .b(n_4627), .o(n_4427) );
BUF_X2 newInst_932 ( .a(newNet_931), .o(newNet_932) );
NAND2_Z01 g58706 ( .a(n_2209), .b(GPR_20__3_), .o(n_2401) );
NOR2_Z1 g34410 ( .a(n_4610), .b(n_3767), .o(n_4128) );
BUF_X2 newInst_1117 ( .a(newNet_1116), .o(newNet_1117) );
NOR2_Z1 g59175 ( .a(n_1873), .b(n_466), .o(n_1931) );
NAND2_Z01 g34651 ( .a(n_3768), .b(n_4551), .o(n_3909) );
BUF_X2 newInst_1624 ( .a(newNet_1623), .o(newNet_1624) );
BUF_X2 newInst_961 ( .a(newNet_734), .o(newNet_961) );
BUF_X2 newInst_1634 ( .a(newNet_1633), .o(newNet_1634) );
INV_X1 g60281 ( .a(n_856), .o(n_855) );
NAND2_Z01 g34702 ( .a(n_3579), .b(GPR_12__6_), .o(n_3863) );
NAND2_Z01 g59704 ( .a(io_do_4), .b(n_1384), .o(n_1426) );
BUF_X2 newInst_1342 ( .a(newNet_1341), .o(newNet_1342) );
NAND2_Z01 g57827 ( .a(n_3049), .b(n_2247), .o(n_3086) );
NOR2_Z1 g35338 ( .a(n_3237), .b(n_3309), .o(n_3332) );
BUF_X2 newInst_894 ( .a(newNet_893), .o(newNet_894) );
NAND2_Z01 g34748 ( .a(n_3594), .b(GPR_7__5_), .o(n_3817) );
INV_X1 g61119 ( .a(n_4685), .o(n_33) );
NOR2_Z1 g59004 ( .a(n_1969), .b(n_1923), .o(n_2103) );
fflopd GPR_reg_3__6_ ( .CK(newNet_936), .D(n_3071), .Q(GPR_3__6_) );
BUF_X2 newInst_158 ( .a(newNet_95), .o(newNet_158) );
INV_X1 g35468 ( .a(pZ_5_), .o(n_3256) );
NAND2_Z01 g59115 ( .a(n_1884), .b(n_1036), .o(n_1994) );
fflopd state_reg_3_ ( .CK(newNet_1596), .D(n_2645), .Q(state_3_) );
NAND2_Z01 g60351 ( .a(n_178), .b(n_567), .o(n_858) );
NOR2_Z1 g59876 ( .a(n_1024), .b(n_1166), .o(n_1251) );
INV_X1 g61043 ( .a(SP_4_), .o(n_109) );
NAND2_Z01 g60036 ( .a(n_771), .b(n_377), .o(n_1094) );
BUF_X2 newInst_1847 ( .a(newNet_1846), .o(newNet_1847) );
NOR2_Z1 g60605 ( .a(n_458), .b(n_250), .o(n_597) );
NAND2_Z01 g59216 ( .a(n_1832), .b(n_1083), .o(n_1889) );
BUF_X2 newInst_1814 ( .a(newNet_1813), .o(newNet_1814) );
BUF_X2 newInst_1176 ( .a(newNet_1175), .o(newNet_1176) );
BUF_X2 newInst_1291 ( .a(newNet_1290), .o(newNet_1291) );
NAND2_Z01 g57987 ( .a(n_2942), .b(n_2193), .o(n_2984) );
NOR3_Z1 g58987 ( .a(n_1756), .b(n_1991), .c(n_1799), .o(n_2120) );
BUF_X2 newInst_1423 ( .a(newNet_1422), .o(newNet_1423) );
INV_X1 g35489 ( .a(pmem_d_2), .o(n_3236) );
AND2_X1 g58109 ( .a(n_2850), .b(n_2156), .o(n_2903) );
NOR2_Z1 g35160 ( .a(n_3201), .b(n_3225), .o(Rd_1_) );
BUF_X2 newInst_1186 ( .a(newNet_1185), .o(newNet_1186) );
NOR4_Z1 g34212 ( .a(n_3961), .b(n_3962), .c(n_4283), .d(n_3950), .o(n_4314) );
BUF_X2 newInst_1349 ( .a(newNet_1348), .o(newNet_1349) );
NAND2_Z01 g60487 ( .a(Rd_2_), .b(n_340), .o(n_659) );
BUF_X2 newInst_983 ( .a(newNet_982), .o(newNet_983) );
NAND2_Z01 g34795 ( .a(n_3585), .b(GPR_13__3_), .o(n_3770) );
INV_X1 g34482 ( .a(n_4059), .o(n_4060) );
BUF_X2 newInst_511 ( .a(newNet_510), .o(newNet_511) );
XOR2_X1 final_adder_mux_R16_278_6_g411 ( .a(n_4448), .b(n_4432), .o(final_adder_mux_R16_278_6_n_38) );
BUF_X2 newInst_1441 ( .a(newNet_1440), .o(newNet_1441) );
NAND2_Z01 final_adder_mux_R16_278_6_g384 ( .a(final_adder_mux_R16_278_6_n_63), .b(final_adder_mux_R16_278_6_n_19), .o(final_adder_mux_R16_278_6_n_65) );
NAND2_Z01 g57927 ( .a(n_2980), .b(n_2250), .o(n_3018) );
BUF_X2 newInst_1028 ( .a(newNet_356), .o(newNet_1028) );
NAND2_Z01 g58739 ( .a(n_2205), .b(GPR_2__4_), .o(n_2368) );
NAND2_Z01 g59400 ( .a(n_1657), .b(n_208), .o(n_1736) );
AND2_X1 g34470 ( .a(n_4058), .b(n_3237), .o(n_4073) );
AND3_X1 g60146 ( .a(n_4534), .b(n_858), .c(SP_10_), .o(n_986) );
INV_X1 drc_bufs61217 ( .a(n_566), .o(n_23) );
NAND4_Z1 g59996 ( .a(n_919), .b(n_888), .c(n_807), .d(n_920), .o(n_1133) );
BUF_X2 newInst_625 ( .a(newNet_534), .o(newNet_625) );
NAND2_Z01 g60255 ( .a(R16_2_), .b(n_571), .o(n_891) );
NAND2_Z01 g60270 ( .a(n_575), .b(GPR_2__5_), .o(n_876) );
AND3_X1 g35373 ( .a(pX_9_), .b(pX_8_), .c(pX_11_), .o(n_3317) );
INV_X1 g35475 ( .a(pmem_d_0), .o(n_3249) );
NAND2_Z01 g34961 ( .a(n_3541), .b(n_4628), .o(n_3601) );
XOR2_X1 g35381 ( .a(pZ_1_), .b(pZ_0_), .o(n_4609) );
BUF_X2 newInst_708 ( .a(newNet_707), .o(newNet_708) );
XOR2_X1 g59597 ( .a(n_1391), .b(n_47), .o(n_1532) );
NAND2_Z01 g34446 ( .a(n_4067), .b(n_3416), .o(dmem_we) );
BUF_X2 newInst_389 ( .a(newNet_388), .o(newNet_389) );
NAND2_Z01 g34525 ( .a(n_3670), .b(n_3944), .o(n_4019) );
NAND4_Z1 g34075 ( .a(n_3413), .b(n_3426), .c(n_4342), .d(n_3412), .o(n_4397) );
BUF_X2 newInst_653 ( .a(newNet_652), .o(newNet_653) );
BUF_X2 newInst_310 ( .a(newNet_309), .o(newNet_310) );
AND2_X1 g60078 ( .a(n_848), .b(n_71), .o(n_1057) );
BUF_X2 newInst_931 ( .a(newNet_930), .o(newNet_931) );
BUF_X2 newInst_393 ( .a(newNet_14), .o(newNet_393) );
AND2_X1 g58389 ( .a(n_2656), .b(n_2205), .o(n_2679) );
BUF_X2 newInst_115 ( .a(newNet_114), .o(newNet_115) );
AND2_X1 g61009 ( .a(n_4441), .b(n_4425), .o(n_131) );
NAND2_Z01 g60198 ( .a(R16_0_), .b(n_571), .o(n_947) );
AND2_X1 g61002 ( .a(n_4629), .b(pmem_d_9), .o(n_137) );
BUF_X2 newInst_531 ( .a(newNet_530), .o(newNet_531) );
NAND2_Z01 g60513 ( .a(n_374), .b(GPR_12__6_), .o(n_633) );
NAND2_Z01 g59865 ( .a(n_474), .b(n_1167), .o(n_1261) );
NAND4_Z1 g34591 ( .a(n_3722), .b(n_3721), .c(n_3737), .d(n_3720), .o(n_3969) );
BUF_X2 newInst_1411 ( .a(newNet_897), .o(newNet_1411) );
NAND4_Z1 g59378 ( .a(n_1478), .b(n_1003), .c(n_1656), .d(n_1338), .o(n_1740) );
NAND2_Z01 g59138 ( .a(n_1872), .b(n_1395), .o(n_1960) );
INV_X1 drc_bufs61137 ( .a(n_30), .o(n_15) );
NAND2_Z01 g60764 ( .a(n_201), .b(pmem_d_1), .o(n_459) );
NAND2_Z01 g60230 ( .a(R16_7_), .b(n_14), .o(n_915) );
NAND2_Z01 g58300 ( .a(n_2698), .b(n_2429), .o(n_2770) );
fflopd GPR_reg_23__7_ ( .CK(newNet_1027), .D(n_3151), .Q(GPR_23__7_) );
NAND2_Z01 g60943 ( .a(io_do_5), .b(n_59), .o(n_208) );
NAND2_Z01 g58554 ( .a(n_2492), .b(pZ_11_), .o(n_2543) );
BUF_X2 newInst_1670 ( .a(newNet_1669), .o(newNet_1670) );
NAND2_Z01 g35277 ( .a(U_14_), .b(n_3275), .o(n_3398) );
NAND2_Z02 g60937 ( .a(pmem_d_9), .b(pmem_d_3), .o(n_250) );
NAND2_Z01 g60930 ( .a(pmem_d_2), .b(pmem_d_0), .o(n_258) );
INV_X1 drc_bufs35551 ( .a(n_4618), .o(n_3204) );
INV_Z1 g16804 ( .a(GPR_20__6_), .o(n_4400) );
fflopd GPR_reg_18__3_ ( .CK(newNet_1350), .D(n_2857), .Q(GPR_18__3_) );
NAND2_Z01 g34219 ( .a(n_4164), .b(GPR_Rd_r_5_), .o(n_4308) );
NAND2_Z01 g34844 ( .a(n_3197), .b(GPR_23__1_), .o(n_3719) );
BUF_X2 newInst_1262 ( .a(newNet_1261), .o(newNet_1262) );
AND2_X1 g58960 ( .a(n_1625), .b(n_2082), .o(n_2143) );
NOR2_Z1 g59722 ( .a(n_1269), .b(n_1352), .o(n_1405) );
NAND2_Z01 g57833 ( .a(n_3043), .b(n_2407), .o(n_3077) );
NAND4_Z1 g34244 ( .a(n_3679), .b(n_3779), .c(n_4171), .d(n_3778), .o(n_4289) );
BUF_X2 newInst_1778 ( .a(newNet_1777), .o(newNet_1778) );
XOR2_X1 final_adder_mux_R16_278_6_g418 ( .a(n_4439), .b(n_4423), .o(final_adder_mux_R16_278_6_n_31) );
NAND2_Z01 g35284 ( .a(n_3299), .b(pX_15_), .o(n_3391) );
BUF_X2 newInst_471 ( .a(newNet_470), .o(newNet_471) );
fflopd GPR_reg_15__6_ ( .CK(newNet_1490), .D(n_3085), .Q(GPR_15__6_) );
BUF_X2 newInst_346 ( .a(newNet_345), .o(newNet_346) );
NAND2_Z01 g60685 ( .a(n_178), .b(n_4536), .o(n_453) );
BUF_X2 newInst_529 ( .a(newNet_528), .o(newNet_529) );
BUF_X2 newInst_325 ( .a(newNet_324), .o(newNet_325) );
BUF_X2 newInst_1711 ( .a(newNet_961), .o(newNet_1711) );
AND2_X1 g61024 ( .a(n_4556), .b(n_4641), .o(n_161) );
AND2_X1 g60743 ( .a(n_124), .b(n_250), .o(n_398) );
NAND2_Z01 g59354 ( .a(n_960), .b(n_1695), .o(n_1759) );
NAND2_Z01 final_adder_mux_R16_278_6_g372 ( .a(final_adder_mux_R16_278_6_n_75), .b(final_adder_mux_R16_278_6_n_24), .o(final_adder_mux_R16_278_6_n_77) );
NOR2_Z1 g58826 ( .a(n_2193), .b(n_1975), .o(n_2352) );
NAND2_Z01 g59917 ( .a(n_1085), .b(n_1084), .o(n_1196) );
NOR4_Z1 g58543 ( .a(n_1459), .b(n_2487), .c(n_2094), .d(n_2119), .o(n_2555) );
NAND2_Z01 g58235 ( .a(n_2755), .b(n_2218), .o(n_2832) );
NAND2_Z01 g34541 ( .a(n_3923), .b(n_3910), .o(pmem_a_3) );
XOR2_X1 g35020 ( .a(n_3513), .b(pZ_3_), .o(n_3556) );
NAND2_Z01 g60217 ( .a(R16_3_), .b(n_571), .o(n_928) );
BUF_X2 newInst_412 ( .a(newNet_411), .o(newNet_412) );
BUF_X2 newInst_1055 ( .a(newNet_1054), .o(newNet_1055) );
INV_X1 g58161 ( .a(n_2850), .o(n_2849) );
BUF_X2 newInst_44 ( .a(newNet_43), .o(newNet_44) );
NOR2_Z1 g34403 ( .a(n_4611), .b(n_3237), .o(n_4135) );
NAND3_Y1 g34435 ( .a(n_3448), .b(n_4065), .c(n_3426), .o(n_4125) );
NOR2_Z1 g34409 ( .a(n_4091), .b(n_3993), .o(n_4129) );
NAND2_Z01 g59685 ( .a(n_1350), .b(n_1192), .o(n_1451) );
NOR2_Z1 g58395 ( .a(n_2644), .b(n_1620), .o(n_2673) );
BUF_X2 newInst_850 ( .a(newNet_849), .o(newNet_850) );
NAND2_Z01 g34320 ( .a(n_4165), .b(n_4537), .o(n_4213) );
BUF_X2 newInst_1530 ( .a(newNet_1529), .o(newNet_1530) );
BUF_X2 newInst_503 ( .a(newNet_502), .o(newNet_503) );
fflopd pZ_reg_6_ ( .CK(newNet_63), .D(n_3112), .Q(pZ_6_) );
BUF_X2 newInst_849 ( .a(newNet_848), .o(newNet_849) );
INV_X1 g59555 ( .a(n_1570), .o(n_1571) );
NAND2_Z01 g34814 ( .a(n_3566), .b(GPR_18__2_), .o(n_3749) );
AND2_X1 g58261 ( .a(n_2752), .b(n_2209), .o(n_2806) );
BUF_X2 newInst_958 ( .a(newNet_957), .o(newNet_958) );
NAND2_Z01 g34885 ( .a(n_3630), .b(pX_11_), .o(n_3678) );
INV_X1 g59211 ( .a(n_1894), .o(n_1893) );
BUF_X2 newInst_185 ( .a(newNet_184), .o(newNet_185) );
BUF_X2 newInst_321 ( .a(newNet_320), .o(newNet_321) );
BUF_X2 newInst_994 ( .a(newNet_993), .o(newNet_994) );
INV_X1 g59419 ( .a(n_1697), .o(n_1698) );
NOR2_Z1 g35345 ( .a(n_4489), .b(n_3231), .o(n_4652) );
AND2_X1 g59427 ( .a(n_1667), .b(PC_7_), .o(n_1692) );
NAND2_Z01 g34761 ( .a(n_3582), .b(GPR_0__4_), .o(n_3804) );
AND2_X1 g60756 ( .a(n_175), .b(n_116), .o(n_387) );
INV_X1 g60528 ( .a(n_613), .o(n_614) );
NAND2_Z01 g59942 ( .a(n_1026), .b(n_458), .o(n_1183) );
XOR2_X1 g34460 ( .a(n_4057), .b(pY_10_), .o(n_4082) );
NAND2_Z01 g35266 ( .a(U_12_), .b(n_3275), .o(n_3407) );
AND2_X1 g61003 ( .a(n_4445), .b(n_4429), .o(n_136) );
BUF_X2 newInst_1391 ( .a(newNet_1390), .o(newNet_1391) );
BUF_X2 newInst_1007 ( .a(newNet_1006), .o(newNet_1007) );
NOR2_Z1 g35213 ( .a(n_3335), .b(n_3332), .o(n_3437) );
INV_Z1 g16796 ( .a(n_4465), .o(n_4419) );
BUF_X2 newInst_976 ( .a(newNet_975), .o(newNet_976) );
BUF_X2 newInst_1838 ( .a(newNet_20), .o(newNet_1838) );
INV_X1 g59908 ( .a(n_1221), .o(n_1222) );
AND2_X1 g59721 ( .a(n_1345), .b(n_1031), .o(n_1406) );
NAND2_Z01 g34168 ( .a(n_4318), .b(n_3351), .o(n_4342) );
BUF_X2 newInst_822 ( .a(newNet_821), .o(newNet_822) );
BUF_X2 newInst_1598 ( .a(newNet_1597), .o(newNet_1598) );
INV_X1 g35110 ( .a(n_3486), .o(n_3487) );
NAND2_Z01 g59168 ( .a(n_1895), .b(n_1870), .o(n_1978) );
BUF_X2 newInst_211 ( .a(newNet_210), .o(newNet_211) );
NOR4_Z1 g35097 ( .a(n_4491), .b(n_3430), .c(n_4634), .d(pmem_d_8), .o(n_4657) );
NOR2_Z1 g59425 ( .a(n_1668), .b(n_595), .o(n_1699) );
NAND2_Z01 g60927 ( .a(n_116), .b(state_3_), .o(n_218) );
NOR3_Z1 g58612 ( .a(n_4615), .b(n_2442), .c(pmem_d_8), .o(n_2486) );
NOR4_Z1 g58019 ( .a(n_2751), .b(n_2849), .c(n_2939), .d(n_2721), .o(n_2953) );
BUF_X2 newInst_948 ( .a(newNet_947), .o(newNet_948) );
NAND2_Z01 g59017 ( .a(n_2059), .b(pmem_d_4), .o(n_2113) );
XOR2_X1 g59498 ( .a(n_1574), .b(n_289), .o(n_1630) );
BUF_X2 newInst_217 ( .a(newNet_216), .o(newNet_217) );
NAND2_Z01 g58471 ( .a(n_2372), .b(n_2585), .o(n_2625) );
BUF_X2 newInst_1434 ( .a(newNet_1088), .o(newNet_1434) );
NAND2_Z01 g60314 ( .a(n_570), .b(pZ_2_), .o(n_812) );
fflopd GPR_reg_12__0_ ( .CK(newNet_1677), .D(n_2637), .Q(GPR_12__0_) );
BUF_X2 newInst_779 ( .a(newNet_778), .o(newNet_779) );
NAND2_Z01 g59877 ( .a(n_1025), .b(n_1170), .o(n_1250) );
fflopd state_reg_0_ ( .CK(newNet_27), .D(n_2722), .Q(state_0_) );
NAND2_Z01 g60297 ( .a(R16_9_), .b(n_571), .o(n_827) );
NAND2_Z01 g58445 ( .a(n_2622), .b(n_2198), .o(n_2648) );
NOR2_Z1 g34328 ( .a(n_4153), .b(n_4178), .o(n_4206) );
NAND2_Z01 g60289 ( .a(R16_1_), .b(n_571), .o(n_835) );
NAND2_Z01 g34782 ( .a(n_3587), .b(GPR_2__3_), .o(n_3783) );
fflopd GPR_reg_13__3_ ( .CK(newNet_1598), .D(n_2862), .Q(GPR_13__3_) );
NOR2_Z1 g35412 ( .a(n_3254), .b(n_3248), .o(n_4686) );
BUF_X2 newInst_1486 ( .a(newNet_1485), .o(newNet_1486) );
BUF_X2 newInst_1825 ( .a(newNet_1824), .o(newNet_1825) );
AND2_X1 g60823 ( .a(n_266), .b(n_173), .o(n_305) );
NAND3_Z1 g34550 ( .a(n_3847), .b(n_3849), .c(n_3848), .o(n_4009) );
fflopd U_reg_9_ ( .CK(newNet_361), .D(n_2866), .Q(U_9_) );
NAND2_Z01 g60444 ( .a(n_353), .b(GPR_10__1_), .o(n_702) );
NAND2_Z01 g34256 ( .a(n_4176), .b(pX_7_), .o(n_4277) );
BUF_X1 drc_bufs61131 ( .a(n_1875), .o(n_18) );
INV_X1 g60531 ( .a(n_606), .o(n_607) );
NAND2_Z02 g58920 ( .a(n_2154), .b(n_1204), .o(n_2202) );
NAND4_Z1 g57915 ( .a(n_1929), .b(n_2524), .c(n_2984), .d(n_2017), .o(n_3024) );
NOR2_Z1 g59984 ( .a(n_1035), .b(rst), .o(n_1144) );
NAND2_Z01 g60420 ( .a(n_347), .b(GPR_9__2_), .o(n_726) );
INV_X2 g61111 ( .a(rst), .o(n_41) );
NOR2_Z1 g35326 ( .a(n_3266), .b(n_3309), .o(n_3343) );
BUF_X2 newInst_827 ( .a(newNet_826), .o(newNet_827) );
fflopd GPR_reg_14__0_ ( .CK(newNet_1578), .D(n_2635), .Q(GPR_14__0_) );
BUF_X2 newInst_1845 ( .a(newNet_1295), .o(newNet_1845) );
NAND2_Z01 g34857 ( .a(n_3567), .b(GPR_6__0_), .o(n_3706) );
BUF_X2 newInst_1222 ( .a(newNet_1221), .o(newNet_1222) );
AND2_X1 g60832 ( .a(n_270), .b(n_144), .o(n_299) );
BUF_X2 newInst_399 ( .a(newNet_398), .o(newNet_399) );
NAND2_Z01 g57922 ( .a(n_2987), .b(n_2301), .o(n_3023) );
fflopd GPR_Rd_r_reg_2_ ( .CK(newNet_1861), .D(io_do_2), .Q(GPR_Rd_r_2_) );
INV_X1 g61069 ( .a(PC_6_), .o(n_83) );
AND2_X1 g35362 ( .a(n_3300), .b(n_3271), .o(n_3326) );
fflopd GPR_reg_14__5_ ( .CK(newNet_1543), .D(n_3017), .Q(GPR_14__5_) );
BUF_X2 newInst_1191 ( .a(newNet_1190), .o(newNet_1191) );
BUF_X2 newInst_1516 ( .a(newNet_1515), .o(newNet_1516) );
NAND2_Z01 g34869 ( .a(n_3582), .b(GPR_0__7_), .o(n_3694) );
NAND2_Z01 g34813 ( .a(n_3567), .b(GPR_6__2_), .o(n_3750) );
NOR3_Z1 g58655 ( .a(n_1911), .b(n_2280), .c(n_1260), .o(n_2447) );
BUF_X2 newInst_1611 ( .a(newNet_1610), .o(newNet_1611) );
NOR2_Z1 g59349 ( .a(n_1703), .b(n_1386), .o(n_1771) );
BUF_X2 newInst_748 ( .a(newNet_747), .o(newNet_748) );
NAND2_Z01 g60700 ( .a(GPR_7__6_), .b(n_183), .o(n_438) );
NAND2_Z01 g59391 ( .a(n_1648), .b(dmem_di_2), .o(n_1724) );
INV_X1 g60169 ( .a(n_968), .o(n_967) );
BUF_X2 newInst_1522 ( .a(newNet_1521), .o(newNet_1522) );
NAND2_Z01 g60071 ( .a(n_841), .b(io_do_6), .o(n_1063) );
BUF_X2 newInst_150 ( .a(newNet_149), .o(newNet_150) );
NAND2_Z01 g59397 ( .a(n_1648), .b(dmem_di_7), .o(n_1718) );
NOR2_Z1 g59789 ( .a(n_1269), .b(n_1161), .o(n_1335) );
NAND2_Z01 g58581 ( .a(n_2480), .b(pZ_13_), .o(n_2517) );
NOR2_Z1 g34719 ( .a(n_3624), .b(n_4410), .o(n_3846) );
NOR2_Z1 g34185 ( .a(n_4324), .b(n_4625), .o(n_4426) );
BUF_X2 newInst_287 ( .a(newNet_202), .o(newNet_287) );
NAND2_Z01 g34600 ( .a(n_3872), .b(n_3871), .o(n_3958) );
INV_Z1 g16803 ( .a(n_4656), .o(n_4412) );
XOR2_X1 g35147 ( .a(n_3450), .b(n_3236), .o(n_3471) );
NAND2_Z01 g59855 ( .a(n_563), .b(n_1170), .o(n_1274) );
NAND2_Z01 g34523 ( .a(n_3960), .b(pZ_6_), .o(n_4027) );
NAND2_Z01 g57883 ( .a(n_3010), .b(n_2198), .o(n_3055) );
NAND2_Z01 g60469 ( .a(n_353), .b(GPR_8__3_), .o(n_677) );
BUF_X2 newInst_149 ( .a(newNet_34), .o(newNet_149) );
AND2_X1 g59130 ( .a(n_1873), .b(pX_14_), .o(n_1985) );
NOR4_Z1 g34194 ( .a(n_4221), .b(n_4254), .c(n_4290), .d(n_4119), .o(n_4329) );
INV_X1 g61086 ( .a(n_4556), .o(n_66) );
BUF_X2 newInst_80 ( .a(newNet_79), .o(newNet_80) );
NAND2_Z01 g34618 ( .a(n_3894), .b(n_3489), .o(n_3942) );
NOR2_Z1 g59266 ( .a(n_1749), .b(n_1328), .o(n_1844) );
XOR2_X1 g34383 ( .a(n_4094), .b(pZ_12_), .o(n_4155) );
fflopd pX_reg_8_ ( .CK(newNet_201), .D(n_2725), .Q(pX_8_) );
NOR2_Z1 g34392 ( .a(n_4611), .b(n_3256), .o(n_4146) );
NAND2_Z01 g57934 ( .a(n_2973), .b(n_2408), .o(n_3008) );
NAND2_Z01 g58902 ( .a(n_2148), .b(n_1839), .o(n_2219) );
NAND2_Z01 g34686 ( .a(n_3597), .b(GPR_17__7_), .o(n_3879) );
INV_X1 g59677 ( .a(n_1446), .o(n_1447) );
NAND2_Z01 g34900 ( .a(n_3590), .b(pY_5_), .o(n_3663) );
AND2_X1 g59717 ( .a(n_1382), .b(PC_9_), .o(n_1409) );
BUF_X2 newInst_1563 ( .a(newNet_1562), .o(newNet_1563) );
NAND2_Z01 g58785 ( .a(n_2200), .b(GPR_7__4_), .o(n_2315) );
fflopd GPR_reg_10__6_ ( .CK(newNet_1723), .D(n_3090), .Q(GPR_10__6_) );
NAND2_Z01 g34190 ( .a(n_4325), .b(n_4466), .o(n_4333) );
NAND2_Z01 g58877 ( .a(n_2153), .b(GPR_8__3_), .o(n_2230) );
NAND2_Z01 g58149 ( .a(n_2816), .b(n_2238), .o(n_2864) );
BUF_X2 newInst_545 ( .a(newNet_544), .o(newNet_545) );
NOR2_Z1 g34420 ( .a(n_4088), .b(n_4028), .o(n_4117) );
BUF_X2 newInst_225 ( .a(newNet_224), .o(newNet_225) );
NAND2_Z01 g34543 ( .a(n_3921), .b(n_3908), .o(pmem_a_1) );
BUF_X2 newInst_1298 ( .a(newNet_1297), .o(newNet_1298) );
XNOR2_X1 g58832 ( .a(n_2162), .b(n_1831), .o(n_2275) );
NOR2_Z2 g34364 ( .a(n_3209), .b(n_4039), .o(n_4176) );
INV_X1 g59454 ( .a(n_1665), .o(n_1666) );
NAND2_Z02 g58911 ( .a(n_2161), .b(n_1202), .o(n_2211) );
NAND2_Z01 g35054 ( .a(n_3505), .b(n_3295), .o(n_3529) );
NAND2_Z01 g59570 ( .a(n_1470), .b(pmem_d_1), .o(n_1558) );
NAND4_Z1 g35014 ( .a(n_3351), .b(n_3464), .c(n_3497), .d(n_3447), .o(n_3558) );
NAND2_Z01 g59335 ( .a(n_1676), .b(SP_12_), .o(n_1779) );
NAND2_Z01 g58461 ( .a(n_2597), .b(n_2261), .o(n_2635) );
NAND2_Z01 g59050 ( .a(n_18), .b(n_4573), .o(n_2057) );
NAND2_Z01 g59151 ( .a(n_1896), .b(n_1122), .o(n_1948) );
AND2_X1 g60056 ( .a(n_845), .b(n_45), .o(n_1078) );
BUF_X2 newInst_886 ( .a(newNet_885), .o(newNet_886) );
NAND2_Z01 g58839 ( .a(n_2159), .b(GPR_10__5_), .o(n_2268) );
NAND2_Z01 g35436 ( .a(n_3243), .b(n_3236), .o(n_3273) );
NAND2_Z01 g60545 ( .a(n_21), .b(Rd_r_2_), .o(n_561) );
AND3_X1 g59195 ( .a(n_615), .b(n_1893), .c(pY_4_), .o(n_1914) );
NAND2_Z01 g34832 ( .a(n_3582), .b(GPR_0__1_), .o(n_3731) );
NOR2_Z2 g60995 ( .a(n_4649), .b(rst), .o(n_178) );
NOR2_Z1 g34642 ( .a(n_3642), .b(n_3435), .o(n_3918) );
NAND2_Z01 g34542 ( .a(n_3922), .b(n_3909), .o(pmem_a_2) );
INV_X2 newInst_1738 ( .a(newNet_19), .o(newNet_1738) );
fflopd GPR_reg_9__1_ ( .CK(newNet_683), .D(n_2735), .Q(GPR_9__1_) );
NOR3_Z1 g59663 ( .a(n_850), .b(n_1344), .c(io_do_2), .o(n_1464) );
XOR2_X1 g60394 ( .a(n_467), .b(pZ_3_), .o(n_752) );
INV_X1 g59128 ( .a(n_1968), .o(n_1969) );
NAND2_Z01 g58844 ( .a(n_2139), .b(GPR_11__4_), .o(n_2263) );
NAND2_Z01 g34864 ( .a(n_3628), .b(GPR_19__0_), .o(n_3699) );
BUF_X2 newInst_1060 ( .a(newNet_1059), .o(newNet_1060) );
AND2_X1 g34507 ( .a(n_4026), .b(n_3210), .o(n_4038) );
BUF_X2 newInst_28 ( .a(newNet_27), .o(newNet_28) );
NAND2_Z01 g60061 ( .a(n_843), .b(pmem_d_7), .o(n_1073) );
NAND2_Z01 g58311 ( .a(n_2682), .b(n_2379), .o(n_2759) );
NAND2_Z01 g60045 ( .a(n_765), .b(n_343), .o(n_1085) );
NAND2_Z01 g35286 ( .a(pZ_14_), .b(n_3199), .o(n_3389) );
BUF_X2 newInst_665 ( .a(newNet_664), .o(newNet_665) );
NAND2_Z01 g59120 ( .a(n_1893), .b(n_1901), .o(n_2058) );
NOR2_Z1 g34827 ( .a(n_3580), .b(n_4406), .o(n_3736) );
fflopd SP_reg_6_ ( .CK(newNet_482), .D(n_1742), .Q(SP_6_) );
NOR2_Z1 g59603 ( .a(n_1442), .b(n_4411), .o(n_1523) );
fflopd GPR_reg_1__4_ ( .CK(newNet_1233), .D(n_2935), .Q(GPR_1__4_) );
BUF_X2 newInst_1306 ( .a(newNet_1305), .o(newNet_1306) );
BUF_X2 newInst_1677 ( .a(newNet_1676), .o(newNet_1677) );
BUF_X2 newInst_282 ( .a(newNet_239), .o(newNet_282) );
BUF_X2 newInst_1812 ( .a(newNet_1811), .o(newNet_1812) );
XOR2_X1 g60865 ( .a(n_4448), .b(n_4432), .o(n_283) );
NAND2_Z01 g58036 ( .a(n_2909), .b(n_2269), .o(n_2949) );
AND2_X1 g57740 ( .a(n_3115), .b(n_2211), .o(n_3132) );
BUF_X2 newInst_1616 ( .a(newNet_1615), .o(newNet_1616) );
fflopd GPR_reg_23__5_ ( .CK(newNet_1037), .D(n_3004), .Q(GPR_23__5_) );
fflopd GPR_reg_9__4_ ( .CK(newNet_675), .D(n_2923), .Q(GPR_9__4_) );
INV_X1 g59912 ( .a(n_1200), .o(n_1201) );
NOR2_Z1 g34996 ( .a(n_3553), .b(n_3484), .o(n_3586) );
AND2_X1 g58520 ( .a(n_2567), .b(n_14), .o(n_2588) );
NAND2_Z01 g58304 ( .a(n_2693), .b(n_2411), .o(n_2766) );
AND3_X1 g59043 ( .a(n_4527), .b(n_1982), .c(pZ_12_), .o(n_2066) );
INV_X1 drc_bufs61182 ( .a(n_969), .o(n_26) );
NAND2_Z01 g59285 ( .a(n_1761), .b(n_1040), .o(n_1823) );
NAND4_Z1 g58942 ( .a(n_1500), .b(n_1908), .c(n_2100), .d(n_1499), .o(n_2165) );
XOR2_X1 final_adder_mux_R16_278_6_g412 ( .a(n_4449), .b(n_4433), .o(final_adder_mux_R16_278_6_n_37) );
NAND2_Z01 g60967 ( .a(n_39), .b(pmem_d_1), .o(n_153) );
BUF_X2 newInst_1394 ( .a(newNet_1393), .o(newNet_1394) );
BUF_X2 newInst_478 ( .a(newNet_477), .o(newNet_478) );
BUF_X2 newInst_1532 ( .a(newNet_1531), .o(newNet_1532) );
NAND2_Z01 g60486 ( .a(n_20), .b(Rd_r_2_), .o(n_660) );
NAND2_Z01 g58798 ( .a(n_2195), .b(U_11_), .o(n_2302) );
NAND2_Z01 g34809 ( .a(n_3599), .b(GPR_5__0_), .o(n_3754) );
BUF_X2 newInst_1581 ( .a(newNet_1580), .o(newNet_1581) );
NAND2_Z01 g58805 ( .a(n_2197), .b(U_3_), .o(n_2295) );
NAND2_Z01 g60512 ( .a(n_361), .b(GPR_5__0_), .o(n_634) );
INV_Z1 g35495 ( .a(pX_0_), .o(n_4574) );
BUF_X2 newInst_1192 ( .a(newNet_1191), .o(newNet_1192) );
BUF_X2 newInst_176 ( .a(newNet_33), .o(newNet_176) );
NAND2_Z01 g58170 ( .a(n_2796), .b(n_2230), .o(n_2840) );
BUF_X2 newInst_1137 ( .a(newNet_1136), .o(newNet_1137) );
NAND3_Z1 g59306 ( .a(n_849), .b(n_1694), .c(n_55), .o(n_1808) );
NAND3_Z1 g58486 ( .a(n_1796), .b(n_2575), .c(n_1096), .o(n_2610) );
NAND2_Z01 final_adder_mux_R16_278_6_g374 ( .a(final_adder_mux_R16_278_6_n_74), .b(final_adder_mux_R16_278_6_n_8), .o(final_adder_mux_R16_278_6_n_75) );
INV_X1 g35513 ( .a(pZ_7_), .o(n_3215) );
fflopd io_sp_reg_3_ ( .CK(newNet_322), .D(n_553), .Q(io_sp_3_) );
NOR2_Z2 g35045 ( .a(n_3526), .b(n_3467), .o(n_3536) );
BUF_X2 newInst_811 ( .a(newNet_810), .o(newNet_811) );
NAND2_Z01 g60322 ( .a(n_577), .b(pZ_14_), .o(n_805) );
INV_X1 g35474 ( .a(SP_7_), .o(n_3250) );
NAND4_Z1 g59252 ( .a(n_1722), .b(n_1683), .c(n_1791), .d(n_1089), .o(n_1860) );
NOR2_Z1 g35347 ( .a(n_3278), .b(pX_2_), .o(n_3356) );
AND2_X1 g60812 ( .a(n_277), .b(pmem_d_13), .o(n_310) );
NAND3_Z1 g59029 ( .a(n_1888), .b(n_2022), .c(n_1424), .o(n_2075) );
NAND4_Z1 g59206 ( .a(n_1278), .b(n_1240), .c(n_1814), .d(n_1746), .o(n_1905) );
AND2_X1 g35124 ( .a(n_3465), .b(n_3274), .o(n_3486) );
INV_X1 g34934 ( .a(n_3632), .o(n_3633) );
NOR2_Z1 g34476 ( .a(n_4647), .b(n_4646), .o(n_4068) );
BUF_X2 newInst_457 ( .a(newNet_456), .o(newNet_457) );
NAND2_Z01 g34638 ( .a(n_3769), .b(pZ_3_), .o(n_3922) );
NAND2_Z01 g58757 ( .a(n_2203), .b(GPR_4__1_), .o(n_2343) );
NOR2_Z1 g59979 ( .a(n_1047), .b(SP_6_), .o(n_1161) );
XOR2_X1 g60671 ( .a(n_171), .b(n_87), .o(n_478) );
NAND2_Z01 g34778 ( .a(n_3572), .b(GPR_4__3_), .o(n_3787) );
NOR2_Z1 g34425 ( .a(n_4088), .b(n_3557), .o(n_4112) );
fflopd GPR_reg_0__5_ ( .CK(newNet_1781), .D(n_2995), .Q(GPR_0__5_) );
BUF_X2 newInst_497 ( .a(newNet_496), .o(newNet_497) );
BUF_X2 newInst_18 ( .a(newNet_17), .o(newNet_18) );
NAND2_Z01 g59506 ( .a(n_1575), .b(n_148), .o(n_1614) );
NAND2_Z01 g60916 ( .a(PC_8_), .b(pmem_d_9), .o(n_262) );
INV_X2 newInst_1315 ( .a(newNet_1314), .o(newNet_1315) );
NAND2_Z01 g57823 ( .a(n_3053), .b(n_2267), .o(n_3090) );
BUF_X2 newInst_587 ( .a(newNet_586), .o(newNet_587) );
NAND2_Z01 g60233 ( .a(n_580), .b(GPR_14__0_), .o(n_912) );
NAND2_Z01 g59316 ( .a(n_1718), .b(n_1102), .o(n_1797) );
BUF_X2 newInst_1822 ( .a(newNet_1821), .o(newNet_1822) );
NAND2_Z01 g58953 ( .a(n_2092), .b(n_54), .o(n_2147) );
NAND2_Z01 g60560 ( .a(n_305), .b(n_273), .o(n_618) );
NAND4_Z1 g34122 ( .a(n_4274), .b(n_4302), .c(n_4312), .d(n_4138), .o(dmem_a_4) );
fflopd GPR_reg_12__4_ ( .CK(newNet_1640), .D(n_2947), .Q(GPR_12__4_) );
NAND2_Z01 g34766 ( .a(n_3591), .b(U_12_), .o(n_3799) );
fflopd PC_reg_5_ ( .CK(newNet_620), .D(n_2283), .Q(PC_5_) );
BUF_X2 newInst_1493 ( .a(newNet_1492), .o(newNet_1493) );
BUF_X2 newInst_297 ( .a(newNet_63), .o(newNet_297) );
INV_X1 g60951 ( .a(n_190), .o(n_191) );
NAND2_Z01 g60203 ( .a(n_575), .b(GPR_2__3_), .o(n_942) );
NOR2_Z1 g35340 ( .a(n_3240), .b(n_3309), .o(n_3331) );
BUF_X2 newInst_167 ( .a(newNet_136), .o(newNet_167) );
BUF_X2 newInst_1148 ( .a(newNet_1147), .o(newNet_1148) );
NAND2_Z01 g34107 ( .a(n_4340), .b(n_4354), .o(n_4446) );
BUF_X2 newInst_717 ( .a(newNet_716), .o(newNet_717) );
NOR2_Z1 g35353 ( .a(n_3311), .b(pmem_d_12), .o(n_3328) );
fflopd pY_reg_14_ ( .CK(newNet_171), .D(n_3141), .Q(pY_14_) );
AND2_X1 g59949 ( .a(n_837), .b(n_1031), .o(n_1179) );
NAND2_Z01 g59836 ( .a(n_1206), .b(io_do_6), .o(n_1289) );
NAND2_Z01 g34534 ( .a(n_3935), .b(n_3911), .o(pmem_a_4) );
NOR2_Z1 g59968 ( .a(n_1042), .b(n_205), .o(n_1170) );
NAND2_Z01 g58038 ( .a(n_2906), .b(n_2235), .o(n_2947) );
BUF_X2 newInst_611 ( .a(newNet_610), .o(newNet_611) );
BUF_X2 newInst_576 ( .a(newNet_429), .o(newNet_576) );
AND2_X1 g35294 ( .a(n_3263), .b(n_3298), .o(n_3381) );
BUF_X2 newInst_257 ( .a(newNet_30), .o(newNet_257) );
INV_X1 g34632 ( .a(n_3928), .o(n_4600) );
NAND2_Z01 g59293 ( .a(n_1772), .b(n_1803), .o(n_1830) );
NAND2_Z01 g34764 ( .a(n_3627), .b(GPR_15__4_), .o(n_3801) );
NAND4_Z1 g34572 ( .a(n_3825), .b(n_3828), .c(n_3827), .d(n_3826), .o(n_3988) );
NOR2_Z1 g35235 ( .a(n_3353), .b(pmem_d_3), .o(n_3433) );
NAND2_Z01 g60082 ( .a(n_589), .b(n_844), .o(n_1109) );
INV_X1 drc_bufs61122 ( .a(n_1701), .o(n_31) );
NAND2_Z02 g60360 ( .a(n_11), .b(n_45), .o(n_848) );
NAND2_Z01 g59628 ( .a(n_17), .b(T), .o(n_1499) );
INV_X1 g60090 ( .a(n_1039), .o(n_1038) );
BUF_X2 newInst_1023 ( .a(newNet_1022), .o(newNet_1023) );
NOR4_Z1 g58142 ( .a(n_2613), .b(n_2789), .c(n_2165), .d(n_1242), .o(n_2871) );
AND3_X1 g35091 ( .a(n_4662), .b(n_4661), .c(n_3318), .o(n_4629) );
NAND2_Z01 g60717 ( .a(n_200), .b(GPR_9__4_), .o(n_421) );
BUF_X2 newInst_1269 ( .a(newNet_1268), .o(newNet_1269) );
NAND2_Z01 g34610 ( .a(n_3691), .b(n_3690), .o(n_3950) );
NAND2_Z01 g60224 ( .a(n_578), .b(GPR_19__2_), .o(n_921) );
NAND3_Z1 g59181 ( .a(n_1752), .b(n_1846), .c(n_27), .o(n_1926) );
fflopd GPR_reg_4__2_ ( .CK(newNet_919), .D(n_2745), .Q(GPR_4__2_) );
NOR3_Z1 g59530 ( .a(n_1130), .b(n_1463), .c(n_885), .o(n_1597) );
INV_Z1 g16810 ( .a(GPR_15__3_), .o(n_4408) );
NAND4_Z1 g58138 ( .a(n_2069), .b(n_2548), .c(n_2830), .d(n_2020), .o(n_2875) );
NAND4_Z1 g59376 ( .a(n_770), .b(n_1475), .c(n_1660), .d(n_1363), .o(n_1742) );
AND2_X1 g58517 ( .a(n_2567), .b(n_2153), .o(n_2579) );
NAND2_Z01 g60496 ( .a(n_353), .b(GPR_8__6_), .o(n_650) );
BUF_X2 newInst_1216 ( .a(newNet_1215), .o(newNet_1216) );
AND2_X1 g59022 ( .a(n_1985), .b(n_1666), .o(n_2080) );
NOR4_Z1 g58651 ( .a(n_2106), .b(n_1458), .c(n_1249), .d(n_2130), .o(n_2450) );
BUF_X2 newInst_1607 ( .a(newNet_1606), .o(newNet_1607) );
NAND2_Z01 g34621 ( .a(n_3891), .b(n_3491), .o(n_3939) );
BUF_X2 newInst_101 ( .a(newNet_100), .o(newNet_101) );
XOR2_X1 g59736 ( .a(n_1225), .b(n_71), .o(n_1394) );
BUF_X2 newInst_106 ( .a(newNet_105), .o(newNet_106) );
NAND2_Z01 g34535 ( .a(n_3934), .b(n_3537), .o(n_4586) );
NAND2_Z01 g60558 ( .a(n_388), .b(n_399), .o(n_548) );
NAND2_Z01 g58159 ( .a(n_2806), .b(n_2401), .o(n_2854) );
NAND4_Z1 g57809 ( .a(n_1917), .b(n_2500), .c(n_3060), .d(n_2029), .o(n_3098) );
INV_X1 g35463 ( .a(pY_1_), .o(n_3261) );
NAND2_Z01 g58595 ( .a(n_2460), .b(pX_5_), .o(n_2500) );
AND2_X1 g57905 ( .a(n_3009), .b(n_2200), .o(n_3033) );
NAND4_Z1 g59547 ( .a(n_756), .b(n_1322), .c(n_1400), .d(n_14), .o(n_1581) );
NAND2_Z01 g58669 ( .a(n_2214), .b(GPR_16__4_), .o(n_2437) );
NAND4_Z1 g60005 ( .a(n_720), .b(n_829), .c(n_671), .d(n_557), .o(n_1124) );
AND2_X1 g58371 ( .a(n_2656), .b(n_2213), .o(n_2700) );
INV_X2 newInst_234 ( .a(newNet_233), .o(newNet_234) );
BUF_X2 newInst_522 ( .a(newNet_521), .o(newNet_522) );
BUF_X2 newInst_786 ( .a(newNet_385), .o(newNet_786) );
AND2_X1 g59712 ( .a(n_1325), .b(n_1311), .o(n_1420) );
NAND2_Z01 g59563 ( .a(n_1482), .b(n_1505), .o(n_1564) );
NAND2_Z01 g58681 ( .a(n_2212), .b(GPR_18__5_), .o(n_2425) );
NOR2_Z1 g35444 ( .a(pZ_1_), .b(pmem_d_1), .o(n_3271) );
BUF_X2 newInst_729 ( .a(newNet_728), .o(newNet_729) );
NAND2_Z01 g34140 ( .a(n_4317), .b(n_4619), .o(n_4368) );
NAND4_Z1 g58131 ( .a(n_1965), .b(n_2477), .c(n_2829), .d(n_2057), .o(n_2882) );
BUF_X2 newInst_188 ( .a(newNet_187), .o(newNet_188) );
NOR2_Z1 g60821 ( .a(n_177), .b(SP_4_), .o(n_306) );
NAND3_Z1 g34554 ( .a(n_3738), .b(n_3740), .c(n_3739), .o(n_4005) );
fflopd GPR_reg_20__2_ ( .CK(newNet_1200), .D(n_2764), .Q(GPR_20__2_) );
NAND2_Z01 g57687 ( .a(n_3157), .b(n_2194), .o(n_3179) );
BUF_X2 newInst_1631 ( .a(newNet_1630), .o(newNet_1631) );
NAND2_Z01 g58322 ( .a(n_2672), .b(n_2334), .o(n_2743) );
AND3_X1 g59190 ( .a(n_864), .b(n_1873), .c(pX_5_), .o(n_1917) );
NAND2_Z01 g35306 ( .a(n_3289), .b(pY_4_), .o(n_3370) );
NAND2_Z03 g34167 ( .a(n_4313), .b(n_3957), .o(io_do_3) );
BUF_X2 newInst_107 ( .a(newNet_106), .o(newNet_107) );
NOR2_Z1 g34965 ( .a(n_3547), .b(pX_9_), .o(n_3634) );
NOR2_Z1 g59390 ( .a(n_28), .b(n_60), .o(n_1725) );
NOR2_Z1 g59006 ( .a(n_1970), .b(n_105), .o(n_2102) );
BUF_X2 newInst_1373 ( .a(newNet_1372), .o(newNet_1373) );
BUF_X2 newInst_368 ( .a(newNet_367), .o(newNet_368) );
INV_X1 g35481 ( .a(pZ_2_), .o(n_3243) );
BUF_X2 newInst_139 ( .a(newNet_138), .o(newNet_139) );
NAND4_Z1 g59990 ( .a(n_816), .b(n_832), .c(n_802), .d(n_870), .o(n_1139) );
NAND4_Z1 g34248 ( .a(n_3666), .b(n_3704), .c(n_4173), .d(n_3703), .o(n_4285) );
BUF_X2 newInst_1071 ( .a(newNet_1070), .o(newNet_1071) );
NAND2_Z01 g58813 ( .a(n_2199), .b(GPR_0__7_), .o(n_2287) );
NAND2_Z01 g34104 ( .a(n_4341), .b(n_4357), .o(n_4445) );
NAND4_Z1 g34587 ( .a(n_3673), .b(n_3745), .c(n_3746), .d(n_3744), .o(n_3973) );
BUF_X2 newInst_636 ( .a(newNet_635), .o(newNet_636) );
INV_Y1 g35385 ( .a(n_3310), .o(n_4529) );
BUF_X2 newInst_1361 ( .a(newNet_1360), .o(newNet_1361) );
AND2_X1 g58106 ( .a(n_2850), .b(n_2158), .o(n_2906) );
NAND2_Z01 g58537 ( .a(n_2530), .b(pZ_15_), .o(n_2560) );
NAND2_Z01 g59465 ( .a(n_1628), .b(n_83), .o(n_1667) );
AND2_X1 g58369 ( .a(n_2657), .b(n_2156), .o(n_2702) );
INV_X1 g61107 ( .a(pmem_d_12), .o(n_45) );
NAND2_Z01 g58478 ( .a(n_2579), .b(n_2233), .o(n_2616) );
NAND2_Z02 g58966 ( .a(n_2088), .b(n_1213), .o(n_2153) );
NOR2_Z1 g34347 ( .a(n_4178), .b(n_4061), .o(n_4187) );
NAND2_Z01 g34131 ( .a(n_4164), .b(GPR_Rd_r_4_), .o(n_4377) );
BUF_X2 newInst_812 ( .a(newNet_811), .o(newNet_812) );
NAND2_Z01 g34115 ( .a(n_4332), .b(n_4346), .o(n_4433) );
NAND2_Z01 g59744 ( .a(n_1315), .b(n_141), .o(n_1378) );
INV_X2 newInst_1221 ( .a(newNet_1220), .o(newNet_1221) );
fflopd GPR_reg_14__2_ ( .CK(newNet_1564), .D(n_2778), .Q(GPR_14__2_) );
NAND2_Z01 g57946 ( .a(n_2961), .b(n_2191), .o(n_2996) );
BUF_X2 newInst_1687 ( .a(newNet_1686), .o(newNet_1687) );
AND2_X1 g58120 ( .a(n_2850), .b(n_2205), .o(n_2892) );
AND2_X1 g58646 ( .a(n_2354), .b(n_1931), .o(n_2461) );
BUF_X2 newInst_1285 ( .a(newNet_1284), .o(newNet_1285) );
NAND2_Z01 g58679 ( .a(n_2212), .b(GPR_18__3_), .o(n_2427) );
NAND2_Z01 g60220 ( .a(n_575), .b(GPR_2__6_), .o(n_925) );
BUF_X2 newInst_671 ( .a(newNet_663), .o(newNet_671) );
NAND2_Z01 g59621 ( .a(n_1415), .b(S), .o(n_1506) );
NOR2_Z1 g60604 ( .a(n_462), .b(n_199), .o(n_598) );
BUF_X2 newInst_1857 ( .a(newNet_1052), .o(newNet_1857) );
NAND2_Z01 g59752 ( .a(n_1312), .b(io_do_1), .o(n_1372) );
AND2_X1 g59584 ( .a(n_1269), .b(n_1484), .o(n_1544) );
BUF_X2 newInst_379 ( .a(newNet_378), .o(newNet_379) );
fflopd GPR_reg_19__5_ ( .CK(newNet_1285), .D(n_3012), .Q(GPR_19__5_) );
XNOR2_X1 g35076 ( .a(n_3493), .b(PC_6_), .o(n_4543) );
NAND2_Z02 g59244 ( .a(n_1828), .b(n_291), .o(n_1873) );
NAND4_Z1 g60380 ( .a(n_396), .b(n_411), .c(n_452), .d(n_456), .o(n_765) );
BUF_X2 newInst_1365 ( .a(newNet_1364), .o(newNet_1365) );
AND3_X1 g59035 ( .a(n_47), .b(n_1867), .c(pmem_d_5), .o(n_2083) );
NOR2_Z1 g34454 ( .a(n_4075), .b(n_4645), .o(n_4087) );
BUF_X2 newInst_198 ( .a(newNet_197), .o(newNet_198) );
NAND2_Z01 g60411 ( .a(n_347), .b(GPR_9__6_), .o(n_735) );
NOR2_Z1 g59972 ( .a(n_1042), .b(n_172), .o(n_1164) );
NAND2_Z01 g59509 ( .a(n_1573), .b(SP_4_), .o(n_1612) );
AND2_X1 g58404 ( .a(n_2656), .b(n_2140), .o(n_2664) );
AND2_X1 g59525 ( .a(n_1269), .b(n_1569), .o(n_1604) );
NAND2_Z01 g58643 ( .a(n_2357), .b(n_2004), .o(n_2463) );
XOR2_X1 g35200 ( .a(n_3322), .b(n_3300), .o(n_3454) );
NAND2_Z01 g35404 ( .a(pZ_7_), .b(pZ_6_), .o(n_4525) );
BUF_X2 newInst_1708 ( .a(newNet_1707), .o(newNet_1708) );
BUF_X2 newInst_1244 ( .a(newNet_1243), .o(newNet_1244) );
NAND2_Z01 g34467 ( .a(n_4647), .b(n_4646), .o(n_4075) );
INV_Z1 g16812 ( .a(GPR_8__4_), .o(n_4405) );
NOR2_Z1 g59503 ( .a(n_1566), .b(n_817), .o(n_1617) );
NAND2_Z01 g59276 ( .a(n_1801), .b(n_1654), .o(n_1851) );
NAND2_Z01 g34682 ( .a(n_3628), .b(GPR_19__7_), .o(n_3883) );
BUF_X2 newInst_1103 ( .a(newNet_366), .o(newNet_1103) );
NAND2_Z01 g60729 ( .a(n_196), .b(n_4484), .o(n_410) );
NAND2_Z01 g59221 ( .a(n_1853), .b(n_1707), .o(n_1885) );
AND2_X1 g58000 ( .a(n_2940), .b(n_2208), .o(n_2971) );
XOR2_X1 final_adder_mux_R16_278_6_g367 ( .a(final_adder_mux_R16_278_6_n_80), .b(final_adder_mux_R16_278_6_n_32), .o(R16_13_) );
XOR2_X1 g60855 ( .a(n_4436), .b(n_4420), .o(n_332) );
BUF_X2 newInst_1014 ( .a(newNet_1013), .o(newNet_1014) );
BUF_X2 newInst_430 ( .a(newNet_429), .o(newNet_430) );
BUF_X2 newInst_1056 ( .a(newNet_1055), .o(newNet_1056) );
NAND4_Z2 g35184 ( .a(n_3333), .b(n_3372), .c(n_3336), .d(n_3387), .o(n_4626) );
NAND2_Z01 g58890 ( .a(n_2140), .b(GPR_9__4_), .o(n_2192) );
BUF_X2 newInst_1468 ( .a(newNet_1467), .o(newNet_1468) );
NOR2_Z1 g34888 ( .a(n_3565), .b(n_3260), .o(n_3675) );
fflopd GPR_reg_6__0_ ( .CK(newNet_833), .D(n_2619), .Q(GPR_6__0_) );
AND3_X1 g34512 ( .a(n_4529), .b(n_3905), .c(state_2_), .o(n_4033) );
INV_X1 g59600 ( .a(n_1527), .o(n_1528) );
INV_X1 g34369 ( .a(n_4164), .o(n_4163) );
XOR2_X1 g34353 ( .a(n_4126), .b(SP_7_), .o(n_4182) );
BUF_X2 newInst_334 ( .a(newNet_333), .o(newNet_334) );
NOR2_Z1 g59170 ( .a(n_1895), .b(n_1205), .o(n_1935) );
AND2_X1 g58510 ( .a(n_2567), .b(n_2206), .o(n_2586) );
INV_X1 g34977 ( .a(n_3580), .o(n_3579) );
fflopd pX_reg_10_ ( .CK(newNet_281), .D(n_2870), .Q(pX_10_) );
BUF_X2 newInst_1114 ( .a(newNet_963), .o(newNet_1114) );
NAND2_Z01 g59931 ( .a(n_1119), .b(n_969), .o(n_1214) );
NAND2_Z01 g34164 ( .a(n_4317), .b(pmem_d_0), .o(n_4344) );
AND2_X1 g35222 ( .a(n_4683), .b(n_3220), .o(n_3434) );
BUF_X2 newInst_595 ( .a(newNet_594), .o(newNet_595) );
INV_X1 g61038 ( .a(pX_11_), .o(n_114) );
NAND3_Z1 g59649 ( .a(n_748), .b(n_1356), .c(n_387), .o(n_1489) );
NAND2_Z01 g58779 ( .a(n_2201), .b(GPR_6__7_), .o(n_2321) );
NAND2_Z01 g60888 ( .a(n_4685), .b(n_32), .o(n_239) );
BUF_X2 newInst_900 ( .a(newNet_594), .o(newNet_900) );
NAND2_Z01 g60227 ( .a(n_575), .b(GPR_2__2_), .o(n_918) );
BUF_X2 newInst_1721 ( .a(newNet_1720), .o(newNet_1721) );
NAND2_Z01 g60260 ( .a(n_590), .b(GPR_6__6_), .o(n_886) );
BUF_X2 newInst_907 ( .a(newNet_906), .o(newNet_907) );
XOR2_X1 g35017 ( .a(n_4515), .b(pX_8_), .o(n_4566) );
NOR2_Z1 g34273 ( .a(n_4613), .b(n_3261), .o(n_4260) );
NAND4_Z1 g57761 ( .a(n_1962), .b(n_2501), .c(n_3104), .d(n_2054), .o(n_3114) );
NAND4_Z1 g59997 ( .a(n_814), .b(n_880), .c(n_819), .d(n_900), .o(n_1132) );
NAND2_Z01 g59464 ( .a(n_10), .b(n_1602), .o(n_1668) );
XOR2_X1 g59366 ( .a(io_do_4), .b(n_1649), .o(n_1770) );
NAND2_Z01 g34739 ( .a(n_3597), .b(GPR_17__5_), .o(n_3826) );
BUF_X2 newInst_774 ( .a(newNet_773), .o(newNet_774) );
NOR2_Z1 g34321 ( .a(n_4612), .b(n_3498), .o(n_4212) );
BUF_X2 newInst_794 ( .a(newNet_793), .o(newNet_794) );
NAND2_Z01 g59587 ( .a(n_1488), .b(n_382), .o(n_1541) );
AND2_X1 g57999 ( .a(n_2940), .b(n_2209), .o(n_2972) );
NAND4_Z2 g35194 ( .a(n_3363), .b(n_3379), .c(n_3368), .d(n_3399), .o(n_4624) );
NAND2_Z02 g34455 ( .a(n_4071), .b(n_3930), .o(n_4088) );
BUF_X2 newInst_1863 ( .a(newNet_1270), .o(newNet_1863) );
NAND2_Z01 g60271 ( .a(n_590), .b(GPR_6__3_), .o(n_875) );
BUF_X2 newInst_1461 ( .a(newNet_1460), .o(newNet_1461) );
BUF_X2 newInst_1338 ( .a(newNet_1337), .o(newNet_1338) );
BUF_X2 newInst_863 ( .a(newNet_620), .o(newNet_863) );
BUF_X2 newInst_1663 ( .a(newNet_1662), .o(newNet_1663) );
NOR2_Z1 g59929 ( .a(n_1111), .b(n_123), .o(n_1217) );
AND2_X1 g58361 ( .a(n_2657), .b(n_2158), .o(n_2710) );
BUF_X2 newInst_138 ( .a(newNet_130), .o(newNet_138) );
NAND2_Z01 g60370 ( .a(n_485), .b(state_1_), .o(n_844) );
BUF_X2 newInst_468 ( .a(newNet_467), .o(newNet_468) );
AND3_X1 g59897 ( .a(n_4559), .b(n_999), .c(rst), .o(n_1232) );
NAND2_Z01 g34675 ( .a(n_3636), .b(GPR_10__7_), .o(n_3890) );
BUF_X2 newInst_1660 ( .a(newNet_1659), .o(newNet_1660) );
NOR2_Z1 g34171 ( .a(n_4324), .b(n_4682), .o(n_4429) );
BUF_X2 newInst_802 ( .a(newNet_801), .o(newNet_802) );
BUF_X2 newInst_637 ( .a(newNet_636), .o(newNet_637) );
NAND2_Z01 g59743 ( .a(n_1224), .b(io_sel_0_), .o(n_1379) );
fflopd GPR_reg_13__4_ ( .CK(newNet_5), .D(n_2946), .Q(GPR_13__4_) );
BUF_X2 newInst_1432 ( .a(newNet_1431), .o(newNet_1432) );
NOR2_Z1 g60791 ( .a(n_199), .b(n_202), .o(n_374) );
INV_X1 g35503 ( .a(pX_10_), .o(n_3224) );
BUF_X2 newInst_365 ( .a(newNet_364), .o(newNet_365) );
BUF_X2 newInst_245 ( .a(newNet_244), .o(newNet_245) );
NAND2_Z01 g59063 ( .a(n_1902), .b(n_4594), .o(n_2044) );
fflopd U_reg_3_ ( .CK(newNet_382), .D(n_2950), .Q(U_3_) );
XOR2_X1 final_adder_mux_R16_278_6_g394 ( .a(final_adder_mux_R16_278_6_n_53), .b(final_adder_mux_R16_278_6_n_39), .o(R16_4_) );
INV_X1 g61095 ( .a(n_4624), .o(n_57) );
AND2_X1 g60342 ( .a(n_589), .b(n_59), .o(n_788) );
XNOR2_X1 g59307 ( .a(n_1736), .b(pmem_d_10), .o(n_1825) );
BUF_X2 newInst_356 ( .a(newNet_355), .o(newNet_356) );
NOR2_Z1 g59954 ( .a(n_989), .b(n_1019), .o(n_1177) );
BUF_X2 newInst_855 ( .a(newNet_854), .o(newNet_855) );
BUF_X2 newInst_1205 ( .a(newNet_1204), .o(newNet_1205) );
fflopd U_reg_11_ ( .CK(newNet_430), .D(n_2951), .Q(U_11_) );
NAND2_Z01 g59630 ( .a(n_1421), .b(n_407), .o(n_1527) );
NOR2_Z1 g34175 ( .a(n_4324), .b(n_4623), .o(n_4425) );
NAND2_Z01 g58851 ( .a(n_2139), .b(GPR_11__5_), .o(n_2256) );
NAND2_Z01 g34720 ( .a(n_3586), .b(GPR_9__0_), .o(n_3845) );
NAND2_Z01 g60703 ( .a(GPR_1__4_), .b(n_183), .o(n_435) );
BUF_X2 newInst_1756 ( .a(newNet_1755), .o(newNet_1756) );
BUF_X2 newInst_1544 ( .a(newNet_985), .o(newNet_1544) );
BUF_X2 newInst_1344 ( .a(newNet_1343), .o(newNet_1344) );
AND2_X1 g57755 ( .a(n_3115), .b(n_2199), .o(n_3117) );
NAND2_Z01 g57719 ( .a(n_3121), .b(n_2321), .o(n_3148) );
BUF_X2 newInst_952 ( .a(newNet_951), .o(newNet_952) );
AND2_X1 g58259 ( .a(n_2752), .b(n_2211), .o(n_2808) );
AND2_X1 g60627 ( .a(n_460), .b(n_197), .o(n_583) );
NAND2_Z01 g58854 ( .a(n_2157), .b(GPR_13__1_), .o(n_2253) );
BUF_X2 newInst_159 ( .a(newNet_137), .o(newNet_159) );
NAND2_Z01 g60893 ( .a(SP_0_), .b(SP_1_), .o(n_275) );
NAND4_Z1 g59564 ( .a(n_568), .b(n_1383), .c(n_1357), .d(n_4660), .o(n_1563) );
INV_X2 newInst_1832 ( .a(newNet_1831), .o(newNet_1832) );
XOR2_X1 g34236 ( .a(n_4280), .b(SP_9_), .o(n_4295) );
AND2_X1 g57729 ( .a(n_3115), .b(n_2159), .o(n_3143) );
BUF_X2 newInst_1326 ( .a(newNet_225), .o(newNet_1326) );
NAND2_Z01 g60960 ( .a(n_63), .b(pmem_d_2), .o(n_157) );
NAND2_Z01 g58802 ( .a(n_2195), .b(U_15_), .o(n_2298) );
AND2_X1 g58270 ( .a(n_2752), .b(n_2200), .o(n_2797) );
NAND2_Z02 g35156 ( .a(n_3198), .b(pmem_d_4), .o(n_3469) );
BUF_X2 newInst_58 ( .a(newNet_57), .o(newNet_58) );
BUF_X2 newInst_43 ( .a(newNet_42), .o(newNet_43) );
AND2_X1 g59228 ( .a(n_1854), .b(io_do_7), .o(n_1892) );
INV_X1 g60771 ( .a(n_366), .o(n_367) );
BUF_X2 newInst_1159 ( .a(newNet_1158), .o(newNet_1159) );
BUF_X2 newInst_622 ( .a(newNet_621), .o(newNet_622) );
NAND2_Z01 g35450 ( .a(n_3214), .b(n_3248), .o(n_3281) );
NAND2_Z01 g60452 ( .a(n_368), .b(GPR_13__3_), .o(n_694) );
BUF_X2 newInst_662 ( .a(newNet_661), .o(newNet_662) );
NAND2_Z01 g58633 ( .a(n_2354), .b(pX_7_), .o(n_2469) );
XOR2_X1 g34517 ( .a(n_3959), .b(n_3223), .o(n_4028) );
NAND2_Z01 g35269 ( .a(U_6_), .b(n_3275), .o(n_3405) );
XOR2_X1 g60008 ( .a(n_866), .b(pZ_5_), .o(n_1122) );
BUF_X2 newInst_1015 ( .a(newNet_1014), .o(newNet_1015) );
BUF_X2 newInst_858 ( .a(newNet_857), .o(newNet_858) );
NAND2_Z01 g34679 ( .a(n_3630), .b(pX_15_), .o(n_3886) );
NAND4_Z1 g60099 ( .a(n_416), .b(n_424), .c(n_449), .d(n_448), .o(n_1020) );
AND3_X1 g59535 ( .a(n_339), .b(n_1551), .c(n_4488), .o(n_1592) );
NOR2_Z1 g58825 ( .a(n_2194), .b(n_1975), .o(n_2354) );
INV_X1 g61091 ( .a(io_do_6), .o(n_61) );
NAND2_Z01 g60406 ( .a(n_457), .b(GPR_16__5_), .o(n_740) );
BUF_X2 newInst_1531 ( .a(newNet_1530), .o(newNet_1531) );
BUF_X2 newInst_296 ( .a(newNet_295), .o(newNet_296) );
AND2_X1 g60349 ( .a(n_177), .b(n_567), .o(n_782) );
NAND2_Z01 g35441 ( .a(n_3256), .b(n_3220), .o(n_3284) );
BUF_X2 newInst_1234 ( .a(newNet_43), .o(newNet_1234) );
INV_X2 g59235 ( .a(n_1873), .o(n_1872) );
AND2_X1 g57990 ( .a(n_2940), .b(n_2158), .o(n_2981) );
BUF_X2 newInst_1797 ( .a(newNet_1796), .o(newNet_1797) );
XOR2_X1 g59737 ( .a(n_1314), .b(n_304), .o(n_1393) );
fflopd io_sp_reg_5_ ( .CK(newNet_308), .D(n_551), .Q(io_sp_5_) );
BUF_X2 newInst_466 ( .a(newNet_114), .o(newNet_466) );
INV_X1 g61084 ( .a(io_do_3), .o(n_68) );
AND2_X1 g59370 ( .a(n_1735), .b(n_853), .o(n_1745) );
fflopd GPR_Rd_r_reg_4_ ( .CK(newNet_1849), .D(io_do_4), .Q(GPR_Rd_r_4_) );
XOR2_X1 g35100 ( .a(n_3466), .b(pZ_5_), .o(n_3499) );
NAND2_Z01 g34644 ( .a(n_4538), .b(n_3768), .o(n_3916) );
NAND3_Z1 g59240 ( .a(n_803), .b(n_1813), .c(n_825), .o(n_1878) );
NOR2_Z1 g59435 ( .a(n_1646), .b(n_1456), .o(n_1684) );
NAND2_Z01 g60887 ( .a(n_42), .b(pmem_d_14), .o(n_277) );
NAND2_Z01 g34879 ( .a(n_3566), .b(GPR_18__7_), .o(n_3684) );
BUF_X2 newInst_1578 ( .a(newNet_1577), .o(newNet_1578) );
NOR2_Z1 g34289 ( .a(n_4163), .b(n_3233), .o(n_4244) );
XNOR2_X1 g34660 ( .a(n_3617), .b(PC_10_), .o(n_4537) );
BUF_X2 newInst_1454 ( .a(newNet_1453), .o(newNet_1454) );
NAND2_Z01 g58789 ( .a(n_2213), .b(GPR_17__2_), .o(n_2311) );
NAND2_Z01 g35300 ( .a(n_3299), .b(pX_9_), .o(n_3375) );
NOR2_Z1 g59083 ( .a(n_1883), .b(n_1848), .o(n_2024) );
BUF_X2 newInst_1449 ( .a(newNet_1448), .o(newNet_1449) );
BUF_X2 newInst_1120 ( .a(newNet_1119), .o(newNet_1120) );
INV_X1 g61063 ( .a(pZ_14_), .o(n_89) );
BUF_X2 newInst_313 ( .a(newNet_312), .o(newNet_313) );
BUF_X2 newInst_1253 ( .a(newNet_786), .o(newNet_1253) );
NAND2_Z01 g60561 ( .a(n_341), .b(pY_7_), .o(n_546) );
NAND2_Z01 g59481 ( .a(n_1602), .b(n_351), .o(n_1644) );
NAND2_Z01 g34149 ( .a(n_4325), .b(n_4682), .o(n_4359) );
fflopd GPR_reg_6__3_ ( .CK(newNet_814), .D(n_2842), .Q(GPR_6__3_) );
NAND2_Z01 g57822 ( .a(n_3055), .b(n_2293), .o(n_3091) );
NAND2_Z01 g35132 ( .a(n_3463), .b(n_3228), .o(n_3485) );
NOR2_Z4 g58530 ( .a(n_2557), .b(n_1590), .o(n_2567) );
BUF_X2 newInst_1320 ( .a(newNet_1319), .o(newNet_1320) );
BUF_X2 newInst_1020 ( .a(newNet_380), .o(newNet_1020) );
BUF_X2 newInst_764 ( .a(newNet_763), .o(newNet_764) );
AND2_X1 g34165 ( .a(n_3195), .b(n_4178), .o(n_4343) );
NAND2_Z01 g34699 ( .a(n_3587), .b(GPR_2__6_), .o(n_3866) );
NOR2_Z1 g60633 ( .a(n_338), .b(n_205), .o(n_501) );
NAND2_Z01 g59818 ( .a(n_1193), .b(n_232), .o(n_1314) );
BUF_X2 newInst_1400 ( .a(newNet_1399), .o(newNet_1400) );
NAND2_Z01 g34781 ( .a(n_3568), .b(GPR_22__3_), .o(n_3784) );
BUF_X2 newInst_1084 ( .a(newNet_1083), .o(newNet_1084) );
NAND2_Z01 g60264 ( .a(n_590), .b(GPR_6__0_), .o(n_882) );
INV_X1 g61031 ( .a(PC_8_), .o(n_121) );
NAND2_Z01 g60901 ( .a(PC_2_), .b(pmem_d_5), .o(n_269) );
NAND2_Z01 g60242 ( .a(n_574), .b(GPR_10__2_), .o(n_903) );
NAND2_Z01 g58286 ( .a(n_2712), .b(n_2187), .o(n_2784) );
NAND2_Z01 g60436 ( .a(n_349), .b(U_3_), .o(n_710) );
AND2_X1 g34490 ( .a(n_4033), .b(state_3_), .o(n_4647) );
NAND2_Z01 g34695 ( .a(n_3636), .b(GPR_10__6_), .o(n_3870) );
BUF_X2 newInst_517 ( .a(newNet_516), .o(newNet_517) );
AND2_X1 g60057 ( .a(n_844), .b(n_48), .o(n_1077) );
BUF_X2 newInst_1377 ( .a(newNet_1376), .o(newNet_1377) );
NAND2_Z01 g34604 ( .a(n_3751), .b(n_3293), .o(n_3959) );
NOR4_Z1 g34245 ( .a(n_3667), .b(n_4031), .c(n_4167), .d(n_4017), .o(n_4288) );
NAND2_Z01 g34897 ( .a(n_3564), .b(pX_0_), .o(n_3666) );
INV_X1 g61112 ( .a(io_do_0), .o(n_40) );
fflopd GPR_reg_22__5_ ( .CK(newNet_1076), .D(n_3005), .Q(GPR_22__5_) );
BUF_X1 mybuffer5 ( .o(io_a_5), .a(pmem_d_10) );
NAND2_Z02 g58922 ( .a(n_2154), .b(n_1202), .o(n_2200) );
NOR4_Z1 g58278 ( .a(n_2570), .b(n_2658), .c(n_2446), .d(n_1247), .o(n_2790) );
NOR2_Z1 g60587 ( .a(n_363), .b(pZ_13_), .o(n_610) );
NAND2_Z01 g59416 ( .a(n_39), .b(n_1664), .o(n_1729) );
fflopd GPR_reg_16__1_ ( .CK(newNet_1473), .D(n_2774), .Q(GPR_16__1_) );
NOR2_Z1 g60828 ( .a(n_199), .b(n_248), .o(n_347) );
NAND3_Z1 g58338 ( .a(n_2472), .b(n_2650), .c(n_2112), .o(n_2731) );
NAND4_Z1 g34123 ( .a(n_4271), .b(n_4298), .c(n_4311), .d(n_4136), .o(dmem_a_2) );
AND2_X1 final_adder_mux_R16_278_6_g437 ( .a(n_4441), .b(n_4425), .o(final_adder_mux_R16_278_6_n_12) );
BUF_X2 newInst_1509 ( .a(newNet_1508), .o(newNet_1509) );
fflopd GPR_reg_21__5_ ( .CK(newNet_1125), .D(n_3006), .Q(GPR_21__5_) );
BUF_X2 newInst_809 ( .a(newNet_808), .o(newNet_809) );
fflopd pZ_reg_12_ ( .CK(newNet_99), .D(n_3026), .Q(pZ_12_) );
NAND2_Z01 g59969 ( .a(n_1026), .b(n_165), .o(n_1152) );
NAND2_Z01 g59791 ( .a(n_1266), .b(n_1170), .o(n_1333) );
NOR2_Z1 g34305 ( .a(n_16064_BAR), .b(n_3765), .o(n_4228) );
NAND2_Z01 g59620 ( .a(n_1413), .b(io_sp_4_), .o(n_1507) );
NAND2_Z01 g35028 ( .a(n_3526), .b(n_3467), .o(n_3553) );
AND3_X1 g35374 ( .a(pY_9_), .b(pY_8_), .c(pY_11_), .o(n_3316) );
BUF_X2 newInst_915 ( .a(newNet_914), .o(newNet_915) );
NAND2_Z01 g58474 ( .a(n_2336), .b(n_2582), .o(n_2620) );
NAND2_Z01 g58680 ( .a(n_2212), .b(GPR_18__4_), .o(n_2426) );
NAND2_Z01 g58047 ( .a(n_2898), .b(n_2409), .o(n_2935) );
BUF_X2 newInst_648 ( .a(newNet_647), .o(newNet_648) );
NAND2_Z01 g34136 ( .a(n_4317), .b(n_4644), .o(n_4372) );
NOR4_Z1 g60662 ( .a(n_59), .b(n_4684), .c(n_4478), .d(pmem_d_12), .o(n_484) );
NAND2_Z01 g34755 ( .a(n_3568), .b(GPR_22__4_), .o(n_3810) );
BUF_X2 newInst_1817 ( .a(newNet_264), .o(newNet_1817) );
NAND2_Z01 g58148 ( .a(n_2817), .b(n_2270), .o(n_2865) );
fflopd GPR_reg_4__3_ ( .CK(newNet_916), .D(n_2844), .Q(GPR_4__3_) );
BUF_X2 newInst_1447 ( .a(newNet_1446), .o(newNet_1447) );
NAND2_Z01 g58871 ( .a(n_2155), .b(GPR_14__1_), .o(n_2236) );
BUF_X2 newInst_722 ( .a(newNet_721), .o(newNet_722) );
NOR2_Z1 g59341 ( .a(n_1708), .b(n_37), .o(n_1776) );
NAND2_Z01 g58678 ( .a(n_2212), .b(GPR_18__2_), .o(n_2428) );
AND2_X1 g59567 ( .a(n_1487), .b(n_93), .o(n_1561) );
NOR2_Z2 g59226 ( .a(n_1829), .b(n_4611), .o(n_1896) );
NOR2_Z1 g34340 ( .a(n_4159), .b(n_3515), .o(n_4194) );
NAND2_Z01 g60751 ( .a(SP_13_), .b(n_180), .o(n_391) );
NAND2_Z01 g34143 ( .a(n_4325), .b(n_4625), .o(n_4365) );
NAND2_Z01 g57691 ( .a(n_3158), .b(n_2193), .o(n_3175) );
fflopd pX_reg_3_ ( .CK(newNet_234), .D(n_2958), .Q(pX_3_) );
AND2_X1 g60934 ( .a(n_4683), .b(n_32), .o(n_214) );
NAND2_Z01 g60216 ( .a(R16_10_), .b(n_14), .o(n_929) );
NAND2_Z01 g58594 ( .a(n_2460), .b(pX_6_), .o(n_2501) );
fflopd GPR_reg_7__3_ ( .CK(newNet_770), .D(n_2841), .Q(GPR_7__3_) );
INV_X1 g61104 ( .a(pmem_d_5), .o(n_48) );
NAND2_Z01 g59697 ( .a(io_do_3), .b(n_1384), .o(n_1433) );
BUF_X2 newInst_618 ( .a(newNet_371), .o(newNet_618) );
AND2_X1 g60335 ( .a(n_612), .b(n_64), .o(n_861) );
XOR2_X1 g60163 ( .a(n_520), .b(pmem_d_0), .o(n_973) );
NOR2_Z1 g35161 ( .a(n_3201), .b(n_3232), .o(Rd_3_) );
BUF_X2 newInst_980 ( .a(newNet_979), .o(newNet_980) );
NAND2_Z01 g34806 ( .a(n_3573), .b(U_2_), .o(n_3757) );
NAND2_Z01 g58464 ( .a(n_2435), .b(n_2593), .o(n_2632) );
NOR3_Z1 g59528 ( .a(n_1123), .b(n_1465), .c(n_933), .o(n_1599) );
INV_X1 g60011 ( .a(n_1118), .o(n_1119) );
NAND2_Z01 g60907 ( .a(PC_3_), .b(pmem_d_6), .o(n_232) );
NAND2_Z01 g34917 ( .a(n_3634), .b(n_3224), .o(n_3646) );
INV_X1 g35260 ( .a(n_4531), .o(n_3414) );
INV_X1 g35480 ( .a(pmem_d_4), .o(n_3244) );
BUF_X2 newInst_427 ( .a(newNet_426), .o(newNet_427) );
XOR2_X1 g34251 ( .a(n_4180), .b(SP_8_), .o(n_4282) );
INV_X1 g34503 ( .a(n_4040), .o(n_4041) );
AND2_X1 g35352 ( .a(n_4482), .b(n_3286), .o(n_3353) );
BUF_X2 newInst_496 ( .a(newNet_495), .o(newNet_496) );
BUF_X2 newInst_684 ( .a(newNet_461), .o(newNet_684) );
BUF_X2 newInst_87 ( .a(newNet_86), .o(newNet_87) );
AND2_X1 g59239 ( .a(n_1831), .b(n_1036), .o(n_1866) );
NAND2_Z02 g35244 ( .a(n_3359), .b(n_3346), .o(n_4651) );
fflopd pY_reg_0_ ( .CK(newNet_193), .D(n_2731), .Q(pY_0_) );
NOR2_Z1 g35168 ( .a(n_3445), .b(n_3358), .o(n_3456) );
NAND2_Z01 g58469 ( .a(n_2388), .b(n_2587), .o(n_2627) );
NAND4_Z1 g59377 ( .a(n_773), .b(n_1474), .c(n_1655), .d(n_1362), .o(n_1741) );
BUF_X2 newInst_1263 ( .a(newNet_1262), .o(newNet_1263) );
BUF_X2 newInst_175 ( .a(newNet_124), .o(newNet_175) );
fflopd SP_reg_0_ ( .CK(newNet_574), .D(n_1594), .Q(SP_0_) );
AND2_X1 g60079 ( .a(n_845), .b(n_59), .o(n_1056) );
INV_X1 g61052 ( .a(pX_10_), .o(n_100) );
NAND2_Z01 g58553 ( .a(n_2494), .b(pY_9_), .o(n_2544) );
NAND2_Z01 g35055 ( .a(n_3504), .b(n_3308), .o(n_3528) );
XOR2_X1 g35382 ( .a(PC_0_), .b(PC_1_), .o(n_4553) );
BUF_X2 newInst_1410 ( .a(newNet_1409), .o(newNet_1410) );
NAND2_Z01 g58042 ( .a(n_2902), .b(n_2437), .o(n_2943) );
BUF_X2 newInst_692 ( .a(newNet_691), .o(newNet_692) );
fflopd GPR_reg_0__1_ ( .CK(newNet_1812), .D(n_2733), .Q(GPR_0__1_) );
NAND2_Z01 g60765 ( .a(n_247), .b(pmem_d_1), .o(n_458) );
BUF_X2 newInst_206 ( .a(newNet_205), .o(newNet_206) );
BUF_X2 newInst_969 ( .a(newNet_968), .o(newNet_969) );
NAND4_Z1 g34592 ( .a(n_3672), .b(n_3719), .c(n_3654), .d(n_3819), .o(n_3968) );
NOR2_Z1 g58342 ( .a(n_2687), .b(n_1735), .o(n_2727) );
AND4_X1 g34499 ( .a(n_3987), .b(n_3989), .c(n_3988), .d(n_3986), .o(n_4045) );
BUF_X2 newInst_624 ( .a(newNet_623), .o(newNet_624) );
BUF_X2 newInst_559 ( .a(newNet_558), .o(newNet_559) );
NAND4_Z1 g34076 ( .a(n_4269), .b(n_4131), .c(n_4379), .d(n_4250), .o(n_4396) );
BUF_X2 newInst_650 ( .a(newNet_444), .o(newNet_650) );
NAND2_Z01 g60197 ( .a(n_640), .b(n_561), .o(n_948) );
fflopd GPR_reg_5__1_ ( .CK(newNet_871), .D(n_2744), .Q(GPR_5__1_) );
NAND2_Z01 final_adder_mux_R16_278_6_g425 ( .a(n_4437), .b(n_4421), .o(final_adder_mux_R16_278_6_n_23) );
BUF_X2 newInst_34 ( .a(newNet_33), .o(newNet_34) );
NAND4_Z1 g58412 ( .a(n_1244), .b(n_2450), .c(n_2576), .d(n_1280), .o(n_2658) );
BUF_X2 newInst_1429 ( .a(newNet_1428), .o(newNet_1429) );
NAND2_Z01 g58788 ( .a(n_2200), .b(GPR_7__7_), .o(n_2312) );
NAND2_Z01 g34725 ( .a(n_3591), .b(U_5_), .o(n_3840) );
NAND2_Z01 g59261 ( .a(n_1786), .b(n_1103), .o(n_1849) );
XOR2_X1 final_adder_mux_R16_278_6_g419 ( .a(n_4440), .b(n_4424), .o(final_adder_mux_R16_278_6_n_30) );
BUF_X2 newInst_1327 ( .a(newNet_1326), .o(newNet_1327) );
AND2_X1 final_adder_mux_R16_278_6_g449 ( .a(n_4447), .b(n_4431), .o(final_adder_mux_R16_278_6_n_0) );
BUF_X2 newInst_276 ( .a(newNet_275), .o(newNet_276) );
NAND2_Z01 g60994 ( .a(n_91), .b(n_47), .o(n_141) );
BUF_X2 newInst_1198 ( .a(newNet_192), .o(newNet_1198) );
AND2_X1 g58111 ( .a(n_2850), .b(n_2213), .o(n_2901) );
XOR2_X1 final_adder_mux_R16_278_6_g402 ( .a(final_adder_mux_R16_278_6_n_36), .b(final_adder_mux_R16_278_6_n_28), .o(R16_1_) );
NAND2_Z01 g35435 ( .a(n_3231), .b(n_3249), .o(n_4490) );
NAND2_Z01 g60944 ( .a(io_do_4), .b(n_65), .o(n_207) );
AND2_X1 g59139 ( .a(n_1893), .b(n_1220), .o(n_1983) );
NOR3_Z1 g58544 ( .a(n_569), .b(n_2527), .c(n_176), .o(n_2554) );
BUF_X2 newInst_1712 ( .a(newNet_1711), .o(newNet_1712) );
NAND2_Z01 g34265 ( .a(n_4176), .b(pX_9_), .o(n_4268) );
NAND2_Z01 g60686 ( .a(n_198), .b(GPR_21__4_), .o(n_452) );
NOR2_Z1 g59938 ( .a(n_1110), .b(n_61), .o(n_1186) );
NAND2_Z01 g58236 ( .a(n_2753), .b(n_2217), .o(n_2831) );
NAND2_Z01 g58163 ( .a(n_2803), .b(n_2377), .o(n_2847) );
NAND2_Z01 g60505 ( .a(Rd_1_), .b(n_345), .o(n_641) );
NAND2_Z01 g58573 ( .a(n_2479), .b(n_2051), .o(n_2523) );
BUF_X2 newInst_1044 ( .a(newNet_1043), .o(newNet_1044) );
BUF_X2 newInst_348 ( .a(newNet_347), .o(newNet_348) );
INV_X1 g59554 ( .a(n_1573), .o(n_1572) );
NAND4_Z1 g60381 ( .a(n_398), .b(n_412), .c(n_415), .d(n_426), .o(n_764) );
NAND2_Z01 g58864 ( .a(n_2156), .b(GPR_15__3_), .o(n_2243) );
BUF_X2 newInst_641 ( .a(newNet_199), .o(newNet_641) );
BUF_X2 newInst_376 ( .a(newNet_375), .o(newNet_376) );
NAND2_Z01 g34296 ( .a(n_4166), .b(n_4541), .o(n_4238) );
BUF_X2 newInst_470 ( .a(newNet_469), .o(newNet_470) );
INV_X1 g58888 ( .a(n_2198), .o(n_2197) );
NAND2_Z01 g58160 ( .a(n_2805), .b(n_2393), .o(n_2853) );
BUF_X2 newInst_502 ( .a(newNet_501), .o(newNet_502) );
NOR2_Z1 g59339 ( .a(n_1701), .b(n_62), .o(n_1777) );
BUF_X2 newInst_5 ( .a(newNet_4), .o(newNet_5) );
NAND2_Z01 g59864 ( .a(n_1164), .b(n_63), .o(n_1262) );
NAND4_Z1 g58490 ( .a(n_1154), .b(n_2074), .c(n_2556), .d(n_1250), .o(n_2606) );
NAND2_Z01 g58691 ( .a(n_2214), .b(GPR_16__3_), .o(n_2415) );
NAND2_Z01 g34404 ( .a(n_3208), .b(pZ_8_), .o(n_4134) );
NAND2_Z01 g61023 ( .a(n_40), .b(n_39), .o(n_162) );
BUF_X2 newInst_1177 ( .a(newNet_1176), .o(newNet_1177) );
AND3_X1 g58569 ( .a(n_1977), .b(n_2504), .c(n_2003), .o(n_2529) );
INV_X1 g60529 ( .a(n_610), .o(n_611) );
AND2_X1 g35427 ( .a(n_3262), .b(state_0_), .o(n_4557) );
BUF_X2 newInst_1129 ( .a(newNet_1128), .o(newNet_1129) );
NAND2_Z01 g58751 ( .a(n_2204), .b(GPR_3__3_), .o(n_2349) );
NAND2_Z01 g58243 ( .a(n_2754), .b(n_2216), .o(n_2824) );
AND2_X1 g57895 ( .a(n_3009), .b(n_2210), .o(n_3043) );
fflopd GPR_reg_7__5_ ( .CK(newNet_756), .D(n_2998), .Q(GPR_7__5_) );
BUF_X2 newInst_418 ( .a(newNet_417), .o(newNet_418) );
NOR2_Z1 g60973 ( .a(n_4444), .b(n_4428), .o(n_149) );
XOR2_X1 g35257 ( .a(n_3277), .b(pX_2_), .o(n_4572) );
BUF_X2 newInst_326 ( .a(newNet_325), .o(newNet_326) );
AND2_X1 g35346 ( .a(n_3297), .b(n_3249), .o(n_3357) );
XNOR2_X1 g35021 ( .a(n_3529), .b(pmem_d_11), .o(n_3555) );
BUF_X2 newInst_1314 ( .a(newNet_1313), .o(newNet_1314) );
AND2_X1 g60640 ( .a(n_177), .b(n_331), .o(n_496) );
AND3_X1 g35139 ( .a(n_4491), .b(n_4634), .c(n_3259), .o(n_3479) );
BUF_X2 newInst_322 ( .a(newNet_321), .o(newNet_322) );
AND2_X1 g58394 ( .a(n_2657), .b(n_2202), .o(n_2674) );
BUF_X2 newInst_528 ( .a(newNet_527), .o(newNet_528) );
BUF_X2 newInst_750 ( .a(newNet_749), .o(newNet_750) );
BUF_X2 newInst_1029 ( .a(newNet_1028), .o(newNet_1029) );
BUF_X2 newInst_837 ( .a(newNet_836), .o(newNet_837) );
INV_X2 newInst_1785 ( .a(newNet_1784), .o(newNet_1785) );
NOR2_Z2 g34920 ( .a(n_3588), .b(rst), .o(n_3769) );
AND3_X1 g60371 ( .a(n_376), .b(n_346), .c(n_71), .o(n_842) );
fflopd GPR_reg_9__5_ ( .CK(newNet_670), .D(n_2996), .Q(GPR_9__5_) );
AND3_X1 g60147 ( .a(n_500), .b(n_346), .c(n_4490), .o(n_1029) );
AND2_X1 g60761 ( .a(n_4624), .b(n_251), .o(n_384) );
fflopd pZ_reg_5_ ( .CK(newNet_74), .D(n_3094), .Q(pZ_5_) );
NAND4_Z1 g59445 ( .a(n_1544), .b(n_1429), .c(n_1618), .d(n_986), .o(n_1677) );
NAND2_Z01 g58623 ( .a(n_2284), .b(n_1795), .o(n_2474) );
NOR2_Z1 g60115 ( .a(n_776), .b(n_450), .o(n_1011) );
AND2_X1 g59176 ( .a(n_1872), .b(n_1875), .o(n_1975) );
BUF_X2 newInst_554 ( .a(newNet_553), .o(newNet_554) );
BUF_X2 newInst_711 ( .a(newNet_710), .o(newNet_711) );
BUF_X2 newInst_745 ( .a(newNet_744), .o(newNet_745) );
BUF_X2 newInst_1116 ( .a(newNet_1115), .o(newNet_1116) );
NAND4_Z1 g59544 ( .a(n_1157), .b(n_1345), .c(n_1401), .d(n_576), .o(n_1584) );
NAND2_Z01 g35276 ( .a(U_1_), .b(n_3275), .o(n_3399) );
NAND2_Z01 g59098 ( .a(n_1871), .b(n_363), .o(n_2010) );
BUF_X2 newInst_960 ( .a(newNet_959), .o(newNet_960) );
NOR4_Z1 g35140 ( .a(n_4652), .b(n_3320), .c(n_4651), .d(n_3327), .o(n_3478) );
BUF_X2 newInst_935 ( .a(newNet_488), .o(newNet_935) );
NOR2_Z1 g34187 ( .a(n_4324), .b(n_4614), .o(n_4428) );
INV_X1 drc_bufs61216 ( .a(n_23), .o(n_11) );
NOR2_Z1 g60354 ( .a(n_564), .b(rst), .o(n_854) );
XNOR2_X1 g60858 ( .a(n_54), .b(n_40), .o(n_286) );
AND2_X1 g58596 ( .a(n_2459), .b(n_94), .o(n_2499) );
BUF_X2 newInst_988 ( .a(newNet_987), .o(newNet_988) );
BUF_X2 newInst_594 ( .a(newNet_593), .o(newNet_594) );
BUF_X2 newInst_38 ( .a(newNet_37), .o(newNet_38) );
BUF_X2 newInst_1801 ( .a(newNet_1800), .o(newNet_1801) );
BUF_X2 newInst_971 ( .a(newNet_970), .o(newNet_971) );
AND2_X1 g59775 ( .a(n_1306), .b(PC_8_), .o(n_1382) );
BUF_X2 newInst_1485 ( .a(newNet_1484), .o(newNet_1485) );
AND2_X1 g60758 ( .a(n_40), .b(n_165), .o(n_385) );
NAND2_Z01 g34870 ( .a(n_3584), .b(GPR_21__3_), .o(n_3693) );
fflopd GPR_reg_19__6_ ( .CK(newNet_1279), .D(n_3081), .Q(GPR_19__6_) );
BUF_X2 newInst_264 ( .a(newNet_263), .o(newNet_264) );
NAND2_Z01 g34650 ( .a(n_3768), .b(n_4549), .o(n_3910) );
fflopd GPR_reg_0__3_ ( .CK(newNet_1793), .D(n_2838), .Q(GPR_0__3_) );
NAND2_Z01 g57839 ( .a(n_3037), .b(n_2346), .o(n_3071) );
NAND2_Z01 g34484 ( .a(n_4041), .b(SP_1_), .o(n_4059) );
NAND3_Z1 g35172 ( .a(n_3248), .b(n_3359), .c(pmem_d_13), .o(n_4641) );
NOR2_Z1 g60308 ( .a(n_615), .b(n_124), .o(n_867) );
NAND2_Z01 g57832 ( .a(n_3044), .b(n_2416), .o(n_3081) );
BUF_X2 newInst_570 ( .a(newNet_569), .o(newNet_570) );
NAND2_Z01 g59703 ( .a(io_do_6), .b(n_1353), .o(n_1427) );
BUF_X2 newInst_1770 ( .a(newNet_1769), .o(newNet_1770) );
NOR2_Z1 g59094 ( .a(n_1869), .b(n_1082), .o(n_2061) );
AND2_X1 g35046 ( .a(n_3525), .b(n_3474), .o(n_4648) );
BUF_X2 newInst_769 ( .a(newNet_768), .o(newNet_769) );
BUF_X2 newInst_1419 ( .a(newNet_1418), .o(newNet_1419) );
BUF_X2 newInst_893 ( .a(newNet_892), .o(newNet_893) );
NAND2_Z01 g57802 ( .a(n_3080), .b(n_13), .o(n_3105) );
BUF_X2 newInst_877 ( .a(newNet_876), .o(newNet_877) );
NAND2_Z01 g60479 ( .a(n_20), .b(Rd_r_3_), .o(n_667) );
NAND2_Z01 g59149 ( .a(n_1896), .b(n_1454), .o(n_1950) );
BUF_X2 newInst_510 ( .a(newNet_509), .o(newNet_510) );
fflopd SP_reg_11_ ( .CK(newNet_555), .D(n_1809), .Q(SP_11_) );
AND2_X1 g58008 ( .a(n_2940), .b(n_2200), .o(n_2963) );
BUF_X2 newInst_1341 ( .a(newNet_1340), .o(newNet_1341) );
NAND2_Z01 g59351 ( .a(n_31), .b(n_62), .o(n_1762) );
INV_X1 g59479 ( .a(n_1647), .o(n_1646) );
BUF_X2 newInst_612 ( .a(newNet_611), .o(newNet_612) );
NAND2_Z01 g34839 ( .a(n_3636), .b(GPR_10__1_), .o(n_3724) );
BUF_X2 newInst_1424 ( .a(newNet_1227), .o(newNet_1424) );
AND3_X1 g59800 ( .a(n_47), .b(n_1208), .c(pmem_d_6), .o(n_1347) );
AND2_X1 g59275 ( .a(n_61), .b(n_6), .o(n_1838) );
fflopd state_reg_2_ ( .CK(newNet_16), .D(n_1376), .Q(state_2_) );
AND2_X1 g57988 ( .a(n_2940), .b(n_2159), .o(n_2983) );
NAND4_Z1 g59807 ( .a(n_648), .b(n_677), .c(n_1176), .d(n_710), .o(n_1321) );
NAND2_Z01 g57826 ( .a(n_3050), .b(n_2249), .o(n_3087) );
AND2_X1 g59782 ( .a(n_1308), .b(n_1270), .o(n_1350) );
BUF_X2 newInst_166 ( .a(newNet_165), .o(newNet_166) );
NAND2_Z01 g59768 ( .a(n_1268), .b(n_976), .o(n_1359) );
fflopd GPR_reg_12__1_ ( .CK(newNet_1667), .D(n_2783), .Q(GPR_12__1_) );
BUF_X2 newInst_1651 ( .a(newNet_1650), .o(newNet_1651) );
BUF_X2 newInst_733 ( .a(newNet_732), .o(newNet_733) );
BUF_X2 newInst_47 ( .a(newNet_46), .o(newNet_47) );
NAND2_Z01 g58602 ( .a(n_2459), .b(n_1945), .o(n_2493) );
NOR3_Z1 g59654 ( .a(n_1127), .b(n_1443), .c(n_1126), .o(n_1471) );
NAND2_Z01 g58295 ( .a(n_2703), .b(n_2244), .o(n_2775) );
AND2_X1 g57898 ( .a(n_3009), .b(n_2207), .o(n_3040) );
NAND2_Z01 g34154 ( .a(n_4317), .b(n_4616), .o(n_4354) );
NAND2_Z01 g60565 ( .a(n_357), .b(pZ_12_), .o(n_543) );
fflopd pY_reg_12_ ( .CK(newNet_175), .D(n_3028), .Q(pY_12_) );
INV_X1 g60280 ( .a(n_858), .o(n_857) );
BUF_X2 newInst_486 ( .a(newNet_485), .o(newNet_486) );
BUF_X2 newInst_925 ( .a(newNet_924), .o(newNet_925) );
BUF_X2 newInst_759 ( .a(newNet_758), .o(newNet_759) );
NAND4_Z1 g58562 ( .a(n_1518), .b(n_1439), .c(n_2448), .d(n_1062), .o(n_2536) );
NAND2_Z01 g57928 ( .a(n_2979), .b(n_2227), .o(n_3017) );
NAND2_Z01 g58290 ( .a(n_2707), .b(n_2251), .o(n_2780) );
AND2_X1 g58269 ( .a(n_2752), .b(n_2201), .o(n_2798) );
NAND4_Z1 g34582 ( .a(n_3678), .b(n_3776), .c(n_3876), .d(n_3775), .o(n_3978) );
BUF_X2 newInst_1539 ( .a(newNet_1538), .o(newNet_1539) );
NAND4_Z1 g60154 ( .a(n_733), .b(n_740), .c(n_736), .d(n_652), .o(n_981) );
NAND3_Z2 g60126 ( .a(n_43), .b(n_605), .c(pmem_d_10), .o(n_1036) );
NAND2_Z01 g58885 ( .a(n_2140), .b(GPR_9__1_), .o(n_2222) );
BUF_X2 newInst_566 ( .a(newNet_451), .o(newNet_566) );
BUF_X2 newInst_577 ( .a(newNet_576), .o(newNet_577) );
NAND3_Z1 g34449 ( .a(n_3855), .b(n_4052), .c(n_3856), .o(n_4091) );
NOR3_Z1 g60133 ( .a(n_4650), .b(n_569), .c(n_4663), .o(n_999) );
AND2_X1 g58383 ( .a(n_2656), .b(n_2208), .o(n_2685) );
NAND2_Z01 g58903 ( .a(n_2123), .b(io_do_5), .o(n_2180) );
fflopd S_reg ( .CK(newNet_454), .D(n_3194), .Q(S) );
NAND2_Z01 g59005 ( .a(n_1990), .b(n_1712), .o(n_2114) );
NOR2_Z1 g34280 ( .a(n_4163), .b(n_3251), .o(n_4253) );
NOR2_Z1 g34315 ( .a(n_16064_BAR), .b(n_3521), .o(n_4218) );
NAND4_Z1 g57654 ( .a(n_1961), .b(n_2469), .c(n_3179), .d(n_2025), .o(n_3188) );
NAND2_Z01 g59403 ( .a(io_do_1), .b(n_1664), .o(n_1713) );
BUF_X2 newInst_312 ( .a(newNet_311), .o(newNet_312) );
AND3_X1 g59991 ( .a(n_113), .b(n_1114), .c(pY_7_), .o(n_1138) );
AND2_X1 g58268 ( .a(n_2752), .b(n_2202), .o(n_2799) );
NOR2_Z2 g60964 ( .a(n_59), .b(pmem_d_3), .o(n_198) );
BUF_X2 newInst_1096 ( .a(newNet_1095), .o(newNet_1096) );
INV_X1 g60530 ( .a(n_608), .o(n_609) );
BUF_X2 newInst_569 ( .a(newNet_568), .o(newNet_569) );
AND2_X1 g57889 ( .a(n_3009), .b(n_2155), .o(n_3049) );
NAND2_Z01 g58693 ( .a(n_2210), .b(GPR_1__0_), .o(n_2413) );
XNOR2_X1 g60852 ( .a(n_4441), .b(n_4425), .o(n_334) );
NAND2_Z01 g34145 ( .a(n_4325), .b(n_4627), .o(n_4363) );
fflopd GPR_reg_15__2_ ( .CK(newNet_1511), .D(n_2775), .Q(GPR_15__2_) );
NAND2_Z01 g58555 ( .a(n_2493), .b(pZ_9_), .o(n_2542) );
BUF_X2 newInst_1068 ( .a(newNet_226), .o(newNet_1068) );
NAND2_Z01 g34330 ( .a(n_4166), .b(n_4553), .o(n_4204) );
NAND2_Z01 g58299 ( .a(n_2697), .b(n_2428), .o(n_2771) );
NOR2_Z1 g59581 ( .a(n_1485), .b(n_1386), .o(n_1550) );
NAND2_Z01 g34393 ( .a(n_3208), .b(pZ_1_), .o(n_4145) );
NAND2_Z01 g34653 ( .a(n_3768), .b(n_4555), .o(n_3907) );
NAND2_Z01 g59750 ( .a(n_1294), .b(n_209), .o(n_1389) );
NOR2_Z1 g35370 ( .a(n_3287), .b(n_3286), .o(n_3320) );
BUF_X2 newInst_1630 ( .a(newNet_851), .o(newNet_1630) );
NAND2_Z01 g34561 ( .a(n_3906), .b(n_3352), .o(n_4649) );
AND2_X1 g59957 ( .a(n_1048), .b(io_do_6), .o(n_1199) );
AND2_X1 final_adder_mux_R16_278_6_g439 ( .a(n_4449), .b(n_4433), .o(final_adder_mux_R16_278_6_n_10) );
NAND2_Z01 g34671 ( .a(n_3619), .b(n_3618), .o(n_3894) );
AND2_X1 g60580 ( .a(n_463), .b(n_68), .o(n_612) );
NAND4_Z1 g59442 ( .a(n_813), .b(n_804), .c(n_1597), .d(n_881), .o(n_1678) );
NAND2_Z01 g60456 ( .a(n_360), .b(GPR_1__0_), .o(n_690) );
XOR2_X1 g35073 ( .a(n_3485), .b(pX_6_), .o(n_3520) );
INV_X1 g35482 ( .a(SP_6_), .o(n_3242) );
BUF_X2 newInst_1717 ( .a(newNet_1716), .o(newNet_1717) );
BUF_X2 newInst_143 ( .a(newNet_142), .o(newNet_143) );
NAND2_Z01 g58237 ( .a(n_2756), .b(n_2217), .o(n_2830) );
INV_X1 g35426 ( .a(n_3275), .o(n_4640) );
INV_X1 g61106 ( .a(n_4521), .o(n_46) );
NOR2_Z1 g59880 ( .a(n_1219), .b(n_344), .o(n_1247) );
NAND2_Z01 g60182 ( .a(n_627), .b(n_703), .o(n_958) );
INV_X1 g58381 ( .a(n_2687), .o(n_2688) );
NOR2_Z1 g58275 ( .a(n_2727), .b(n_2728), .o(n_2792) );
BUF_X2 newInst_7 ( .a(newNet_6), .o(newNet_7) );
NAND2_Z01 g35030 ( .a(n_3518), .b(n_3464), .o(n_3541) );
fflopd pY_reg_9_ ( .CK(newNet_121), .D(n_2876), .Q(pY_9_) );
NAND2_Z01 g59932 ( .a(n_1045), .b(n_969), .o(n_1212) );
NAND2_Z01 g57653 ( .a(n_3181), .b(n_1771), .o(n_3189) );
AND2_X1 g59028 ( .a(n_1904), .b(n_1619), .o(n_2076) );
BUF_X2 newInst_1352 ( .a(newNet_1351), .o(newNet_1352) );
BUF_X2 newInst_509 ( .a(newNet_508), .o(newNet_509) );
NAND4_Z2 g35181 ( .a(n_3367), .b(n_3378), .c(n_3361), .d(n_3400), .o(n_4616) );
NOR2_Z1 g59290 ( .a(n_19), .b(n_1738), .o(n_1820) );
INV_Z1 g16813 ( .a(GPR_1__0_), .o(n_4410) );
BUF_X2 newInst_839 ( .a(newNet_838), .o(newNet_839) );
NAND2_Z01 g60741 ( .a(SP_12_), .b(n_180), .o(n_399) );
AND2_X1 g59526 ( .a(n_1571), .b(pX_12_), .o(n_1603) );
NAND2_Z01 g58246 ( .a(n_2755), .b(n_2198), .o(n_2821) );
NAND2_Z01 g35246 ( .a(n_3356), .b(n_3263), .o(n_3428) );
NOR2_Z1 g34267 ( .a(n_4175), .b(n_3253), .o(n_4266) );
NAND2_Z01 g34875 ( .a(n_3571), .b(GPR_20__7_), .o(n_3688) );
INV_X1 g60092 ( .a(n_1033), .o(n_1034) );
BUF_X2 newInst_1147 ( .a(newNet_1146), .o(newNet_1147) );
BUF_X2 newInst_754 ( .a(newNet_753), .o(newNet_754) );
BUF_X2 newInst_1601 ( .a(newNet_1600), .o(newNet_1601) );
BUF_X2 newInst_519 ( .a(newNet_518), .o(newNet_519) );
NAND3_Z1 g59410 ( .a(n_145), .b(n_1608), .c(n_4627), .o(n_1708) );
BUF_X2 newInst_1433 ( .a(newNet_1432), .o(newNet_1433) );
XOR2_X1 g35104 ( .a(n_4622), .b(n_3236), .o(n_4467) );
BUF_X2 newInst_762 ( .a(newNet_761), .o(newNet_762) );
NAND2_Z01 g35411 ( .a(pY_5_), .b(pmem_d_13), .o(n_3293) );
XOR2_X1 g34657 ( .a(n_3593), .b(n_3222), .o(n_4587) );
BUF_X2 newInst_1190 ( .a(newNet_1189), .o(newNet_1190) );
NAND2_Z01 g34842 ( .a(n_3586), .b(GPR_9__1_), .o(n_3721) );
NAND2_Z01 g60339 ( .a(n_11), .b(pmem_d_3), .o(n_791) );
NAND2_Z01 g58626 ( .a(n_2353), .b(n_2014), .o(n_2483) );
fflopd GPR_reg_17__2_ ( .CK(newNet_1400), .D(n_2777), .Q(GPR_17__2_) );
BUF_X2 newInst_434 ( .a(newNet_433), .o(newNet_434) );
NAND2_Z01 g60313 ( .a(n_570), .b(pZ_6_), .o(n_813) );
NAND2_Z01 g57981 ( .a(n_2941), .b(n_2218), .o(n_2991) );
NAND2_Z01 g59939 ( .a(n_1109), .b(pmem_d_3), .o(n_1185) );
INV_X2 newInst_892 ( .a(newNet_891), .o(newNet_892) );
NOR3_Z1 g58491 ( .a(n_315), .b(n_2574), .c(n_386), .o(n_2605) );
BUF_X2 newInst_702 ( .a(newNet_701), .o(newNet_702) );
NAND2_Z01 g34157 ( .a(n_4317), .b(n_4622), .o(n_4351) );
BUF_X2 newInst_690 ( .a(newNet_689), .o(newNet_690) );
NAND2_Z01 g60296 ( .a(n_598), .b(GPR_15__5_), .o(n_828) );
INV_X1 g59910 ( .a(n_1212), .o(n_1213) );
AND2_X1 g35348 ( .a(n_4633), .b(pmem_d_9), .o(n_4491) );
NAND2_Z01 g60257 ( .a(n_596), .b(GPR_3__2_), .o(n_889) );
fflopd GPR_reg_11__0_ ( .CK(newNet_1710), .D(n_2638), .Q(GPR_11__0_) );
BUF_X2 newInst_878 ( .a(newNet_396), .o(newNet_878) );
NOR2_Z1 g34430 ( .a(n_4610), .b(n_4609), .o(n_4107) );
fflopd SP_reg_4_ ( .CK(newNet_492), .D(n_1674), .Q(SP_4_) );
NAND2_Z01 g58880 ( .a(n_2155), .b(GPR_14__5_), .o(n_2227) );
BUF_X2 newInst_944 ( .a(newNet_943), .o(newNet_944) );
AND2_X1 g59122 ( .a(n_55), .b(n_1877), .o(n_1989) );
fflopd GPR_reg_20__0_ ( .CK(newNet_1209), .D(n_2629), .Q(GPR_20__0_) );
NAND2_Z01 g59093 ( .a(n_1872), .b(n_1486), .o(n_2014) );
NOR2_Z1 g59110 ( .a(n_1893), .b(n_1447), .o(n_1999) );
BUF_X2 newInst_1197 ( .a(newNet_1196), .o(newNet_1197) );
AND2_X1 g34407 ( .a(n_4082), .b(n_4088), .o(n_4131) );
NAND2_Z01 g59514 ( .a(n_1549), .b(pmem_d_8), .o(n_1625) );
AND2_X1 g61020 ( .a(n_4489), .b(pmem_d_1), .o(n_165) );
XOR2_X1 g59904 ( .a(n_970), .b(pmem_d_2), .o(n_1226) );
NAND2_Z01 g35265 ( .a(U_11_), .b(n_3275), .o(n_3408) );
NAND2_Z01 g59147 ( .a(n_1871), .b(n_610), .o(n_1952) );
NAND2_Z01 g34466 ( .a(n_4060), .b(SP_2_), .o(n_4076) );
INV_X1 g61034 ( .a(SP_2_), .o(n_118) );
NAND2_Z01 g58600 ( .a(n_2479), .b(n_1958), .o(n_2495) );
NAND2_Z01 g58668 ( .a(n_2214), .b(GPR_16__2_), .o(n_2438) );
AND3_X1 g59042 ( .a(n_51), .b(n_1983), .c(pY_11_), .o(n_2067) );
BUF_X2 newInst_584 ( .a(newNet_583), .o(newNet_584) );
NAND2_Z01 g60288 ( .a(R16_5_), .b(n_14), .o(n_836) );
fflopd GPR_reg_8__4_ ( .CK(newNet_703), .D(n_2924), .Q(GPR_8__4_) );
fflopd GPR_reg_23__1_ ( .CK(newNet_1056), .D(n_2759), .Q(GPR_23__1_) );
BUF_X2 newInst_402 ( .a(newNet_401), .o(newNet_402) );
fflopd U_reg_0_ ( .CK(newNet_442), .D(n_2719), .Q(U_0_) );
AND2_X1 g58393 ( .a(n_2656), .b(n_2203), .o(n_2675) );
BUF_X2 newInst_1446 ( .a(newNet_1445), .o(newNet_1446) );
BUF_X2 newInst_1783 ( .a(newNet_1782), .o(newNet_1783) );
NAND2_Z01 g60481 ( .a(n_374), .b(GPR_12__7_), .o(n_665) );
BUF_X2 newInst_1336 ( .a(newNet_845), .o(newNet_1336) );
BUF_X2 newInst_923 ( .a(newNet_615), .o(newNet_923) );
INV_X1 g35093 ( .a(n_3499), .o(n_4605) );
NAND4_Z1 g60143 ( .a(n_629), .b(n_695), .c(n_656), .d(n_669), .o(n_989) );
NOR2_Z1 g61004 ( .a(io_do_0), .b(pmem_d_0), .o(n_135) );
NAND2_Z01 g34765 ( .a(n_3631), .b(GPR_11__4_), .o(n_3800) );
NAND2_Z01 g34914 ( .a(n_3633), .b(pZ_10_), .o(n_3649) );
BUF_X2 newInst_1459 ( .a(newNet_1458), .o(newNet_1459) );
BUF_X2 newInst_1057 ( .a(newNet_737), .o(newNet_1057) );
NAND3_Z1 g35192 ( .a(n_3377), .b(n_3436), .c(n_3410), .o(n_4627) );
BUF_X2 newInst_1553 ( .a(newNet_1552), .o(newNet_1553) );
NAND4_Z1 g34576 ( .a(n_3658), .b(n_3805), .c(n_3807), .d(n_3806), .o(n_3984) );
AND2_X1 g57993 ( .a(n_2940), .b(n_2156), .o(n_2978) );
NOR2_Z1 g59867 ( .a(n_1162), .b(pmem_d_0), .o(n_1270) );
BUF_X2 newInst_1019 ( .a(newNet_506), .o(newNet_1019) );
NAND2_Z01 g58296 ( .a(n_2701), .b(n_2439), .o(n_2774) );
AND3_X1 g60124 ( .a(n_109), .b(n_609), .c(SP_5_), .o(n_1003) );
BUF_X2 newInst_505 ( .a(newNet_504), .o(newNet_505) );
NAND2_Z01 g34816 ( .a(n_3568), .b(GPR_22__2_), .o(n_3747) );
XOR2_X1 g35258 ( .a(n_3276), .b(pY_2_), .o(n_3420) );
NAND4_Z1 g58015 ( .a(n_2067), .b(n_2545), .c(n_2915), .d(n_2052), .o(n_2957) );
BUF_X2 newInst_1356 ( .a(newNet_1355), .o(newNet_1356) );
BUF_X2 newInst_681 ( .a(newNet_680), .o(newNet_681) );
INV_X1 g59383 ( .a(n_1730), .o(n_1731) );
NOR4_Z1 g59375 ( .a(n_4490), .b(n_346), .c(n_1592), .d(pmem_d_7), .o(n_1743) );
fflopd GPR_reg_18__5_ ( .CK(newNet_1338), .D(n_3013), .Q(GPR_18__5_) );
fflopd GPR_reg_2__2_ ( .CK(newNet_1012), .D(n_2749), .Q(GPR_2__2_) );
fflopd pY_reg_1_ ( .CK(newNet_158), .D(n_2878), .Q(pY_1_) );
NOR2_Z1 g35025 ( .a(n_3527), .b(n_3216), .o(n_3554) );
NAND2_Z01 g60196 ( .a(n_641), .b(n_558), .o(n_949) );
NAND3_Z1 g34556 ( .a(n_3695), .b(n_3697), .c(n_3696), .o(n_4003) );
NOR3_Z1 g35141 ( .a(n_3254), .b(n_3446), .c(pmem_d_3), .o(n_4665) );
XOR2_X1 g57661 ( .a(n_3158), .b(n_3078), .o(n_3181) );
AND2_X1 g57894 ( .a(n_3009), .b(n_2211), .o(n_3044) );
BUF_X2 newInst_274 ( .a(newNet_273), .o(newNet_274) );
NAND2_Z01 g58328 ( .a(n_2666), .b(n_2231), .o(n_2737) );
NAND2_Z01 g59231 ( .a(n_1833), .b(n_1014), .o(n_1881) );
INV_X1 g59345 ( .a(n_1767), .o(n_1768) );
INV_X1 g35469 ( .a(pY_8_), .o(n_3255) );
INV_X1 g35324 ( .a(n_3345), .o(n_4596) );
NAND2_Z01 g60463 ( .a(n_457), .b(GPR_16__0_), .o(n_683) );
NAND4_Z1 g59809 ( .a(n_683), .b(n_684), .c(n_1174), .d(n_651), .o(n_1319) );
NOR3_Z1 g59802 ( .a(n_1167), .b(n_1032), .c(n_1164), .o(n_1346) );
BUF_X2 newInst_933 ( .a(newNet_932), .o(newNet_933) );
NAND2_Z01 g34830 ( .a(n_3572), .b(GPR_4__1_), .o(n_3733) );
AND2_X1 g60754 ( .a(n_109), .b(n_204), .o(n_388) );
BUF_X2 newInst_1775 ( .a(newNet_688), .o(newNet_1775) );
BUF_X2 newInst_843 ( .a(newNet_842), .o(newNet_843) );
BUF_X2 newInst_1803 ( .a(newNet_1802), .o(newNet_1803) );
BUF_X2 newInst_1700 ( .a(newNet_1699), .o(newNet_1700) );
NAND2_Z01 g58821 ( .a(n_31), .b(n_2164), .o(n_2284) );
INV_X1 g60539 ( .a(n_581), .o(n_580) );
NOR3_Z1 g58940 ( .a(n_1819), .b(n_2095), .c(n_1797), .o(n_2167) );
BUF_X2 newInst_295 ( .a(newNet_294), .o(newNet_295) );
AND2_X1 g58002 ( .a(n_2940), .b(n_2206), .o(n_2969) );
NOR2_Z1 g34206 ( .a(n_4296), .b(n_4178), .o(n_4320) );
NAND2_Z01 g58865 ( .a(n_2155), .b(GPR_14__3_), .o(n_2242) );
AND2_X1 g60797 ( .a(n_177), .b(n_275), .o(n_369) );
INV_X1 g60774 ( .a(n_352), .o(n_351) );
NAND2_Z01 g59409 ( .a(n_1647), .b(n_1163), .o(n_1709) );
INV_Y1 g35383 ( .a(n_3311), .o(n_4685) );
fflopd GPR_reg_11__4_ ( .CK(newNet_1693), .D(n_2948), .Q(GPR_11__4_) );
NAND2_Z01 g35165 ( .a(n_3431), .b(n_4660), .o(n_3464) );
NAND4_Z1 g59670 ( .a(n_1055), .b(n_1290), .c(n_1367), .d(n_1067), .o(n_1458) );
BUF_X2 newInst_997 ( .a(newNet_996), .o(newNet_997) );
AND2_X1 g34485 ( .a(n_4038), .b(n_3255), .o(n_4056) );
XOR2_X1 g34385 ( .a(n_4099), .b(SP_4_), .o(n_4153) );
BUF_X2 newInst_652 ( .a(newNet_83), .o(newNet_652) );
BUF_X2 newInst_4 ( .a(newNet_3), .o(newNet_4) );
BUF_X2 newInst_1830 ( .a(newNet_1829), .o(newNet_1830) );
INV_X1 g61046 ( .a(pX_13_), .o(n_106) );
AND2_X1 g60820 ( .a(n_253), .b(n_4529), .o(n_352) );
NAND4_Z1 g34077 ( .a(n_4255), .b(n_4268), .c(n_4380), .d(n_4127), .o(n_4395) );
NAND4_Z1 g34588 ( .a(n_3843), .b(n_3742), .c(n_3884), .d(n_3741), .o(n_3972) );
NAND2_Z01 g58571 ( .a(n_2483), .b(pX_11_), .o(n_2525) );
NOR2_Z1 g34184 ( .a(n_4324), .b(n_4621), .o(n_4424) );
INV_X1 g61060 ( .a(GPR_18__0_), .o(n_92) );
BUF_X2 newInst_1536 ( .a(newNet_142), .o(newNet_1536) );
NAND2_Z01 g57935 ( .a(n_2972), .b(n_2399), .o(n_3007) );
NAND2_Z01 g34763 ( .a(n_3571), .b(GPR_20__4_), .o(n_3802) );
AND2_X1 g58388 ( .a(n_2657), .b(n_2205), .o(n_2680) );
INV_X1 g60171 ( .a(n_963), .o(n_962) );
NAND2_Z01 g59002 ( .a(n_1912), .b(PC_0_), .o(n_2105) );
NAND4_Z1 g60001 ( .a(n_821), .b(n_897), .c(n_899), .d(n_896), .o(n_1128) );
NAND2_Z01 g59265 ( .a(n_1450), .b(n_1805), .o(n_1845) );
NAND2_Z01 g60241 ( .a(R16_6_), .b(n_14), .o(n_904) );
NAND2_Z01 g60885 ( .a(n_4645), .b(n_4646), .o(n_241) );
NAND2_Z01 g35337 ( .a(pZ_0_), .b(n_3199), .o(n_3333) );
NAND2_Z01 g60232 ( .a(n_598), .b(GPR_15__7_), .o(n_913) );
BUF_X2 newInst_1854 ( .a(newNet_1853), .o(newNet_1854) );
NAND2_Z01 g59434 ( .a(n_1647), .b(n_1397), .o(n_1685) );
fflopd pY_reg_5_ ( .CK(newNet_141), .D(n_3096), .Q(pY_5_) );
NAND4_Z1 g60139 ( .a(n_743), .b(n_712), .c(n_735), .d(n_636), .o(n_993) );
BUF_X2 newInst_512 ( .a(newNet_511), .o(newNet_512) );
AND2_X1 g60579 ( .a(n_68), .b(n_458), .o(n_532) );
NAND2_Z01 g35158 ( .a(n_3432), .b(pmem_d_9), .o(n_4656) );
fflopd PC_reg_9_ ( .CK(newNet_602), .D(n_2533), .Q(PC_9_) );
NAND2_Z01 g58671 ( .a(n_2212), .b(GPR_18__0_), .o(n_2435) );
NAND2_Z01 g58330 ( .a(n_2665), .b(n_2222), .o(n_2735) );
XOR2_X1 final_adder_mux_R16_278_6_g416 ( .a(n_4437), .b(n_4421), .o(final_adder_mux_R16_278_6_n_33) );
NAND2_Z01 g60055 ( .a(n_863), .b(n_153), .o(n_1079) );
NAND4_Z1 g60158 ( .a(n_531), .b(n_533), .c(n_532), .d(n_530), .o(n_977) );
BUF_X2 newInst_1305 ( .a(newNet_1304), .o(newNet_1305) );
NAND2_Z01 g34548 ( .a(n_4537), .b(n_3768), .o(n_4010) );
NAND2_Z01 g60645 ( .a(n_214), .b(n_310), .o(n_573) );
NAND2_Z01 g34620 ( .a(n_3892), .b(n_3481), .o(n_3940) );
NAND2_Z01 g59406 ( .a(io_do_4), .b(n_1649), .o(n_1710) );
NAND2_Z01 g60748 ( .a(SP_14_), .b(n_180), .o(n_394) );
NOR2_Z1 g34896 ( .a(n_3578), .b(n_3265), .o(n_3667) );
NAND2_Z01 g59389 ( .a(n_1669), .b(n_187), .o(n_1726) );
BUF_X2 newInst_1746 ( .a(newNet_1745), .o(newNet_1746) );
fflopd GPR_reg_3__5_ ( .CK(newNet_946), .D(n_3002), .Q(GPR_3__5_) );
NAND3_Z1 g59593 ( .a(n_1339), .b(n_1528), .c(n_321), .o(n_1536) );
XOR2_X1 g35379 ( .a(pY_0_), .b(n_3249), .o(n_3314) );
NOR2_Z1 g59112 ( .a(n_1895), .b(n_1448), .o(n_1997) );
NAND4_Z1 g34228 ( .a(n_4273), .b(n_4201), .c(n_4202), .d(n_4203), .o(n_4303) );
INV_X1 g59309 ( .a(n_1801), .o(n_1802) );
NAND2_Z01 g59075 ( .a(n_1875), .b(n_4566), .o(n_2032) );
NAND2_Z01 g60488 ( .a(n_358), .b(GPR_0__7_), .o(n_658) );
NOR2_Z1 g59355 ( .a(n_19), .b(n_758), .o(n_1758) );
INV_X1 g60780 ( .a(n_323), .o(n_324) );
AND2_X1 g35361 ( .a(n_4489), .b(pmem_d_3), .o(n_4487) );
NOR2_Z1 g34323 ( .a(n_4159), .b(n_3904), .o(n_4210) );
fflopd GPR_reg_22__7_ ( .CK(newNet_1067), .D(n_3154), .Q(GPR_22__7_) );
BUF_X2 newInst_1123 ( .a(newNet_1122), .o(newNet_1123) );
BUF_X2 newInst_688 ( .a(newNet_687), .o(newNet_688) );
NAND2_Z01 g58312 ( .a(n_2681), .b(n_2378), .o(n_2758) );
INV_X1 g61062 ( .a(SP_8_), .o(n_90) );
INV_X1 g60772 ( .a(n_365), .o(n_364) );
NAND2_Z01 g58578 ( .a(n_2481), .b(pX_13_), .o(n_2520) );
NAND2_Z01 g60455 ( .a(n_357), .b(pY_15_), .o(n_691) );
NAND2_Z01 g59219 ( .a(n_1842), .b(n_1241), .o(n_1887) );
AND2_X1 g34453 ( .a(n_4072), .b(n_4645), .o(n_4089) );
NAND2_Z01 g35155 ( .a(n_3450), .b(n_3273), .o(n_3457) );
INV_X1 g61067 ( .a(SP_13_), .o(n_85) );
fflopd io_sel_reg_1_ ( .CK(newNet_338), .D(n_1012), .Q(io_sel_1_) );
BUF_X2 newInst_1043 ( .a(newNet_1042), .o(newNet_1043) );
NOR2_Z1 g34299 ( .a(n_4612), .b(n_3927), .o(n_4235) );
NAND2_Z01 g34756 ( .a(n_3566), .b(GPR_18__4_), .o(n_3809) );
AND3_X1 g59797 ( .a(n_4524), .b(n_1220), .c(n_88), .o(n_1349) );
NAND2_Z01 g59824 ( .a(n_1171), .b(dmem_di_4), .o(n_1300) );
NAND3_Z1 g59033 ( .a(n_965), .b(n_1868), .c(n_963), .o(n_2086) );
NAND2_Z01 g58771 ( .a(n_2202), .b(GPR_5__7_), .o(n_2329) );
NOR3_Z1 g59536 ( .a(n_501), .b(n_1563), .c(n_1010), .o(n_1591) );
BUF_X2 newInst_71 ( .a(newNet_70), .o(newNet_71) );
BUF_X2 newInst_1034 ( .a(newNet_1033), .o(newNet_1034) );
BUF_X2 newInst_1031 ( .a(newNet_1030), .o(newNet_1031) );
BUF_X2 newInst_355 ( .a(newNet_354), .o(newNet_355) );
NOR2_Z1 g34367 ( .a(n_4120), .b(n_3469), .o(n_4168) );
NAND2_Z01 g58046 ( .a(n_2899), .b(n_2418), .o(n_2936) );
BUF_X2 newInst_792 ( .a(newNet_791), .o(newNet_792) );
NAND2_Z01 g59820 ( .a(n_1171), .b(dmem_di_2), .o(n_1304) );
XOR2_X1 g59242 ( .a(n_61), .b(n_6), .o(n_1876) );
BUF_X2 newInst_153 ( .a(newNet_152), .o(newNet_153) );
BUF_X2 newInst_395 ( .a(newNet_394), .o(newNet_395) );
BUF_X2 newInst_453 ( .a(newNet_452), .o(newNet_453) );
fflopd pZ_reg_9_ ( .CK(newNet_36), .D(n_2872), .Q(pZ_9_) );
BUF_X2 newInst_62 ( .a(newNet_61), .o(newNet_62) );
INV_X1 g35037 ( .a(n_3536), .o(n_3535) );
BUF_X2 newInst_617 ( .a(newNet_616), .o(newNet_617) );
fflopd GPR_reg_2__6_ ( .CK(newNet_988), .D(n_3072), .Q(GPR_2__6_) );
NAND2_Z01 g58635 ( .a(n_2360), .b(pY_2_), .o(n_2467) );
NAND2_Z01 g59681 ( .a(n_1377), .b(n_263), .o(n_1452) );
AND2_X1 g60343 ( .a(n_568), .b(n_59), .o(n_860) );
AND2_X1 g35007 ( .a(n_4650), .b(n_3525), .o(n_3569) );
NAND4_Z1 g58828 ( .a(n_1685), .b(n_1787), .c(n_2166), .d(n_2076), .o(n_2279) );
BUF_X2 newInst_596 ( .a(newNet_595), .o(newNet_596) );
NAND2_Z01 g59081 ( .a(n_1871), .b(n_4602), .o(n_2026) );
NOR4_Z1 g35048 ( .a(n_4584), .b(n_4484), .c(n_3479), .d(pmem_d_7), .o(n_4650) );
BUF_X2 newInst_1250 ( .a(newNet_1249), .o(newNet_1250) );
INV_X1 g61027 ( .a(pZ_0_), .o(n_125) );
NOR3_Z1 g59658 ( .a(n_1000), .b(n_1321), .c(n_959), .o(n_1468) );
NOR2_Z1 g35311 ( .a(n_3223), .b(n_3288), .o(n_3365) );
BUF_X2 newInst_1696 ( .a(newNet_1695), .o(newNet_1696) );
NAND2_Z01 g58804 ( .a(n_2197), .b(U_2_), .o(n_2296) );
NAND2_Z01 g58856 ( .a(n_2157), .b(GPR_13__2_), .o(n_2251) );
NAND2_Z01 g60789 ( .a(n_187), .b(n_264), .o(n_318) );
BUF_X2 newInst_331 ( .a(newNet_330), .o(newNet_331) );
NAND2_Z01 g60396 ( .a(n_441), .b(n_438), .o(n_750) );
fflopd GPR_reg_3__2_ ( .CK(newNet_960), .D(n_2747), .Q(GPR_3__2_) );
NAND2_Z01 g60272 ( .a(R16_12_), .b(n_14), .o(n_874) );
AND2_X1 g59773 ( .a(n_1238), .b(n_4664), .o(n_1356) );
INV_X1 g61098 ( .a(io_do_7), .o(n_54) );
NAND2_Z01 g34475 ( .a(n_4045), .b(Rd_0_), .o(n_4066) );
BUF_X2 newInst_629 ( .a(newNet_628), .o(newNet_629) );
BUF_X2 newInst_1070 ( .a(newNet_1069), .o(newNet_1070) );
NAND2_Z01 g60065 ( .a(n_841), .b(io_do_0), .o(n_1069) );
fflopd pX_reg_13_ ( .CK(newNet_257), .D(n_3093), .Q(pX_13_) );
NAND2_Z01 g60440 ( .a(n_368), .b(GPR_15__4_), .o(n_706) );
NAND2_Z02 g58921 ( .a(n_2154), .b(n_1203), .o(n_2201) );
BUF_X2 newInst_183 ( .a(newNet_182), .o(newNet_183) );
NAND2_Z01 g58792 ( .a(n_2199), .b(GPR_0__2_), .o(n_2308) );
NAND2_Z01 g59569 ( .a(n_1467), .b(pmem_d_1), .o(n_1559) );
INV_X1 g59708 ( .a(n_1421), .o(n_1422) );
fflopd C_reg ( .CK(newNet_1827), .D(n_2919), .Q(C) );
NAND4_Z1 g59998 ( .a(n_911), .b(n_912), .c(n_910), .d(n_882), .o(n_1131) );
BUF_X2 newInst_965 ( .a(newNet_964), .o(newNet_965) );
BUF_X2 newInst_383 ( .a(newNet_256), .o(newNet_383) );
XNOR2_X1 g34516 ( .a(n_3960), .b(pZ_6_), .o(n_4029) );
NAND2_Z01 g58733 ( .a(n_2206), .b(GPR_23__7_), .o(n_2374) );
XOR2_X1 g60822 ( .a(io_do_0), .b(io_do_1), .o(n_350) );
NAND3_Z1 g35375 ( .a(n_3258), .b(n_3240), .c(n_3218), .o(n_3315) );
NAND4_Z1 g34230 ( .a(n_4183), .b(n_4184), .c(n_4239), .d(n_4247), .o(n_4301) );
NAND2_Z01 g58689 ( .a(n_2211), .b(GPR_19__5_), .o(n_2417) );
BUF_X2 newInst_1507 ( .a(newNet_1506), .o(newNet_1507) );
INV_X1 g35506 ( .a(PC_6_), .o(n_3221) );
BUF_X2 newInst_308 ( .a(newNet_307), .o(newNet_308) );
AND2_X1 g59764 ( .a(n_1228), .b(pmem_d_1), .o(n_1361) );
NAND2_Z01 g58584 ( .a(n_2465), .b(pY_6_), .o(n_2514) );
BUF_X2 newInst_464 ( .a(newNet_463), .o(newNet_464) );
AND2_X1 g60935 ( .a(n_104), .b(state_3_), .o(n_253) );
NAND2_Z01 g60910 ( .a(PC_4_), .b(pmem_d_4), .o(n_231) );
INV_Z1 g16811 ( .a(GPR_17__0_), .o(n_4409) );
NOR2_Z1 g35116 ( .a(n_3206), .b(pmem_d_7), .o(n_4470) );
INV_X1 g60769 ( .a(n_378), .o(n_377) );
NAND2_Z01 g58683 ( .a(n_2212), .b(GPR_18__7_), .o(n_2423) );
NAND2_Z01 g59220 ( .a(n_1812), .b(io_do_4), .o(n_1886) );
BUF_X2 newInst_1185 ( .a(newNet_1184), .o(newNet_1185) );
NAND2_Z01 g58701 ( .a(n_2210), .b(GPR_1__7_), .o(n_2405) );
fflopd U_reg_13_ ( .CK(newNet_415), .D(n_3092), .Q(U_13_) );
NAND2_Z01 g60023 ( .a(n_822), .b(n_269), .o(n_1120) );
BUF_X2 newInst_35 ( .a(newNet_34), .o(newNet_35) );
NAND2_Z01 g34114 ( .a(n_4333), .b(n_4347), .o(n_4432) );
NAND2_Z01 g58439 ( .a(n_2622), .b(n_2218), .o(n_2654) );
fflopd GPR_reg_4__5_ ( .CK(newNet_900), .D(n_3001), .Q(GPR_4__5_) );
NOR2_Z1 g34849 ( .a(n_3574), .b(n_3239), .o(n_3714) );
INV_X2 g60283 ( .a(n_850), .o(n_849) );
BUF_X2 newInst_1481 ( .a(newNet_1480), .o(newNet_1481) );
NAND2_Z01 g60631 ( .a(n_66), .b(n_335), .o(n_579) );
AND3_X1 g59203 ( .a(n_1486), .b(n_1873), .c(pX_11_), .o(n_1907) );
NOR2_Z1 g59950 ( .a(n_1118), .b(n_969), .o(n_1203) );
NAND2_Z01 g59943 ( .a(n_1039), .b(n_848), .o(n_1206) );
INV_X1 g60543 ( .a(n_564), .o(n_565) );
BUF_X2 newInst_1683 ( .a(newNet_1682), .o(newNet_1683) );
NAND2_Z01 g58639 ( .a(n_2358), .b(pZ_0_), .o(n_2457) );
NAND4_Z1 g60375 ( .a(n_445), .b(n_408), .c(n_444), .d(n_443), .o(n_769) );
NOR2_Z1 g59980 ( .a(n_1043), .b(n_4638), .o(n_1147) );
NOR2_Z1 g60608 ( .a(n_322), .b(n_193), .o(n_515) );
BUF_X2 newInst_862 ( .a(newNet_861), .o(newNet_862) );
XOR2_X1 g60861 ( .a(n_4439), .b(n_4423), .o(n_285) );
NOR2_Z1 g35354 ( .a(n_4560), .b(state_1_), .o(n_3352) );
NAND3_Z3 g59890 ( .a(n_4649), .b(n_1028), .c(n_41), .o(n_1269) );
BUF_X2 newInst_1414 ( .a(newNet_1413), .o(newNet_1414) );
AND2_X1 g35397 ( .a(n_3213), .b(pmem_d_14), .o(n_4684) );
BUF_X2 newInst_1811 ( .a(newNet_1810), .o(newNet_1811) );
BUF_X2 newInst_1323 ( .a(newNet_1322), .o(newNet_1323) );
NAND4_Z1 g58566 ( .a(n_1342), .b(n_2099), .c(n_2447), .d(n_1061), .o(n_2532) );
NAND2_Z01 g58933 ( .a(n_2138), .b(n_849), .o(n_2174) );
NOR2_Z1 g35118 ( .a(n_3203), .b(pmem_d_1), .o(n_4474) );
NAND2_Z01 g59486 ( .a(n_27), .b(n_1534), .o(n_1639) );
BUF_X2 newInst_621 ( .a(newNet_157), .o(newNet_621) );
NOR2_Z1 g34848 ( .a(n_3576), .b(n_4403), .o(n_3715) );
NAND2_Z01 g60475 ( .a(n_370), .b(GPR_20__5_), .o(n_671) );
NAND2_Z01 g58754 ( .a(n_2204), .b(GPR_3__6_), .o(n_2346) );
NAND2_Z02 g58923 ( .a(n_2152), .b(n_1172), .o(n_2199) );
NOR2_Z1 g60589 ( .a(n_378), .b(Z), .o(n_524) );
NAND2_Z01 g60716 ( .a(n_198), .b(GPR_21__1_), .o(n_422) );
BUF_X2 newInst_1403 ( .a(newNet_1402), .o(newNet_1403) );
NOR2_Z1 g34342 ( .a(n_4612), .b(n_3344), .o(n_4192) );
AND2_X1 g58128 ( .a(n_2850), .b(n_2199), .o(n_2884) );
BUF_X2 newInst_564 ( .a(newNet_563), .o(newNet_564) );
BUF_X2 newInst_141 ( .a(newNet_140), .o(newNet_141) );
BUF_X2 newInst_92 ( .a(newNet_91), .o(newNet_92) );
BUF_X2 newInst_57 ( .a(newNet_9), .o(newNet_57) );
BUF_X2 newInst_1428 ( .a(newNet_1427), .o(newNet_1428) );
NAND2_Z01 g58868 ( .a(n_2158), .b(GPR_12__6_), .o(n_2239) );
NAND2_Z01 g60449 ( .a(n_341), .b(pZ_1_), .o(n_697) );
fflopd GPR_reg_1__5_ ( .CK(newNet_1228), .D(n_3008), .Q(GPR_1__5_) );
NAND2_Z01 g60246 ( .a(n_591), .b(GPR_22__7_), .o(n_899) );
BUF_X2 newInst_799 ( .a(newNet_546), .o(newNet_799) );
NAND2_Z01 final_adder_mux_R16_278_6_g432 ( .a(n_4445), .b(n_4429), .o(final_adder_mux_R16_278_6_n_17) );
NAND2_Z01 g60052 ( .a(n_866), .b(pZ_5_), .o(n_1112) );
BUF_X2 newInst_304 ( .a(newNet_303), .o(newNet_304) );
NOR2_Z1 g34284 ( .a(n_4613), .b(n_3255), .o(n_4249) );
BUF_X2 newInst_123 ( .a(newNet_122), .o(newNet_123) );
BUF_X2 newInst_99 ( .a(newNet_9), .o(newNet_99) );
BUF_X2 newInst_898 ( .a(newNet_897), .o(newNet_898) );
NOR2_Z1 g60374 ( .a(n_4556), .b(n_481), .o(n_841) );
NAND2_Z01 g60476 ( .a(n_358), .b(GPR_0__6_), .o(n_670) );
BUF_X2 newInst_1733 ( .a(newNet_1732), .o(newNet_1733) );
AND2_X1 final_adder_mux_R16_278_6_g445 ( .a(n_4438), .b(n_4422), .o(final_adder_mux_R16_278_6_n_4) );
NAND2_Z01 g60894 ( .a(C), .b(pmem_d_12), .o(n_274) );
NAND2_Z01 g60506 ( .a(Rd_2_), .b(n_345), .o(n_640) );
NAND2_Z01 g60909 ( .a(PC_4_), .b(pmem_d_7), .o(n_263) );
NAND2_Z01 g34134 ( .a(n_4317), .b(n_4615), .o(n_4374) );
NAND2_Z01 g34524 ( .a(n_3809), .b(n_3945), .o(n_4020) );
BUF_X2 newInst_977 ( .a(newNet_976), .o(newNet_977) );
NOR3_Z1 g60847 ( .a(n_4647), .b(n_4418), .c(n_241), .o(n_291) );
INV_X1 g59638 ( .a(n_1491), .o(n_1490) );
AND3_X1 g58606 ( .a(n_1997), .b(n_2480), .c(n_1996), .o(n_2505) );
NAND2_Z01 g60112 ( .a(n_779), .b(n_778), .o(n_1014) );
INV_X1 g34356 ( .a(n_4176), .o(n_4175) );
XOR2_X1 g34502 ( .a(n_4649), .b(SP_0_), .o(n_4042) );
AND2_X1 g58409 ( .a(n_2656), .b(n_14), .o(n_2690) );
NAND2_Z01 g58716 ( .a(n_2208), .b(GPR_21__5_), .o(n_2391) );
NOR2_Z1 g59921 ( .a(n_1101), .b(n_4415), .o(n_1194) );
BUF_X2 newInst_578 ( .a(newNet_577), .o(newNet_578) );
AND3_X1 g34065 ( .a(n_3544), .b(n_4397), .c(rst), .o(pmem_ce) );
BUF_X2 newInst_989 ( .a(newNet_955), .o(newNet_989) );
NOR2_Z1 g59729 ( .a(n_161), .b(n_1379), .o(n_1413) );
NAND2_Z01 g34774 ( .a(n_3584), .b(GPR_21__4_), .o(n_3791) );
NAND2_Z01 g34137 ( .a(n_4325), .b(n_4619), .o(n_4371) );
BUF_X2 newInst_1655 ( .a(newNet_1654), .o(newNet_1655) );
NAND2_Z01 g59508 ( .a(n_1564), .b(n_1387), .o(n_1613) );
NAND2_Z01 g59886 ( .a(n_1164), .b(n_61), .o(n_1241) );
NAND2_Z01 g58690 ( .a(n_2211), .b(GPR_19__6_), .o(n_2416) );
NAND2_Z01 g34873 ( .a(n_3573), .b(U_7_), .o(n_3690) );
NAND2_Z01 g58055 ( .a(n_2889), .b(n_2332), .o(n_2927) );
BUF_X2 newInst_1058 ( .a(newNet_1057), .o(newNet_1058) );
NAND3_Z1 g59193 ( .a(n_572), .b(n_1902), .c(n_77), .o(n_1971) );
NAND2_Z01 g34685 ( .a(n_3599), .b(GPR_5__7_), .o(n_3880) );
XOR2_X1 g35074 ( .a(n_3488), .b(pZ_6_), .o(n_3519) );
BUF_X2 newInst_1824 ( .a(newNet_1823), .o(newNet_1824) );
NAND2_Z02 g58928 ( .a(n_2132), .b(n_1979), .o(n_2198) );
INV_X1 g59963 ( .a(n_1159), .o(n_1160) );
NOR2_Z1 g60790 ( .a(V), .b(n_252), .o(n_317) );
BUF_X2 newInst_974 ( .a(newNet_973), .o(newNet_974) );
XOR2_X1 g34661 ( .a(n_3638), .b(n_3319), .o(n_3904) );
NAND2_Z01 g58062 ( .a(n_2908), .b(n_868), .o(n_2941) );
NOR2_Z1 g60307 ( .a(n_599), .b(n_95), .o(n_817) );
NAND2_Z01 g34667 ( .a(n_3613), .b(n_3614), .o(n_3898) );
NAND2_Z01 g59269 ( .a(n_1223), .b(n_6), .o(n_1842) );
NOR2_Z1 g59879 ( .a(n_1160), .b(n_568), .o(n_1248) );
NOR3_Z2 g59494 ( .a(n_1601), .b(n_10), .c(n_595), .o(n_1647) );
BUF_X2 newInst_1102 ( .a(newNet_1101), .o(newNet_1102) );
NAND2_Z01 g57688 ( .a(n_3157), .b(n_2216), .o(n_3178) );
BUF_X2 newInst_723 ( .a(newNet_722), .o(newNet_723) );
NAND2_Z01 g58978 ( .a(n_2085), .b(n_1209), .o(n_2129) );
NAND2_Z01 g57878 ( .a(n_3010), .b(n_2218), .o(n_3061) );
INV_Z1 g16814 ( .a(GPR_8__0_), .o(n_4403) );
INV_X1 g35066 ( .a(n_3520), .o(n_4568) );
NAND2_Z01 g34740 ( .a(n_3584), .b(GPR_21__5_), .o(n_3825) );
NAND2_Z01 g59331 ( .a(n_1736), .b(n_211), .o(n_1782) );
BUF_X2 newInst_1724 ( .a(newNet_1139), .o(newNet_1724) );
NAND2_Z01 g35205 ( .a(n_4533), .b(SP_7_), .o(n_39083_BAR) );
NOR2_Z1 g59751 ( .a(n_1307), .b(n_52), .o(n_1373) );
BUF_X2 newInst_1808 ( .a(newNet_1807), .o(newNet_1808) );
BUF_X2 newInst_196 ( .a(newNet_195), .o(newNet_196) );
NOR2_Z1 g60353 ( .a(n_524), .b(n_507), .o(n_781) );
NOR2_Z1 g34368 ( .a(n_4113), .b(n_3469), .o(n_4167) );
BUF_X2 newInst_1294 ( .a(newNet_1293), .o(newNet_1294) );
NAND2_Z01 g60267 ( .a(n_588), .b(GPR_7__5_), .o(n_879) );
NAND2_Z01 g34533 ( .a(n_3936), .b(n_3539), .o(n_4563) );
NAND2_Z01 g58355 ( .a(n_2655), .b(n_25), .o(n_2716) );
NAND2_Z01 g34625 ( .a(n_3769), .b(pZ_5_), .o(n_3935) );
INV_X1 g35477 ( .a(pY_5_), .o(n_3247) );
NOR2_Z1 g59014 ( .a(n_1921), .b(n_63), .o(n_2094) );
AND3_X1 g34498 ( .a(n_3964), .b(n_4003), .c(n_4014), .o(n_4046) );
AND2_X1 g58506 ( .a(n_2567), .b(n_2210), .o(n_2591) );
NAND2_Z01 g59429 ( .a(n_1647), .b(n_478), .o(n_1690) );
NAND3_Z1 g59246 ( .a(n_1767), .b(n_1833), .c(n_4666), .o(n_1864) );
BUF_X2 newInst_1622 ( .a(newNet_590), .o(newNet_1622) );
BUF_X2 newInst_1266 ( .a(newNet_1265), .o(newNet_1266) );
NAND2_Z01 g58998 ( .a(n_1975), .b(n_4574), .o(n_2109) );
NAND2_Z01 g35226 ( .a(n_3359), .b(n_3220), .o(n_4634) );
XOR2_X1 g60165 ( .a(n_612), .b(io_do_4), .o(n_1024) );
BUF_X2 newInst_1469 ( .a(newNet_1468), .o(newNet_1469) );
BUF_X2 newInst_1849 ( .a(newNet_1848), .o(newNet_1849) );
NOR2_Z1 g34276 ( .a(n_4613), .b(n_3235), .o(n_4257) );
INV_X1 g61058 ( .a(pZ_8_), .o(n_94) );
NAND4_Z2 g35183 ( .a(n_3342), .b(n_3380), .c(n_3374), .d(n_3388), .o(n_4622) );
XOR2_X1 g35201 ( .a(n_3324), .b(n_3301), .o(n_3453) );
NAND2_Z01 g34264 ( .a(n_4176), .b(pX_10_), .o(n_4269) );
NAND2_Z01 g34530 ( .a(n_3662), .b(n_3940), .o(n_4015) );
NAND2_Z01 g60226 ( .a(n_588), .b(GPR_7__0_), .o(n_919) );
AND2_X1 g60836 ( .a(n_175), .b(n_272), .o(n_345) );
NAND2_Z01 g59274 ( .a(io_do_2), .b(n_1766), .o(n_1839) );
BUF_X2 newInst_1360 ( .a(newNet_1359), .o(newNet_1360) );
NAND3_Z1 g60646 ( .a(n_4622), .b(n_186), .c(pmem_d_2), .o(n_494) );
NAND2_Z01 g34807 ( .a(n_3581), .b(GPR_16__2_), .o(n_3756) );
NAND2_Z01 g35003 ( .a(n_3509), .b(n_3552), .o(n_3576) );
BUF_X2 newInst_487 ( .a(newNet_486), .o(newNet_487) );
INV_X1 g59907 ( .a(io_sel_1_), .o(n_1224) );
NAND2_Z01 g35084 ( .a(n_3481), .b(n_3469), .o(n_3510) );
NAND2_Z01 g60722 ( .a(U_1_), .b(n_249), .o(n_416) );
NAND2_Z01 g58317 ( .a(n_2678), .b(n_2351), .o(n_2748) );
XOR2_X1 g60010 ( .a(n_861), .b(io_do_5), .o(n_1155) );
BUF_X2 newInst_1010 ( .a(newNet_1009), .o(newNet_1010) );
INV_X1 g60873 ( .a(n_255), .o(n_254) );
NAND2_Z01 g57706 ( .a(n_3135), .b(n_2433), .o(n_3163) );
BUF_X2 newInst_384 ( .a(newNet_383), .o(newNet_384) );
BUF_X2 newInst_1364 ( .a(newNet_1363), .o(newNet_1364) );
fflopd GPR_reg_2__7_ ( .CK(newNet_983), .D(n_3153), .Q(GPR_2__7_) );
NAND2_Z01 g60034 ( .a(n_4600), .b(n_856), .o(n_1096) );
NOR2_Z1 g34422 ( .a(n_4610), .b(n_3499), .o(n_4115) );
fflopd GPR_reg_3__4_ ( .CK(newNet_948), .D(n_2929), .Q(GPR_3__4_) );
NOR2_Z1 g59566 ( .a(n_1486), .b(n_114), .o(n_1570) );
AND2_X1 g58379 ( .a(n_2657), .b(n_2209), .o(n_2692) );
BUF_X2 newInst_1286 ( .a(newNet_451), .o(newNet_1286) );
BUF_X2 newInst_104 ( .a(newNet_103), .o(newNet_104) );
NAND2_Z01 g58558 ( .a(n_2504), .b(pY_14_), .o(n_2540) );
NAND4_Z1 g59414 ( .a(n_877), .b(n_902), .c(n_1617), .d(n_876), .o(n_1706) );
BUF_X2 newInst_177 ( .a(newNet_141), .o(newNet_177) );
BUF_X2 newInst_1841 ( .a(newNet_1840), .o(newNet_1841) );
AND3_X1 g58831 ( .a(n_4644), .b(n_2143), .c(n_4615), .o(n_2276) );
AND2_X1 g34224 ( .a(n_4282), .b(n_4178), .o(n_4306) );
NAND2_Z01 g58699 ( .a(n_2210), .b(GPR_1__6_), .o(n_2407) );
INV_X1 g35505 ( .a(pY_10_), .o(n_3222) );
NAND2_Z01 g57846 ( .a(n_872), .b(n_3056), .o(n_3080) );
INV_X1 g60954 ( .a(n_178), .o(n_177) );
BUF_X2 newInst_981 ( .a(newNet_980), .o(newNet_981) );
XOR2_X1 g60867 ( .a(n_4440), .b(n_4424), .o(n_281) );
NAND2_Z01 g34681 ( .a(n_3599), .b(GPR_5__2_), .o(n_3884) );
INV_X1 drc_bufs61245 ( .a(n_3), .o(n_4) );
INV_X2 g61117 ( .a(pmem_d_1), .o(n_35) );
NAND3_Z1 g60816 ( .a(n_4518), .b(n_4517), .c(n_88), .o(n_354) );
NAND3_Z1 g60101 ( .a(n_697), .b(n_696), .c(n_698), .o(n_1019) );
BUF_X2 newInst_1612 ( .a(newNet_1611), .o(newNet_1612) );
BUF_X2 newInst_124 ( .a(newNet_123), .o(newNet_124) );
BUF_X2 newInst_719 ( .a(newNet_718), .o(newNet_719) );
NOR2_Z1 g35245 ( .a(n_3347), .b(n_4683), .o(n_4666) );
BUF_X2 newInst_1524 ( .a(newNet_1523), .o(newNet_1524) );
NAND2_Z01 g34117 ( .a(n_4330), .b(n_4344), .o(n_4435) );
NOR2_Z1 g60799 ( .a(n_199), .b(n_258), .o(n_368) );
INV_X1 g35127 ( .a(n_3482), .o(n_3481) );
BUF_X2 newInst_1567 ( .a(newNet_1566), .o(newNet_1567) );
NAND2_Z01 g60682 ( .a(GPR_7__2_), .b(n_183), .o(n_455) );
INV_X1 g61076 ( .a(pZ_13_), .o(n_76) );
NAND2_Z01 g60611 ( .a(n_325), .b(n_169), .o(n_512) );
BUF_X2 newInst_237 ( .a(newNet_173), .o(newNet_237) );
BUF_X2 newInst_137 ( .a(newNet_136), .o(newNet_137) );
INV_X1 g61037 ( .a(pX_2_), .o(n_115) );
NOR2_Z1 g34349 ( .a(n_16064_BAR), .b(pY_0_), .o(n_4185) );
BUF_X2 newInst_956 ( .a(newNet_955), .o(newNet_956) );
BUF_X2 newInst_1204 ( .a(newNet_1203), .o(newNet_1204) );
BUF_X2 newInst_899 ( .a(newNet_898), .o(newNet_899) );
AND2_X1 g57734 ( .a(n_3115), .b(n_2155), .o(n_3138) );
BUF_X2 newInst_277 ( .a(newNet_276), .o(newNet_277) );
INV_Z1 g16798 ( .a(n_4583), .o(io_we) );
BUF_X2 newInst_1535 ( .a(newNet_1534), .o(newNet_1535) );
BUF_X2 newInst_1637 ( .a(newNet_1636), .o(newNet_1637) );
NAND2_Z01 g34837 ( .a(n_3566), .b(GPR_18__1_), .o(n_3726) );
NOR2_Z1 g58950 ( .a(n_2089), .b(n_964), .o(n_2161) );
NAND2_Z01 g60073 ( .a(n_841), .b(io_do_5), .o(n_1061) );
NAND2_Z01 g35394 ( .a(SP_2_), .b(SP_3_), .o(n_4536) );
NAND2_Z01 g59473 ( .a(n_1603), .b(n_219), .o(n_1651) );
NAND2_Z01 g34646 ( .a(n_3768), .b(n_4541), .o(n_3914) );
fflopd GPR_reg_7__0_ ( .CK(newNet_785), .D(n_2618), .Q(GPR_7__0_) );
NAND2_Z01 g60300 ( .a(n_577), .b(pZ_15_), .o(n_824) );
NAND2_Z01 g34329 ( .a(n_4165), .b(n_4538), .o(n_4205) );
BUF_X2 newInst_739 ( .a(newNet_738), .o(newNet_739) );
NAND2_Z01 g58100 ( .a(n_2852), .b(n_2196), .o(n_2913) );
NAND3_Z1 g59975 ( .a(n_562), .b(n_1030), .c(n_654), .o(n_1150) );
BUF_X2 newInst_1382 ( .a(newNet_1381), .o(newNet_1382) );
BUF_X2 newInst_1039 ( .a(newNet_1038), .o(newNet_1039) );
NAND4_Z1 g34573 ( .a(n_3820), .b(n_3824), .c(n_3823), .d(n_3821), .o(n_3987) );
NAND4_Z1 g58133 ( .a(n_1916), .b(n_2497), .c(n_2827), .d(n_2041), .o(n_2880) );
NAND2_Z01 g35341 ( .a(n_3287), .b(pmem_d_12), .o(n_3330) );
NOR2_Z1 g59688 ( .a(n_1348), .b(n_76), .o(n_1448) );
NAND2_Z01 g34427 ( .a(n_4098), .b(n_4607), .o(n_4110) );
NOR2_Z1 g59356 ( .a(n_1701), .b(n_1226), .o(n_1757) );
AND2_X1 g58374 ( .a(n_2656), .b(n_2212), .o(n_2697) );
NAND2_Z01 g59586 ( .a(n_1268), .b(n_1484), .o(n_1542) );
INV_X1 g61051 ( .a(PC_7_), .o(n_101) );
NAND2_Z01 g58810 ( .a(n_2195), .b(U_8_), .o(n_2290) );
NAND2_Z01 g60039 ( .a(n_856), .b(n_4608), .o(n_1091) );
BUF_X2 newInst_781 ( .a(newNet_780), .o(newNet_781) );
NAND2_Z01 g59395 ( .a(n_1648), .b(dmem_di_5), .o(n_1720) );
INV_X1 g60088 ( .a(n_1047), .o(n_1046) );
AND2_X1 g59713 ( .a(n_1385), .b(pmem_d_6), .o(n_1411) );
NAND2_Z01 g59001 ( .a(n_2007), .b(n_1245), .o(n_2106) );
BUF_X1 drc_bufs61251 ( .a(n_2568), .o(n_0) );
INV_X1 drc_bufs35583 ( .a(n_4647), .o(n_3207) );
AND2_X1 g57899 ( .a(n_3009), .b(n_2206), .o(n_3039) );
BUF_X2 newInst_696 ( .a(newNet_695), .o(newNet_696) );
NAND4_Z1 g59250 ( .a(n_1719), .b(n_1709), .c(n_1789), .d(n_1086), .o(n_1862) );
BUF_X2 newInst_344 ( .a(newNet_343), .o(newNet_344) );
INV_X1 g34976 ( .a(n_3583), .o(n_3584) );
NAND2_Z01 g57880 ( .a(n_3011), .b(n_2215), .o(n_3059) );
BUF_X2 newInst_1587 ( .a(newNet_1586), .o(newNet_1587) );
NAND2_Z01 g34810 ( .a(n_3636), .b(GPR_10__2_), .o(n_3753) );
NAND2_Z01 g58975 ( .a(n_2084), .b(n_1213), .o(n_2132) );
BUF_X2 newInst_919 ( .a(newNet_918), .o(newNet_919) );
AND2_X1 g60081 ( .a(n_848), .b(n_35), .o(n_1054) );
NOR2_Z1 g34988 ( .a(n_3550), .b(n_3482), .o(n_3594) );
BUF_X2 newInst_1073 ( .a(newNet_1072), .o(newNet_1073) );
NAND3_Z1 g60804 ( .a(n_4519), .b(n_4520), .c(n_110), .o(n_363) );
NAND2_Z01 g60570 ( .a(n_341), .b(pY_6_), .o(n_540) );
AND2_X1 g58012 ( .a(n_2940), .b(n_2199), .o(n_2960) );
fflopd GPR_reg_6__6_ ( .CK(newNet_798), .D(n_3068), .Q(GPR_6__6_) );
AND3_X1 g58982 ( .a(n_120), .b(n_1983), .c(pY_9_), .o(n_2125) );
NAND3_Z1 g60119 ( .a(n_4532), .b(n_857), .c(n_73), .o(n_1008) );
BUF_X2 newInst_1729 ( .a(newNet_1649), .o(newNet_1729) );
BUF_X2 newInst_1236 ( .a(newNet_1235), .o(newNet_1236) );
AND2_X1 g57743 ( .a(n_3115), .b(n_2208), .o(n_3128) );
BUF_X2 newInst_597 ( .a(newNet_596), .o(newNet_597) );
AND2_X1 g35298 ( .a(n_3253), .b(n_3298), .o(n_3377) );
AND2_X1 g57744 ( .a(n_3115), .b(n_2207), .o(n_3127) );
NAND2_Z01 g34291 ( .a(n_4164), .b(pmem_d_3), .o(n_4242) );
BUF_X2 newInst_1035 ( .a(newNet_1034), .o(newNet_1035) );
BUF_X2 newInst_912 ( .a(newNet_911), .o(newNet_912) );
BUF_X2 newInst_84 ( .a(newNet_83), .o(newNet_84) );
NAND2_Z01 g60689 ( .a(n_198), .b(GPR_16__1_), .o(n_449) );
AND2_X1 g58254 ( .a(n_2752), .b(n_2155), .o(n_2813) );
BUF_X2 newInst_414 ( .a(newNet_413), .o(newNet_414) );
NAND2_Z01 g34878 ( .a(n_3567), .b(GPR_6__7_), .o(n_3685) );
NOR2_Z1 g35264 ( .a(n_4535), .b(n_3242), .o(n_4533) );
fflopd SP_reg_8_ ( .CK(newNet_474), .D(n_1576), .Q(SP_8_) );
INV_X1 g35389 ( .a(n_4668), .o(n_3302) );
NAND2_Z01 g60886 ( .a(n_34), .b(n_4451), .o(n_240) );
INV_X2 newInst_610 ( .a(newNet_562), .o(newNet_610) );
BUF_X2 newInst_905 ( .a(newNet_904), .o(newNet_905) );
NAND2_Z01 g59835 ( .a(n_1206), .b(io_do_5), .o(n_1290) );
NAND2_Z01 g34716 ( .a(n_3197), .b(GPR_23__6_), .o(n_3849) );
NAND2_Z01 g59523 ( .a(n_1548), .b(n_41), .o(n_1619) );
AND3_X1 g35047 ( .a(n_4655), .b(n_4654), .c(n_3449), .o(n_3530) );
NOR2_X2 g60653 ( .a(n_4556), .b(n_461), .o(n_571) );
NAND2_Z02 g58909 ( .a(n_2161), .b(n_1204), .o(n_2213) );
AND2_X1 g35089 ( .a(n_3480), .b(pY_6_), .o(n_3506) );
INV_X1 g35388 ( .a(n_4514), .o(n_3305) );
BUF_X2 newInst_852 ( .a(newNet_851), .o(newNet_852) );
NOR2_Z1 g60621 ( .a(n_344), .b(H), .o(n_507) );
fflopd GPR_reg_23__4_ ( .CK(newNet_1041), .D(n_2931), .Q(GPR_23__4_) );
XNOR2_X1 g59738 ( .a(n_1283), .b(pmem_d_10), .o(n_1392) );
NAND2_Z01 g58772 ( .a(n_2201), .b(GPR_6__0_), .o(n_2328) );
NOR2_Z1 g58648 ( .a(n_2355), .b(n_1935), .o(n_2459) );
BUF_X2 newInst_1764 ( .a(newNet_889), .o(newNet_1764) );
BUF_X2 newInst_1689 ( .a(newNet_651), .o(newNet_1689) );
BUF_X2 newInst_640 ( .a(newNet_639), .o(newNet_640) );
NAND2_Z01 final_adder_mux_R16_278_6_g377 ( .a(final_adder_mux_R16_278_6_n_71), .b(final_adder_mux_R16_278_6_n_12), .o(final_adder_mux_R16_278_6_n_72) );
NOR2_Z1 g34183 ( .a(n_4324), .b(n_4619), .o(n_4423) );
INV_X1 g35092 ( .a(n_4592), .o(n_3500) );
NAND2_Z01 g60544 ( .a(n_342), .b(GPR_17__7_), .o(n_562) );
BUF_X2 newInst_1657 ( .a(newNet_582), .o(newNet_1657) );
AND2_X1 g58819 ( .a(n_2218), .b(n_1978), .o(n_2357) );
NAND2_Z01 g58875 ( .a(n_2153), .b(GPR_8__1_), .o(n_2232) );
NOR2_Z1 g59485 ( .a(n_1619), .b(n_1393), .o(n_1640) );
BUF_X2 newInst_14 ( .a(newNet_13), .o(newNet_14) );
NAND4_Z1 g60663 ( .a(n_62), .b(n_4653), .c(n_4412), .d(pmem_d_1), .o(n_483) );
BUF_X2 newInst_265 ( .a(newNet_172), .o(newNet_265) );
INV_X1 g61097 ( .a(io_do_5), .o(n_55) );
NAND2_Z01 g58838 ( .a(n_2159), .b(GPR_10__4_), .o(n_2269) );
BUF_X2 newInst_1299 ( .a(newNet_1298), .o(newNet_1299) );
NAND4_Z1 g34567 ( .a(n_3859), .b(n_3860), .c(n_3857), .d(n_3858), .o(n_3993) );
fflopd GPR_reg_1__2_ ( .CK(newNet_1252), .D(n_2766), .Q(GPR_1__2_) );
NOR2_Z1 g34907 ( .a(n_3562), .b(n_3245), .o(n_3656) );
NOR2_Z1 g60929 ( .a(n_4685), .b(n_45), .o(n_216) );
NAND2_Z01 g58473 ( .a(n_2344), .b(n_2583), .o(n_2623) );
NAND2_Z01 g59613 ( .a(n_1414), .b(io_di_1), .o(n_1514) );
BUF_X2 newInst_1270 ( .a(newNet_89), .o(newNet_1270) );
BUF_X2 newInst_215 ( .a(newNet_32), .o(newNet_215) );
NAND2_Z01 g60906 ( .a(PC_9_), .b(pmem_d_9), .o(n_265) );
NAND3_Z1 g58610 ( .a(n_2147), .b(n_2285), .c(n_849), .o(n_2488) );
AND2_X1 g60109 ( .a(n_4556), .b(n_842), .o(n_1043) );
NAND2_Z01 g34613 ( .a(n_3899), .b(n_3483), .o(n_3947) );
NAND2_Z01 g57937 ( .a(n_2970), .b(n_2383), .o(n_3005) );
NAND2_Z01 g60046 ( .a(n_764), .b(n_364), .o(n_1084) );
AND2_X1 g60736 ( .a(n_97), .b(n_204), .o(n_403) );
BUF_X2 newInst_1802 ( .a(newNet_1325), .o(newNet_1802) );
NAND2_Z01 g59087 ( .a(n_1871), .b(n_4600), .o(n_2020) );
NAND2_Z01 g59092 ( .a(n_1900), .b(pmem_d_11), .o(n_2015) );
NOR2_Z1 g59765 ( .a(n_1311), .b(rst), .o(n_1387) );
BUF_X2 newInst_1005 ( .a(newNet_1004), .o(newNet_1005) );
INV_X1 g61085 ( .a(n_4614), .o(n_67) );
BUF_X2 newInst_746 ( .a(newNet_745), .o(newNet_746) );
NAND2_Z01 g58766 ( .a(n_2202), .b(GPR_5__2_), .o(n_2334) );
NAND2_Z01 g34741 ( .a(n_3586), .b(GPR_9__5_), .o(n_3824) );
fflopd GPR_reg_21__0_ ( .CK(newNet_1166), .D(n_2628), .Q(GPR_21__0_) );
NOR2_Z1 g60596 ( .a(n_338), .b(n_172), .o(n_521) );
NOR2_Z1 g34279 ( .a(n_4613), .b(n_3210), .o(n_4254) );
NAND2_Z01 g60900 ( .a(PC_0_), .b(pmem_d_0), .o(n_270) );
NAND2_Z01 g60183 ( .a(n_623), .b(n_725), .o(n_957) );
NAND2_Z01 g35120 ( .a(n_3464), .b(n_3330), .o(n_4661) );
INV_X1 drc_bufs61132 ( .a(n_16), .o(n_17) );
BUF_X2 newInst_824 ( .a(newNet_823), .o(newNet_824) );
NAND2_Z01 g59579 ( .a(n_1490), .b(n_573), .o(n_1552) );
AND3_X1 g59986 ( .a(n_333), .b(n_801), .c(n_119), .o(n_1158) );
NAND2_Z01 g60519 ( .a(n_371), .b(GPR_23__1_), .o(n_627) );
XOR2_X1 g35019 ( .a(n_3528), .b(n_3329), .o(n_3557) );
BUF_X2 newInst_583 ( .a(newNet_582), .o(newNet_583) );
NAND3_Z1 g35250 ( .a(n_4668), .b(n_3200), .c(pmem_d_13), .o(n_4558) );
NOR3_Z1 g58523 ( .a(n_333), .b(n_2554), .c(n_175), .o(n_2574) );
BUF_X1 mybuffer4 ( .o(io_a_4), .a(pmem_d_9) );
NAND2_Z01 g58645 ( .a(n_2359), .b(n_2011), .o(n_2462) );
BUF_X2 newInst_419 ( .a(newNet_418), .o(newNet_419) );
NOR2_Z1 g59819 ( .a(n_1219), .b(n_56), .o(n_1305) );
XOR2_X1 final_adder_mux_R16_278_6_g364 ( .a(final_adder_mux_R16_278_6_n_83), .b(final_adder_mux_R16_278_6_n_33), .o(R16_14_) );
BUF_X2 newInst_370 ( .a(newNet_369), .o(newNet_370) );
NAND2_Z01 g58841 ( .a(n_2159), .b(GPR_10__7_), .o(n_2266) );
BUF_X2 newInst_113 ( .a(newNet_112), .o(newNet_113) );
BUF_X2 newInst_1164 ( .a(newNet_1163), .o(newNet_1164) );
BUF_X2 newInst_1739 ( .a(newNet_1738), .o(newNet_1739) );
BUF_X2 newInst_39 ( .a(newNet_38), .o(newNet_39) );
BUF_X2 newInst_1477 ( .a(newNet_1476), .o(newNet_1477) );
AND2_X1 g59857 ( .a(n_1208), .b(pmem_d_4), .o(n_1307) );
NAND2_Z01 g58099 ( .a(n_2851), .b(n_2216), .o(n_2914) );
BUF_X2 newInst_548 ( .a(newNet_547), .o(newNet_548) );
AND2_X1 g35293 ( .a(n_3241), .b(n_3298), .o(n_3382) );
fflopd pZ_reg_3_ ( .CK(newNet_77), .D(n_2954), .Q(pZ_3_) );
NAND2_Z01 g59602 ( .a(n_1413), .b(io_sp_7_), .o(n_1524) );
BUF_X2 newInst_1277 ( .a(newNet_1276), .o(newNet_1277) );
BUF_X2 newInst_1337 ( .a(newNet_637), .o(newNet_1337) );
BUF_X2 newInst_426 ( .a(newNet_425), .o(newNet_426) );
INV_X1 g59209 ( .a(n_1897), .o(n_1898) );
BUF_X2 newInst_772 ( .a(newNet_629), .o(newNet_772) );
NOR2_Z1 g60702 ( .a(n_4416), .b(n_159), .o(n_436) );
BUF_X2 newInst_205 ( .a(newNet_204), .o(newNet_205) );
XOR2_X1 g58989 ( .a(n_1984), .b(pmem_d_11), .o(n_2138) );
NAND2_Z01 g35398 ( .a(state_0_), .b(state_1_), .o(n_3310) );
BUF_X2 newInst_8 ( .a(newNet_7), .o(newNet_8) );
NAND2_Z01 g59148 ( .a(n_1896), .b(n_971), .o(n_1951) );
INV_X1 g59346 ( .a(n_1766), .o(n_1765) );
NAND2_Z01 g34639 ( .a(n_3769), .b(pZ_2_), .o(n_3921) );
INV_X1 g59417 ( .a(n_1703), .o(n_1704) );
fflopd GPR_reg_19__2_ ( .CK(newNet_1309), .D(n_2768), .Q(GPR_19__2_) );
XOR2_X1 g34928 ( .a(n_3547), .b(pX_9_), .o(n_3766) );
fflopd pX_reg_6_ ( .CK(newNet_213), .D(n_3114), .Q(pX_6_) );
BUF_X2 newInst_151 ( .a(newNet_150), .o(newNet_151) );
BUF_X2 newInst_537 ( .a(newNet_536), .o(newNet_537) );
NAND2_Z01 g34785 ( .a(n_3566), .b(GPR_18__3_), .o(n_3780) );
NAND2_Z01 g57801 ( .a(n_3079), .b(n_2218), .o(n_3106) );
BUF_X2 newInst_163 ( .a(newNet_162), .o(newNet_163) );
NAND2_Z01 g34401 ( .a(n_3208), .b(pZ_3_), .o(n_4137) );
NOR2_Z1 g35355 ( .a(n_4637), .b(state_2_), .o(n_3351) );
NAND3_Z1 g34555 ( .a(n_3716), .b(n_3718), .c(n_3717), .o(n_4004) );
NAND2_Z01 g57805 ( .a(n_3079), .b(n_2216), .o(n_3102) );
AND2_X1 g58003 ( .a(n_2940), .b(n_2205), .o(n_2968) );
BUF_X2 newInst_810 ( .a(newNet_809), .o(newNet_810) );
NAND2_Z01 g59625 ( .a(n_17), .b(H), .o(n_1502) );
NAND2_Z01 g34955 ( .a(n_3536), .b(GPR_21__2_), .o(n_3607) );
BUF_X2 newInst_390 ( .a(newNet_389), .o(newNet_390) );
AND3_X1 g59039 ( .a(n_4514), .b(n_1982), .c(pZ_10_), .o(n_2069) );
NOR2_Z1 g34374 ( .a(n_4103), .b(n_4088), .o(n_4156) );
AND2_X1 g58402 ( .a(n_2656), .b(n_2153), .o(n_2666) );
NAND2_Z01 g58894 ( .a(n_2134), .b(n_1784), .o(n_2188) );
BUF_X2 newInst_258 ( .a(newNet_172), .o(newNet_258) );
NAND3_Z1 g60125 ( .a(n_36), .b(n_605), .c(pmem_d_11), .o(n_1039) );
BUF_X2 newInst_1510 ( .a(newNet_1509), .o(newNet_1510) );
BUF_X2 newInst_448 ( .a(newNet_447), .o(newNet_448) );
fflopd GPR_reg_18__2_ ( .CK(newNet_1358), .D(n_2771), .Q(GPR_18__2_) );
INV_X1 g35483 ( .a(pX_11_), .o(n_3241) );
BUF_X2 newInst_1580 ( .a(newNet_1579), .o(newNet_1580) );
NAND2_Z01 g60896 ( .a(state_0_), .b(state_3_), .o(n_272) );
NAND4_Z1 g58532 ( .a(n_1179), .b(n_2133), .c(n_2491), .d(n_1256), .o(n_2565) );
INV_X1 g34796 ( .a(n_3767), .o(n_4601) );
BUF_X2 newInst_1674 ( .a(newNet_1673), .o(newNet_1674) );
AND2_X1 g58514 ( .a(n_2567), .b(n_2202), .o(n_2582) );
NAND3_Z1 g59347 ( .a(n_1093), .b(n_1658), .c(n_800), .o(n_1773) );
NAND2_Z01 g34322 ( .a(n_4166), .b(n_4551), .o(n_4211) );
BUF_X2 newInst_1215 ( .a(newNet_246), .o(newNet_1215) );
BUF_X2 newInst_350 ( .a(newNet_349), .o(newNet_350) );
AND4_X1 g59850 ( .a(state_2_), .b(n_862), .c(n_150), .d(state_3_), .o(n_1310) );
NAND2_Z01 g59699 ( .a(io_do_4), .b(n_1353), .o(n_1431) );
NAND2_Z01 g34151 ( .a(n_4317), .b(n_4682), .o(n_4357) );
NAND2_Z01 g34144 ( .a(n_4317), .b(n_4623), .o(n_4364) );
NAND2_Z01 g35449 ( .a(n_3232), .b(n_3225), .o(n_3269) );
NAND2_Z01 g58463 ( .a(n_2431), .b(n_2595), .o(n_2633) );
BUF_X2 newInst_286 ( .a(newNet_285), .o(newNet_286) );
NAND2_Z01 g35442 ( .a(n_3265), .b(n_3236), .o(n_3283) );
NAND4_Z1 g58346 ( .a(n_2077), .b(n_2511), .c(n_2651), .d(n_2035), .o(n_2724) );
NAND2_Z01 g59846 ( .a(n_1157), .b(n_1032), .o(n_1280) );
INV_X1 drc_bufs61220 ( .a(n_9), .o(n_10) );
AND2_X1 g60064 ( .a(n_848), .b(n_65), .o(n_1070) );
NAND2_Z01 final_adder_mux_R16_278_6_g395 ( .a(final_adder_mux_R16_278_6_n_53), .b(final_adder_mux_R16_278_6_n_0), .o(final_adder_mux_R16_278_6_n_54) );
NAND2_Z01 g60417 ( .a(n_370), .b(GPR_20__7_), .o(n_729) );
BUF_X2 newInst_1705 ( .a(newNet_1704), .o(newNet_1705) );
AND2_X1 g57989 ( .a(n_2940), .b(n_2139), .o(n_2982) );
BUF_X2 newInst_223 ( .a(newNet_222), .o(newNet_223) );
BUF_X2 newInst_1519 ( .a(newNet_1518), .o(newNet_1519) );
XNOR2_X1 g34933 ( .a(n_3537), .b(pY_12_), .o(n_4585) );
NAND2_Z01 g59104 ( .a(n_1894), .b(n_615), .o(n_2005) );
fflopd GPR_reg_6__7_ ( .CK(newNet_794), .D(n_3148), .Q(GPR_6__7_) );
NAND3_Z1 g59724 ( .a(n_1095), .b(n_1246), .c(n_535), .o(n_1403) );
BUF_X2 newInst_949 ( .a(newNet_744), .o(newNet_949) );
BUF_X2 newInst_801 ( .a(newNet_800), .o(newNet_801) );
BUF_X2 newInst_244 ( .a(newNet_243), .o(newNet_244) );
NAND2_Z01 g60691 ( .a(n_200), .b(GPR_13__1_), .o(n_447) );
AND2_X1 g58112 ( .a(n_2850), .b(n_2212), .o(n_2900) );
NOR2_Z1 g59152 ( .a(n_1873), .b(n_1665), .o(n_1947) );
NAND2_Z01 g60467 ( .a(n_370), .b(GPR_20__0_), .o(n_679) );
fflopd pX_reg_1_ ( .CK(newNet_247), .D(n_2882), .Q(pX_1_) );
INV_X1 g58748 ( .a(n_2352), .o(n_2353) );
BUF_X2 newInst_1431 ( .a(newNet_1430), .o(newNet_1431) );
NAND2_Z01 g58440 ( .a(n_2621), .b(n_2217), .o(n_2653) );
NAND2_Z01 g58480 ( .a(n_2588), .b(n_947), .o(n_2622) );
BUF_X2 newInst_1827 ( .a(newNet_1826), .o(newNet_1827) );
NOR2_Z1 g59870 ( .a(n_760), .b(n_1166), .o(n_1257) );
NAND2_Z01 g34179 ( .a(n_4325), .b(n_4474), .o(n_4337) );
NAND2_Z01 g34883 ( .a(n_3630), .b(pX_12_), .o(n_3680) );
BUF_X2 newInst_829 ( .a(newNet_828), .o(newNet_829) );
NAND2_Z01 g58583 ( .a(n_2464), .b(pY_5_), .o(n_2515) );
BUF_X2 newInst_366 ( .a(newNet_110), .o(newNet_366) );
NAND2_Z01 g34824 ( .a(n_3629), .b(GPR_3__2_), .o(n_3739) );
NOR2_Z1 g34991 ( .a(n_3548), .b(n_3484), .o(n_3591) );
INV_X1 drc_bufs35532 ( .a(n_4624), .o(n_3203) );
AND2_X1 g59133 ( .a(n_1873), .b(n_4573), .o(n_1965) );
AND2_X1 g60984 ( .a(n_4616), .b(pmem_d_7), .o(n_145) );
NAND2_Z01 g35057 ( .a(n_3501), .b(n_4530), .o(n_3526) );
NAND2_Z01 g57718 ( .a(n_3122), .b(n_2329), .o(n_3149) );
NAND2_Z01 g59842 ( .a(n_1168), .b(n_1182), .o(n_1284) );
BUF_X2 newInst_1130 ( .a(newNet_1129), .o(newNet_1130) );
BUF_X2 newInst_450 ( .a(newNet_449), .o(newNet_450) );
BUF_X2 newInst_1552 ( .a(newNet_1551), .o(newNet_1552) );
BUF_X2 newInst_815 ( .a(newNet_305), .o(newNet_815) );
fflopd GPR_Rd_r_reg_3_ ( .CK(newNet_1856), .D(io_do_3), .Q(GPR_Rd_r_3_) );
NAND2_Z01 g57660 ( .a(n_3171), .b(n_1771), .o(n_3182) );
fflopd SP_reg_3_ ( .CK(newNet_503), .D(n_1673), .Q(SP_3_) );
NAND2_Z01 g60415 ( .a(n_329), .b(n_4435), .o(n_731) );
NAND2_Z01 g60275 ( .a(n_582), .b(GPR_11__6_), .o(n_871) );
INV_X1 g35458 ( .a(pZ_6_), .o(n_3266) );
INV_X1 drc_bufs35520 ( .a(n_4089), .o(n_3208) );
NAND2_Z01 g60555 ( .a(n_402), .b(n_391), .o(n_551) );
XOR2_X1 g60384 ( .a(n_282), .b(n_140), .o(n_762) );
BUF_X2 newInst_1002 ( .a(newNet_1001), .o(newNet_1002) );
XNOR2_X1 g60859 ( .a(SP_0_), .b(SP_1_), .o(n_331) );
NAND2_Z01 g58947 ( .a(n_2108), .b(n_1553), .o(n_2150) );
BUF_X2 newInst_1280 ( .a(newNet_642), .o(newNet_1280) );
NOR2_X2 g34968 ( .a(n_3548), .b(n_3492), .o(n_3630) );
BUF_X2 newInst_663 ( .a(newNet_662), .o(newNet_663) );
BUF_X2 newInst_1591 ( .a(newNet_1590), .o(newNet_1591) );
NAND2_Z01 g59565 ( .a(n_1526), .b(n_213), .o(n_1562) );
NAND2_Z01 g34257 ( .a(n_4176), .b(pX_6_), .o(n_4276) );
NAND2_Z01 g58787 ( .a(n_2200), .b(GPR_7__6_), .o(n_2313) );
NOR3_Z1 g59796 ( .a(n_85), .b(n_1200), .c(n_93), .o(n_1328) );
INV_X2 newInst_1691 ( .a(newNet_1690), .o(newNet_1691) );
BUF_X2 newInst_526 ( .a(newNet_525), .o(newNet_526) );
AND2_X1 g58969 ( .a(n_2086), .b(n_1214), .o(n_2137) );
AND2_X1 g59928 ( .a(n_1107), .b(n_235), .o(n_1189) );
XOR2_X1 g60676 ( .a(io_do_0), .b(n_271), .o(n_473) );
BUF_X2 newInst_1128 ( .a(newNet_1127), .o(newNet_1128) );
fflopd GPR_reg_20__3_ ( .CK(newNet_1198), .D(n_2854), .Q(GPR_20__3_) );
INV_X1 g35511 ( .a(pmem_d_3), .o(n_3217) );
BUF_X2 newInst_1525 ( .a(newNet_299), .o(newNet_1525) );
BUF_X2 newInst_1399 ( .a(newNet_332), .o(newNet_1399) );
INV_X1 g35064 ( .a(n_3522), .o(n_4663) );
NAND2_Z01 g34940 ( .a(n_3551), .b(GPR_13__7_), .o(n_3622) );
BUF_X2 newInst_1021 ( .a(newNet_1020), .o(newNet_1021) );
AND2_X1 g35304 ( .a(n_4574), .b(n_3298), .o(n_3372) );
NAND2_Z01 g35451 ( .a(n_3252), .b(n_3227), .o(n_3280) );
NAND2_Z01 g35414 ( .a(pZ_1_), .b(pmem_d_1), .o(n_3291) );
NAND2_Z01 g60468 ( .a(n_380), .b(GPR_4__0_), .o(n_678) );
BUF_X2 newInst_1392 ( .a(newNet_1391), .o(newNet_1392) );
NOR2_Z1 g34416 ( .a(n_4610), .b(n_3533), .o(n_4121) );
NAND2_Z01 g60299 ( .a(n_585), .b(GPR_23__5_), .o(n_825) );
NAND2_Z01 g57930 ( .a(n_2977), .b(n_2436), .o(n_3015) );
NAND2_Z01 g59513 ( .a(n_1570), .b(pX_12_), .o(n_1626) );
INV_X1 g35510 ( .a(pZ_11_), .o(n_3218) );
NAND2_Z01 g58759 ( .a(n_2203), .b(GPR_4__3_), .o(n_2341) );
INV_X1 g34973 ( .a(n_3598), .o(n_3599) );
BUF_X2 newInst_1804 ( .a(newNet_1803), .o(newNet_1804) );
BUF_X2 newInst_1560 ( .a(newNet_567), .o(newNet_1560) );
fflopd GPR_reg_14__3_ ( .CK(newNet_1559), .D(n_2861), .Q(GPR_14__3_) );
NAND4_Z1 g59548 ( .a(n_1304), .b(n_1520), .c(n_1512), .d(n_1066), .o(n_1580) );
BUF_X2 newInst_553 ( .a(newNet_552), .o(newNet_553) );
AND2_X1 g60634 ( .a(n_337), .b(n_4488), .o(n_500) );
BUF_X2 newInst_1769 ( .a(newNet_1768), .o(newNet_1769) );
NOR2_Z2 g34921 ( .a(n_3589), .b(rst), .o(n_3768) );
BUF_X2 newInst_220 ( .a(newNet_219), .o(newNet_220) );
XOR2_X1 g35099 ( .a(n_3462), .b(pY_5_), .o(n_4592) );
AND2_X1 g59517 ( .a(n_1569), .b(SP_12_), .o(n_1622) );
BUF_X2 newInst_433 ( .a(newNet_432), .o(newNet_433) );
NAND2_Z01 g59146 ( .a(n_1896), .b(n_49), .o(n_1953) );
AND2_X1 g58010 ( .a(n_2940), .b(n_2140), .o(n_2961) );
NAND2_Z01 g58601 ( .a(n_2479), .b(n_1954), .o(n_2494) );
AND3_X1 g59659 ( .a(n_992), .b(n_1320), .c(n_958), .o(n_1467) );
NOR2_Z1 g60118 ( .a(n_848), .b(n_139), .o(n_1009) );
fflopd GPR_reg_8__3_ ( .CK(newNet_713), .D(n_2840), .Q(GPR_8__3_) );
INV_X1 g35461 ( .a(pX_3_), .o(n_3263) );
NAND2_Z01 g59089 ( .a(n_1875), .b(n_4563), .o(n_2018) );
NAND2_Z01 g60188 ( .a(n_647), .b(n_622), .o(n_965) );
BUF_X2 newInst_964 ( .a(newNet_963), .o(newNet_964) );
NAND2_Z01 g57925 ( .a(n_2982), .b(n_2256), .o(n_3020) );
NAND2_Z01 g58866 ( .a(n_2156), .b(GPR_15__6_), .o(n_2241) );
BUF_X2 newInst_1111 ( .a(newNet_1110), .o(newNet_1111) );
fflopd Rd_r_reg_0_ ( .CK(newNet_600), .D(n_953), .Q(Rd_r_0_) );
NAND2_Z01 g58734 ( .a(n_2206), .b(GPR_23__6_), .o(n_2373) );
BUF_X2 newInst_616 ( .a(newNet_615), .o(newNet_616) );
NOR2_Z1 g34408 ( .a(n_4610), .b(n_3928), .o(n_4130) );
NOR2_Z1 g59003 ( .a(n_1970), .b(n_84), .o(n_2104) );
BUF_X2 newInst_945 ( .a(newNet_944), .o(newNet_945) );
AND2_X1 g58399 ( .a(n_2657), .b(n_2200), .o(n_2669) );
NAND2_Z01 g34815 ( .a(n_3635), .b(GPR_14__2_), .o(n_3748) );
NAND2_Z01 g58579 ( .a(n_2463), .b(pZ_7_), .o(n_2519) );
BUF_X2 newInst_924 ( .a(newNet_923), .o(newNet_924) );
BUF_X2 newInst_996 ( .a(newNet_995), .o(newNet_996) );
BUF_X2 newInst_1484 ( .a(newNet_1483), .o(newNet_1484) );
AND2_X1 g59749 ( .a(n_1313), .b(n_102), .o(n_1390) );
NAND2_Z01 g59758 ( .a(n_1312), .b(io_do_7), .o(n_1366) );
BUF_X2 newInst_3 ( .a(newNet_2), .o(newNet_3) );
NOR2_Z1 g59926 ( .a(n_1011), .b(n_376), .o(n_1191) );
NAND2_Z01 g60051 ( .a(n_846), .b(pmem_d_15), .o(n_1081) );
BUF_X2 newInst_1413 ( .a(newNet_1412), .o(newNet_1413) );
NOR2_Z1 g60757 ( .a(n_268), .b(n_104), .o(n_386) );
NAND4_Z1 g34064 ( .a(n_4272), .b(n_4216), .c(n_4394), .d(n_4262), .o(n_4399) );
BUF_X2 newInst_991 ( .a(newNet_990), .o(newNet_991) );
NAND2_Z01 g58860 ( .a(n_2155), .b(GPR_14__6_), .o(n_2247) );
BUF_X2 newInst_691 ( .a(newNet_690), .o(newNet_691) );
BUF_X2 newInst_403 ( .a(newNet_402), .o(newNet_403) );
AND2_X1 g58392 ( .a(n_2657), .b(n_2203), .o(n_2676) );
NOR2_X2 g34970 ( .a(n_3548), .b(n_3482), .o(n_3628) );
NOR2_Z1 g60796 ( .a(n_197), .b(n_202), .o(n_370) );
BUF_X2 newInst_1119 ( .a(newNet_152), .o(newNet_1119) );
BUF_X2 newInst_204 ( .a(newNet_203), .o(newNet_204) );
NAND2_Z01 g58572 ( .a(n_2483), .b(pX_12_), .o(n_2524) );
NAND4_Z1 g60144 ( .a(n_689), .b(n_690), .c(n_630), .d(n_688), .o(n_988) );
BUF_X2 newInst_1018 ( .a(newNet_1017), .o(newNet_1018) );
BUF_X2 newInst_585 ( .a(newNet_122), .o(newNet_585) );
NAND2_Z01 g60687 ( .a(GPR_1__5_), .b(n_183), .o(n_451) );
NOR2_Z1 g34207 ( .a(n_4295), .b(n_4178), .o(n_4319) );
INV_X1 g61118 ( .a(n_4435), .o(n_34) );
NAND2_Z01 g57821 ( .a(n_3057), .b(n_2300), .o(n_3092) );
AND2_X1 g35279 ( .a(n_3234), .b(n_4640), .o(n_3396) );
NAND2_Z01 g59511 ( .a(n_1536), .b(SP_3_), .o(n_1611) );
NAND2_Z01 g58327 ( .a(n_2667), .b(n_2232), .o(n_2738) );
NOR2_Z1 g60620 ( .a(n_462), .b(n_182), .o(n_588) );
XOR2_X1 final_adder_mux_R16_278_6_g362 ( .a(final_adder_mux_R16_278_6_n_86), .b(final_adder_mux_R16_278_6_n_34), .o(R16_15_) );
NOR2_Z1 g60610 ( .a(n_431), .b(n_132), .o(n_513) );
NAND2_Z01 g58708 ( .a(n_2209), .b(GPR_20__5_), .o(n_2399) );
BUF_X2 newInst_788 ( .a(newNet_787), .o(newNet_788) );
BUF_X2 newInst_36 ( .a(newNet_35), .o(newNet_36) );
BUF_X2 newInst_1335 ( .a(newNet_1334), .o(newNet_1335) );
NAND2_Z01 g57694 ( .a(n_3158), .b(n_2196), .o(n_3172) );
NOR2_Z1 g59683 ( .a(n_1381), .b(n_4471), .o(n_1442) );
NAND2_Z01 g60024 ( .a(n_828), .b(n_879), .o(n_1104) );
BUF_X2 newInst_1609 ( .a(newNet_1608), .o(newNet_1609) );
AND4_X1 g34078 ( .a(n_4215), .b(n_4248), .c(n_4382), .d(n_4146), .o(dmem_a_5) );
BUF_X2 newInst_508 ( .a(newNet_507), .o(newNet_508) );
NAND4_Z1 g57850 ( .a(n_1254), .b(n_1540), .c(n_2993), .d(n_1253), .o(n_3078) );
NOR2_Z1 g34120 ( .a(n_4326), .b(n_4178), .o(n_4383) );
BUF_X2 newInst_844 ( .a(newNet_843), .o(newNet_844) );
BUF_X2 newInst_709 ( .a(newNet_708), .o(newNet_709) );
fflopd GPR_reg_18__4_ ( .CK(newNet_1345), .D(n_2937), .Q(GPR_18__4_) );
BUF_X2 newInst_1355 ( .a(newNet_1354), .o(newNet_1355) );
XOR2_X1 g60383 ( .a(n_348), .b(io_do_3), .o(n_837) );
BUF_X2 newInst_1664 ( .a(newNet_1663), .o(newNet_1664) );
NOR2_Z1 g35336 ( .a(n_3255), .b(n_3288), .o(n_3334) );
INV_X1 g34386 ( .a(n_4151), .o(n_4152) );
NOR2_Z1 g34623 ( .a(n_3639), .b(n_3640), .o(n_3937) );
INV_X1 g60170 ( .a(n_965), .o(n_964) );
BUF_X2 newInst_959 ( .a(newNet_958), .o(newNet_959) );
NAND2_Z01 g34886 ( .a(n_3564), .b(pX_2_), .o(n_3677) );
INV_X1 g59455 ( .a(n_1663), .o(n_1664) );
BUF_X2 newInst_1086 ( .a(newNet_161), .o(newNet_1086) );
NAND2_Z01 g59173 ( .a(n_55), .b(n_1878), .o(n_1933) );
NAND2_Z01 g58276 ( .a(n_2751), .b(n_24), .o(n_2834) );
AND3_X1 g59891 ( .a(n_4584), .b(n_1043), .c(n_47), .o(n_1267) );
AND4_X1 g60000 ( .a(n_170), .b(n_276), .c(n_482), .d(pmem_d_12), .o(n_1129) );
BUF_X2 newInst_345 ( .a(newNet_344), .o(newNet_345) );
AND2_X1 g58127 ( .a(n_2850), .b(n_2140), .o(n_2885) );
BUF_X2 newInst_1776 ( .a(newNet_1775), .o(newNet_1776) );
fflopd GPR_reg_13__1_ ( .CK(newNet_1609), .D(n_2781), .Q(GPR_13__1_) );
NAND4_Z1 g59808 ( .a(n_701), .b(n_702), .c(n_1177), .d(n_700), .o(n_1320) );
fflopd pY_reg_13_ ( .CK(newNet_174), .D(n_3097), .Q(pY_13_) );
INV_X1 g61082 ( .a(n_4617), .o(n_70) );
NOR2_Z1 g60997 ( .a(n_4628), .b(n_4632), .o(n_176) );
NAND4_Z1 g59474 ( .a(n_1195), .b(n_1198), .c(n_1559), .d(n_1097), .o(n_1663) );
AND2_X1 g35157 ( .a(n_3445), .b(n_3238), .o(n_3468) );
INV_X1 g58593 ( .a(n_2502), .o(n_2503) );
BUF_X2 newInst_504 ( .a(newNet_401), .o(newNet_504) );
BUF_X2 newInst_698 ( .a(newNet_697), .o(newNet_698) );
BUF_X2 newInst_558 ( .a(newNet_557), .o(newNet_558) );
XOR2_X1 g35142 ( .a(n_3428), .b(pX_4_), .o(n_3477) );
NAND4_Z1 g59549 ( .a(n_799), .b(n_1296), .c(n_1498), .d(n_1073), .o(n_1579) );
BUF_X2 newInst_1196 ( .a(newNet_1195), .o(newNet_1196) );
NAND2_Z01 g34188 ( .a(n_4325), .b(n_4464), .o(n_4335) );
NAND2_Z01 g34700 ( .a(n_3568), .b(GPR_22__6_), .o(n_3865) );
NAND2_Z01 g58169 ( .a(n_2797), .b(n_2317), .o(n_2841) );
NAND2_Z01 g60945 ( .a(io_do_6), .b(n_36), .o(n_206) );
NAND2_Z01 g34394 ( .a(n_3208), .b(pZ_11_), .o(n_4144) );
AND2_X1 g59487 ( .a(n_1622), .b(n_1269), .o(n_1638) );
AND2_X1 final_adder_mux_R16_278_6_g404 ( .a(final_adder_mux_R16_278_6_n_28), .b(final_adder_mux_R16_278_6_n_5), .o(final_adder_mux_R16_278_6_n_45) );
NOR2_Z1 g58820 ( .a(n_2217), .b(n_1978), .o(n_2355) );
NOR2_Z1 g59866 ( .a(n_1165), .b(io_do_1), .o(n_1260) );
AND3_X1 g59590 ( .a(n_108), .b(n_1420), .c(rst), .o(n_1538) );
XOR2_X1 g59739 ( .a(n_1315), .b(PC_4_), .o(n_1391) );
AND2_X1 g58267 ( .a(n_2752), .b(n_2203), .o(n_2800) );
NAND2_Z01 g60895 ( .a(PC_1_), .b(pmem_d_4), .o(n_273) );
AND2_X1 g60362 ( .a(n_587), .b(n_274), .o(n_778) );
AND2_X1 g58382 ( .a(n_2657), .b(n_2208), .o(n_2686) );
BUF_X2 newInst_1575 ( .a(newNet_1574), .o(newNet_1575) );
BUF_X2 newInst_913 ( .a(newNet_912), .o(newNet_913) );
NAND2_Z01 g59436 ( .a(n_1647), .b(n_851), .o(n_1683) );
BUF_X2 newInst_411 ( .a(newNet_410), .o(newNet_411) );
NAND2_Z01 g60254 ( .a(n_575), .b(GPR_2__7_), .o(n_892) );
XNOR2_X1 g35259 ( .a(n_3312), .b(PC_2_), .o(n_4551) );
NAND3_Z1 g58354 ( .a(n_1509), .b(n_2607), .c(n_1185), .o(n_2717) );
NAND4_Z1 g60006 ( .a(n_903), .b(n_944), .c(n_931), .d(n_907), .o(n_1123) );
NAND2_Z01 g59580 ( .a(n_1490), .b(n_1275), .o(n_1545) );
INV_X1 g59599 ( .a(n_1529), .o(n_1530) );
NOR2_Z1 g59780 ( .a(n_1308), .b(n_1271), .o(n_1353) );
NAND2_Z01 g34142 ( .a(n_4317), .b(n_4621), .o(n_4366) );
NOR2_Z1 g59881 ( .a(n_981), .b(n_1124), .o(n_1246) );
AND2_X1 g57888 ( .a(n_3009), .b(n_2157), .o(n_3050) );
NAND2_Z01 g58692 ( .a(n_2211), .b(GPR_19__7_), .o(n_2414) );
NAND4_Z1 g60131 ( .a(n_724), .b(n_739), .c(n_706), .d(n_543), .o(n_1001) );
NOR2_Z1 g35031 ( .a(n_3526), .b(Rd_2_), .o(n_3549) );
NAND4_Z1 g34088 ( .a(n_4211), .b(n_4376), .c(n_4321), .d(n_4213), .o(dmem_do_2) );
BUF_X2 newInst_1324 ( .a(newNet_1323), .o(newNet_1324) );
NAND2_Z01 g60457 ( .a(n_372), .b(U_8_), .o(n_689) );
BUF_X2 newInst_1069 ( .a(newNet_1068), .o(newNet_1069) );
BUF_X2 newInst_387 ( .a(newNet_386), .o(newNet_387) );
XNOR2_X1 g60860 ( .a(n_4442), .b(n_4426), .o(n_330) );
NAND2_Z01 g60920 ( .a(n_80), .b(pX_10_), .o(n_222) );
AND3_X1 g59443 ( .a(n_1398), .b(n_1616), .c(n_1137), .o(n_1696) );
NAND2_Z01 g34664 ( .a(n_3622), .b(n_3623), .o(n_3901) );
BUF_X2 newInst_263 ( .a(newNet_262), .o(newNet_263) );
fflopd GPR_reg_18__0_ ( .CK(newNet_1370), .D(n_2632), .Q(GPR_18__0_) );
BUF_X2 newInst_1260 ( .a(newNet_1259), .o(newNet_1260) );
NAND2_Z01 g59273 ( .a(io_do_6), .b(n_1764), .o(n_1840) );
BUF_X2 newInst_482 ( .a(newNet_481), .o(newNet_482) );
AND2_X1 final_adder_mux_R16_278_6_g438 ( .a(n_4444), .b(n_4428), .o(final_adder_mux_R16_278_6_n_11) );
NAND2_Z01 g60957 ( .a(n_41), .b(pmem_d_0), .o(n_204) );
NOR2_Z1 g59291 ( .a(n_19), .b(n_1737), .o(n_1819) );
INV_X1 g35425 ( .a(n_3277), .o(n_3278) );
BUF_X2 newInst_1855 ( .a(newNet_1854), .o(newNet_1855) );
BUF_X2 newInst_1118 ( .a(newNet_1117), .o(newNet_1118) );
INV_X1 g59911 ( .a(n_1210), .o(n_1211) );
AND2_X1 g58122 ( .a(n_2850), .b(n_2203), .o(n_2890) );
NAND2_Z01 g58238 ( .a(n_2755), .b(n_2194), .o(n_2829) );
NAND3_Z1 g59798 ( .a(n_72), .b(n_1205), .c(pZ_12_), .o(n_1348) );
NAND2_Z01 g60273 ( .a(R16_11_), .b(n_571), .o(n_873) );
NOR2_Z1 g60740 ( .a(n_280), .b(n_96), .o(n_468) );
NAND2_Z01 g60404 ( .a(n_372), .b(U_15_), .o(n_742) );
INV_X1 g60282 ( .a(n_852), .o(n_853) );
NAND2_Z01 g58245 ( .a(n_2756), .b(n_2196), .o(n_2822) );
NAND2_Z01 g34656 ( .a(n_3643), .b(n_4561), .o(n_4645) );
NAND4_Z2 g35193 ( .a(n_3337), .b(n_3385), .c(n_3362), .d(n_3397), .o(n_4614) );
BUF_X2 newInst_122 ( .a(newNet_8), .o(newNet_122) );
NAND4_Z1 g34598 ( .a(n_3694), .b(n_3689), .c(n_3687), .d(n_3688), .o(n_3962) );
NAND2_Z01 g34271 ( .a(n_4162), .b(pY_12_), .o(n_4262) );
INV_X1 g60093 ( .a(n_1031), .o(n_1032) );
BUF_X2 newInst_753 ( .a(newNet_752), .o(newNet_753) );
INV_X1 g35150 ( .a(n_3464), .o(n_4630) );
XNOR2_X1 g2 ( .a(n_4294), .b(SP_11_), .o(n_3195) );
AND2_X1 g57991 ( .a(n_2940), .b(n_2157), .o(n_2980) );
BUF_X2 newInst_761 ( .a(newNet_760), .o(newNet_761) );
NAND2_Z01 g58052 ( .a(n_2892), .b(n_2368), .o(n_2930) );
BUF_X2 newInst_518 ( .a(newNet_517), .o(newNet_518) );
NAND2_Z01 final_adder_mux_R16_278_6_g387 ( .a(final_adder_mux_R16_278_6_n_60), .b(final_adder_mux_R16_278_6_n_17), .o(final_adder_mux_R16_278_6_n_62) );
BUF_X2 newInst_1097 ( .a(newNet_526), .o(newNet_1097) );
AND2_X1 g58410 ( .a(n_2657), .b(n_571), .o(n_2689) );
NAND2_Z01 g34652 ( .a(n_3768), .b(n_4553), .o(n_3908) );
NAND2_Z01 g34634 ( .a(n_3769), .b(pZ_9_), .o(n_3926) );
NAND2_Z01 g60235 ( .a(n_582), .b(GPR_11__0_), .o(n_910) );
NAND3_Z1 g57652 ( .a(n_2560), .b(n_3176), .c(n_2145), .o(n_3190) );
NAND2_Z01 g58677 ( .a(n_2212), .b(GPR_18__1_), .o(n_2429) );
NAND2_Z01 g59401 ( .a(n_1633), .b(SP_11_), .o(n_1715) );
NOR2_Z1 g59118 ( .a(n_1891), .b(n_86), .o(n_1991) );
NAND2_Z01 g34843 ( .a(n_3591), .b(U_9_), .o(n_3720) );
NAND2_Z01 g60447 ( .a(n_361), .b(GPR_7__4_), .o(n_699) );
NAND4_Z1 g57951 ( .a(n_1004), .b(n_1406), .c(n_2921), .d(n_1064), .o(n_2994) );
BUF_X2 newInst_1351 ( .a(newNet_1102), .o(newNet_1351) );
BUF_X2 newInst_701 ( .a(newNet_700), .o(newNet_701) );
BUF_X2 newInst_1412 ( .a(newNet_1411), .o(newNet_1412) );
NAND3_Z1 g35189 ( .a(n_3382), .b(n_3438), .c(n_3408), .o(n_4621) );
NOR2_Z1 g35215 ( .a(n_4660), .b(n_3238), .o(n_3449) );
NAND2_Z01 g58791 ( .a(n_2199), .b(GPR_0__1_), .o(n_2309) );
BUF_X2 newInst_1542 ( .a(newNet_1541), .o(newNet_1542) );
NAND2_Z01 g34350 ( .a(n_4158), .b(n_3313), .o(n_4184) );
NAND2_Z01 g59847 ( .a(n_1164), .b(n_54), .o(n_1279) );
NAND4_Z1 g60145 ( .a(n_678), .b(n_679), .c(n_680), .d(n_541), .o(n_987) );
NAND4_Z1 g34580 ( .a(n_3785), .b(n_3787), .c(n_3784), .d(n_3786), .o(n_3980) );
NAND2_Z01 g57982 ( .a(n_2941), .b(n_2194), .o(n_2990) );
INV_X1 drc_bufs61142 ( .a(n_1648), .o(n_28) );
NAND2_Z01 g34156 ( .a(n_4317), .b(n_4618), .o(n_4352) );
NOR4_Z1 g35179 ( .a(n_3233), .b(n_3231), .c(n_3297), .d(pmem_d_0), .o(n_3455) );
NAND2_Z01 g59080 ( .a(n_1875), .b(n_4570), .o(n_2027) );
BUF_X2 newInst_1450 ( .a(newNet_1449), .o(newNet_1450) );
BUF_X2 newInst_485 ( .a(newNet_484), .o(newNet_485) );
NAND2_Z01 g59467 ( .a(n_1586), .b(SP_5_), .o(n_1656) );
AND2_X1 g59707 ( .a(n_1364), .b(SP_0_), .o(n_1423) );
NOR2_Z1 g59223 ( .a(n_1841), .b(PC_0_), .o(n_1883) );
AND2_X1 g59568 ( .a(n_1494), .b(SP_9_), .o(n_1560) );
INV_X1 g34465 ( .a(n_4076), .o(n_4077) );
NOR2_Z1 g60355 ( .a(n_601), .b(n_8), .o(n_780) );
NAND2_Z01 g34162 ( .a(n_4317), .b(pmem_d_2), .o(n_4346) );
BUF_X2 newInst_668 ( .a(newNet_667), .o(newNet_668) );
BUF_X2 newInst_1203 ( .a(newNet_1070), .o(newNet_1203) );
NAND2_Z01 g59642 ( .a(io_do_3), .b(n_1418), .o(n_1479) );
NAND2_Z01 g58315 ( .a(n_2680), .b(n_2371), .o(n_2750) );
AND2_X1 g58373 ( .a(n_2657), .b(n_2212), .o(n_2698) );
NAND2_Z01 g34254 ( .a(n_4161), .b(n_4563), .o(n_4279) );
NOR2_Z1 g34287 ( .a(n_4163), .b(n_3232), .o(n_4246) );
NAND2_Z01 g58283 ( .a(n_2715), .b(n_2272), .o(n_2787) );
NOR4_Z1 g34231 ( .a(n_4218), .b(n_4220), .c(n_4253), .d(n_4118), .o(n_4300) );
AND2_X1 g60766 ( .a(n_4651), .b(n_158), .o(n_383) );
NAND2_Z01 g60200 ( .a(n_584), .b(GPR_18__3_), .o(n_945) );
NOR2_Z1 g60632 ( .a(n_376), .b(C), .o(n_502) );
AND2_X1 g58005 ( .a(n_2940), .b(n_2203), .o(n_2966) );
BUF_X2 newInst_1600 ( .a(newNet_1599), .o(newNet_1600) );
BUF_X2 newInst_303 ( .a(newNet_302), .o(newNet_303) );
NOR4_Z1 g58608 ( .a(n_1684), .b(n_2188), .c(n_2104), .d(n_2177), .o(n_2489) );
NAND2_Z01 g58688 ( .a(n_2211), .b(GPR_19__4_), .o(n_2418) );
BUF_X2 newInst_1296 ( .a(newNet_1232), .o(newNet_1296) );
fflopd GPR_reg_10__0_ ( .CK(newNet_1763), .D(n_2640), .Q(GPR_10__0_) );
NOR2_Z1 g60629 ( .a(n_326), .b(n_179), .o(n_503) );
BUF_X2 newInst_891 ( .a(newNet_890), .o(newNet_891) );
BUF_X2 newInst_339 ( .a(newNet_218), .o(newNet_339) );
BUF_X2 newInst_307 ( .a(newNet_306), .o(newNet_307) );
INV_X1 g35039 ( .a(n_3533), .o(n_4603) );
BUF_X2 newInst_1682 ( .a(newNet_1681), .o(newNet_1682) );
INV_X1 g59477 ( .a(n_1650), .o(n_1649) );
NOR2_Z1 g60586 ( .a(n_8), .b(N), .o(n_526) );
BUF_X2 newInst_1618 ( .a(newNet_1617), .o(newNet_1618) );
XOR2_X1 g34235 ( .a(n_4230), .b(SP_10_), .o(n_4296) );
NAND2_Z01 g58156 ( .a(n_2809), .b(n_2427), .o(n_2857) );
BUF_X2 newInst_363 ( .a(newNet_362), .o(newNet_363) );
NAND3_Z1 g59202 ( .a(n_849), .b(n_1825), .c(n_61), .o(n_1908) );
NAND2_Z01 g58682 ( .a(n_2212), .b(GPR_18__6_), .o(n_2424) );
NOR3_Z1 g34492 ( .a(n_4009), .b(n_3992), .c(n_4022), .o(n_4052) );
NAND2_Z01 g58293 ( .a(n_2700), .b(n_2311), .o(n_2777) );
NAND3_Z1 g60123 ( .a(n_566), .b(io_do_7), .c(pmem_d_11), .o(n_1004) );
NOR2_Z1 g34915 ( .a(n_3562), .b(n_4635), .o(n_3648) );
NAND2_Z01 g59944 ( .a(n_1026), .b(n_462), .o(n_1182) );
BUF_X2 newInst_1445 ( .a(newNet_1444), .o(newNet_1445) );
NAND2_Z01 g34713 ( .a(n_3597), .b(GPR_17__6_), .o(n_3852) );
AND2_X1 g60363 ( .a(n_609), .b(SP_4_), .o(n_777) );
NOR2_Z1 g60607 ( .a(n_352), .b(rst), .o(n_594) );
NOR2_Z1 g59364 ( .a(n_1697), .b(n_1269), .o(n_1749) );
BUF_X2 newInst_1734 ( .a(newNet_1733), .o(newNet_1734) );
NAND4_Z1 g58139 ( .a(n_2039), .b(n_2475), .c(n_2832), .d(n_1946), .o(n_2874) );
NAND2_Z01 g58289 ( .a(n_2708), .b(n_2253), .o(n_2781) );
BUF_X2 newInst_861 ( .a(newNet_860), .o(newNet_861) );
NAND3_Z1 g58567 ( .a(n_1985), .b(n_2503), .c(n_2002), .o(n_2531) );
NAND2_Z01 g58948 ( .a(n_2107), .b(n_1852), .o(n_2162) );
NOR2_Z1 g59787 ( .a(n_1269), .b(n_847), .o(n_1337) );
NAND2_Z01 g34825 ( .a(n_3594), .b(GPR_7__2_), .o(n_3738) );
NAND2_Z01 g34486 ( .a(n_4037), .b(pZ_8_), .o(n_4055) );
BUF_X2 newInst_803 ( .a(newNet_802), .o(newNet_803) );
NAND2_Z01 g58932 ( .a(n_2142), .b(n_2083), .o(n_2193) );
BUF_X2 newInst_1799 ( .a(newNet_1798), .o(newNet_1799) );
NAND2_Z01 g59759 ( .a(n_1284), .b(io_do_7), .o(n_1365) );
fflopd GPR_reg_2__5_ ( .CK(newNet_991), .D(n_3003), .Q(GPR_2__5_) );
fflopd GPR_reg_5__0_ ( .CK(newNet_877), .D(n_2620), .Q(GPR_5__0_) );
NAND4_Z1 g59956 ( .a(n_384), .b(n_186), .c(n_513), .d(n_172), .o(n_1175) );
AND2_X1 g59408 ( .a(n_54), .b(n_1661), .o(n_1733) );
BUF_X2 newInst_620 ( .a(newNet_619), .o(newNet_620) );
BUF_X2 newInst_946 ( .a(newNet_945), .o(newNet_946) );
BUF_X2 newInst_1810 ( .a(newNet_1809), .o(newNet_1810) );
INV_X2 newInst_1644 ( .a(newNet_1643), .o(newNet_1644) );
INV_X1 g61033 ( .a(state_1_), .o(n_119) );
NAND2_Z01 g35137 ( .a(n_3462), .b(n_3247), .o(n_3480) );
NAND2_Z01 g34159 ( .a(n_4317), .b(pmem_d_6), .o(n_4349) );
AND2_X1 g57902 ( .a(n_3009), .b(n_2203), .o(n_3036) );
NAND2_Z01 g58525 ( .a(n_2559), .b(n_1989), .o(n_2572) );
BUF_X2 newInst_1175 ( .a(newNet_1174), .o(newNet_1175) );
INV_X1 drc_bufs61201 ( .a(n_12), .o(n_13) );
BUF_X2 newInst_1430 ( .a(newNet_1429), .o(newNet_1430) );
XOR2_X1 g58492 ( .a(n_2572), .b(n_1876), .o(n_2604) );
BUF_X2 newInst_1745 ( .a(newNet_1744), .o(newNet_1745) );
NAND2_Z01 g34135 ( .a(n_4325), .b(n_4617), .o(n_4373) );
NAND2_Z01 g58870 ( .a(n_2156), .b(GPR_15__5_), .o(n_2237) );
NAND2_Z01 g59052 ( .a(n_18), .b(n_4571), .o(n_2055) );
INV_X2 newInst_140 ( .a(newNet_139), .o(newNet_140) );
BUF_X2 newInst_1559 ( .a(newNet_1558), .o(newNet_1559) );
BUF_X2 newInst_89 ( .a(newNet_0), .o(newNet_89) );
XNOR2_X1 g35016 ( .a(n_4520), .b(pZ_8_), .o(n_3561) );
NAND2_Z01 g60507 ( .a(n_21), .b(Rd_r_3_), .o(n_639) );
AND2_X1 g58504 ( .a(n_2567), .b(n_2212), .o(n_2593) );
BUF_X2 newInst_840 ( .a(newNet_428), .o(newNet_840) );
NAND2_Z01 g34529 ( .a(n_3655), .b(n_3941), .o(n_4016) );
INV_X1 g60538 ( .a(n_583), .o(n_584) );
NAND2_Z01 g58638 ( .a(n_2361), .b(n_2005), .o(n_2464) );
NAND2_Z01 g57770 ( .a(n_3101), .b(n_2299), .o(n_3111) );
NAND2_Z01 g35119 ( .a(Rd_3_), .b(pmem_d_5), .o(n_3492) );
NAND2_Z01 g34862 ( .a(n_3591), .b(U_8_), .o(n_3701) );
NAND2_Z01 g59388 ( .a(n_1648), .b(dmem_di_0), .o(n_1727) );
BUF_X2 newInst_1304 ( .a(newNet_1303), .o(newNet_1304) );
BUF_X2 newInst_561 ( .a(newNet_560), .o(newNet_561) );
NOR2_Z1 g34895 ( .a(n_3578), .b(n_3261), .o(n_3668) );
BUF_X2 newInst_236 ( .a(newNet_235), .o(newNet_236) );
NOR2_Z1 g34776 ( .a(n_3574), .b(n_3234), .o(n_3789) );
AND2_X1 g60788 ( .a(n_160), .b(pmem_d_1), .o(n_376) );
NAND2_Z01 g34722 ( .a(n_3197), .b(GPR_23__2_), .o(n_3843) );
BUF_X2 newInst_1862 ( .a(newNet_1537), .o(newNet_1862) );
XOR2_X1 final_adder_mux_R16_278_6_g417 ( .a(n_4438), .b(n_4422), .o(final_adder_mux_R16_278_6_n_32) );
NAND2_Z01 final_adder_mux_R16_278_6_g424 ( .a(n_4440), .b(n_4424), .o(final_adder_mux_R16_278_6_n_24) );
BUF_X2 newInst_1462 ( .a(newNet_1297), .o(newNet_1462) );
NAND2_Z01 g58670 ( .a(n_2214), .b(GPR_16__5_), .o(n_2436) );
BUF_X2 newInst_897 ( .a(newNet_896), .o(newNet_897) );
BUF_X2 newInst_1537 ( .a(newNet_1536), .o(newNet_1537) );
INV_X1 g61061 ( .a(PC_4_), .o(n_91) );
BUF_X2 newInst_1259 ( .a(newNet_1258), .o(newNet_1259) );
AND2_X1 g61013 ( .a(n_4443), .b(n_4427), .o(n_168) );
NAND2_Z01 g35271 ( .a(n_3299), .b(pX_13_), .o(n_3403) );
BUF_X2 newInst_1151 ( .a(newNet_730), .o(newNet_1151) );
NAND2_Z01 g59074 ( .a(n_1871), .b(n_4601), .o(n_2033) );
NAND2_Z01 g58045 ( .a(n_2900), .b(n_2426), .o(n_2937) );
NAND2_Z01 g60195 ( .a(n_620), .b(n_666), .o(n_950) );
BUF_X2 newInst_495 ( .a(newNet_494), .o(newNet_495) );
NAND2_Z01 g34731 ( .a(n_3629), .b(GPR_2__5_), .o(n_3834) );
BUF_X2 newInst_689 ( .a(newNet_304), .o(newNet_689) );
fflopd GPR_reg_1__1_ ( .CK(newNet_1260), .D(n_2767), .Q(GPR_1__1_) );
NAND2_Z01 g59631 ( .a(n_1440), .b(n_210), .o(n_1526) );
BUF_X2 newInst_542 ( .a(newNet_541), .o(newNet_542) );
NAND2_Z01 g34707 ( .a(n_3630), .b(pX_14_), .o(n_3858) );
NOR2_Z1 g34338 ( .a(n_4612), .b(n_3763), .o(n_4196) );
NAND2_Z01 g57711 ( .a(n_3129), .b(n_2397), .o(n_3156) );
NAND2_Z01 g60941 ( .a(io_do_3), .b(n_71), .o(n_210) );
AND2_X1 g35315 ( .a(n_4640), .b(n_3251), .o(n_4638) );
XOR2_X1 g58991 ( .a(n_2012), .b(n_379), .o(n_2117) );
BUF_X2 newInst_1209 ( .a(newNet_1208), .o(newNet_1209) );
INV_X1 g60773 ( .a(n_356), .o(n_355) );
NAND2_Z01 g59218 ( .a(n_1854), .b(io_do_7), .o(n_1900) );
BUF_X2 newInst_793 ( .a(newNet_792), .o(newNet_793) );
BUF_X2 newInst_1421 ( .a(newNet_1420), .o(newNet_1421) );
INV_X1 g60015 ( .a(n_1106), .o(n_1107) );
NAND2_Z01 g60325 ( .a(n_597), .b(pX_13_), .o(n_802) );
BUF_X2 newInst_1289 ( .a(newNet_1288), .o(newNet_1289) );
NAND2_Z01 g60581 ( .a(io_do_4), .b(n_364), .o(n_531) );
BUF_X2 newInst_1718 ( .a(newNet_1717), .o(newNet_1718) );
NAND2_Z01 g60454 ( .a(n_368), .b(GPR_13__6_), .o(n_692) );
NAND3_Z1 g34068 ( .a(n_4392), .b(n_4387), .c(n_4214), .o(dmem_do_3) );
NAND4_Z1 g60157 ( .a(n_246), .b(n_385), .c(n_528), .d(n_529), .o(n_978) );
INV_X1 g61088 ( .a(io_do_4), .o(n_64) );
BUF_X2 newInst_154 ( .a(newNet_153), .o(newNet_154) );
fflopd GPR_reg_5__6_ ( .CK(newNet_839), .D(n_3069), .Q(GPR_5__6_) );
BUF_X2 newInst_1697 ( .a(newNet_1134), .o(newNet_1697) );
NAND2_Z01 g60680 ( .a(n_4490), .b(n_252), .o(n_471) );
NAND2_Z01 g60407 ( .a(n_370), .b(GPR_22__4_), .o(n_739) );
NAND2_Z01 g58456 ( .a(n_2601), .b(n_2273), .o(n_2640) );
BUF_X2 newInst_292 ( .a(newNet_291), .o(newNet_292) );
BUF_X2 newInst_72 ( .a(newNet_71), .o(newNet_72) );
NAND2_Z01 g60834 ( .a(n_195), .b(n_59), .o(n_346) );
NAND3_Z1 g35376 ( .a(n_3232), .b(n_3275), .c(n_3251), .o(n_4483) );
NAND2_Z01 g60520 ( .a(n_358), .b(GPR_0__3_), .o(n_626) );
fflopd GPR_reg_7__4_ ( .CK(newNet_765), .D(n_2925), .Q(GPR_7__4_) );
INV_X1 g35130 ( .a(n_3476), .o(n_4606) );
NAND2_Z01 g60047 ( .a(n_820), .b(n_225), .o(n_1115) );
NAND2_Z01 g60576 ( .a(n_357), .b(pY_13_), .o(n_535) );
NAND4_Z1 g59671 ( .a(n_1057), .b(n_1293), .c(n_1369), .d(n_1059), .o(n_1457) );
BUF_X2 newInst_315 ( .a(newNet_314), .o(newNet_315) );
BUF_X2 newInst_1251 ( .a(newNet_1250), .o(newNet_1251) );
NAND2_Z01 g35006 ( .a(n_3536), .b(n_3489), .o(n_3570) );
BUF_X2 newInst_1042 ( .a(newNet_842), .o(newNet_1042) );
NAND4_Z1 g59374 ( .a(n_1620), .b(n_1623), .c(n_1625), .d(n_1029), .o(n_1744) );
XNOR2_X1 g60673 ( .a(n_278), .b(pZ_2_), .o(n_476) );
BUF_X2 newInst_1158 ( .a(newNet_880), .o(newNet_1158) );
NAND2_Z01 g59719 ( .a(n_1350), .b(n_782), .o(n_1416) );
BUF_X2 newInst_1228 ( .a(newNet_1227), .o(newNet_1228) );
NOR2_Z1 g34428 ( .a(n_4610), .b(n_3422), .o(n_4109) );
NAND2_Z01 g60480 ( .a(n_371), .b(GPR_21__5_), .o(n_666) );
NOR2_Z1 g59111 ( .a(n_1901), .b(n_112), .o(n_1998) );
INV_X1 g35149 ( .a(n_3467), .o(Rd_2_) );
NAND2_Z01 g34474 ( .a(n_4054), .b(n_3279), .o(n_4067) );
NAND2_Z01 g34519 ( .a(n_3877), .b(n_3949), .o(n_4024) );
NAND4_Z1 g59537 ( .a(n_1303), .b(n_1497), .c(n_1519), .d(n_1071), .o(n_1590) );
BUF_X2 newInst_1453 ( .a(newNet_1452), .o(newNet_1453) );
NOR2_Z1 g60814 ( .a(n_175), .b(state_3_), .o(n_356) );
NOR2_Z1 g59113 ( .a(n_1870), .b(n_76), .o(n_1996) );
NAND4_Z1 g59999 ( .a(n_908), .b(n_884), .c(n_805), .d(n_883), .o(n_1130) );
XOR2_X1 g35049 ( .a(n_3507), .b(n_3260), .o(n_4567) );
fflopd GPR_reg_8__1_ ( .CK(newNet_725), .D(n_2738), .Q(GPR_8__1_) );
AND2_X1 g35349 ( .a(n_4488), .b(n_4490), .o(n_4484) );
NAND2_Z01 g58625 ( .a(n_2360), .b(pY_0_), .o(n_2472) );
BUF_X2 newInst_82 ( .a(newNet_56), .o(newNet_82) );
NAND2_Z01 g58634 ( .a(n_2352), .b(pX_8_), .o(n_2468) );
BUF_X2 newInst_91 ( .a(newNet_90), .o(newNet_91) );
BUF_X2 newInst_15 ( .a(newNet_14), .o(newNet_15) );
fflopd GPR_reg_9__6_ ( .CK(newNet_669), .D(n_3065), .Q(GPR_9__6_) );
NAND2_Z01 g58335 ( .a(n_2690), .b(n_891), .o(n_2754) );
AND2_X1 g58364 ( .a(n_2656), .b(n_2157), .o(n_2707) );
AND2_X1 g58515 ( .a(n_2567), .b(n_2201), .o(n_2581) );
NAND2_Z01 g59825 ( .a(n_1171), .b(dmem_di_5), .o(n_1299) );
BUF_X2 newInst_1840 ( .a(newNet_1839), .o(newNet_1840) );
NAND2_Z01 g58150 ( .a(n_2815), .b(n_2257), .o(n_2863) );
NOR2_Z2 g59243 ( .a(n_1829), .b(n_4612), .o(n_1875) );
NAND3_Z1 g34166 ( .a(n_4293), .b(n_4308), .c(n_4225), .o(dmem_do_5) );
NAND2_Z01 g35225 ( .a(n_3360), .b(n_3220), .o(n_3443) );
NAND2_Z01 g57834 ( .a(n_3042), .b(n_2398), .o(n_3076) );
NAND2_Z01 g58891 ( .a(n_2140), .b(GPR_9__5_), .o(n_2191) );
NOR2_Z1 g59353 ( .a(n_1730), .b(n_351), .o(n_1760) );
NAND2_Z01 g59396 ( .a(n_1648), .b(dmem_di_6), .o(n_1719) );
NAND2_Z01 g58811 ( .a(n_2195), .b(U_9_), .o(n_2289) );
fflopd GPR_reg_5__7_ ( .CK(newNet_837), .D(n_3149), .Q(GPR_5__7_) );
fflopd GPR_reg_10__7_ ( .CK(newNet_1721), .D(n_3168), .Q(GPR_10__7_) );
BUF_X2 newInst_628 ( .a(newNet_627), .o(newNet_628) );
NOR2_Z1 g35437 ( .a(pZ_1_), .b(pZ_0_), .o(n_3285) );
NAND2_Z01 g57800 ( .a(n_3080), .b(n_2217), .o(n_3107) );
NOR2_Z1 g35342 ( .a(n_3311), .b(n_3233), .o(n_3360) );
NAND2_Z01 g58667 ( .a(n_2214), .b(GPR_16__1_), .o(n_2439) );
INV_X1 g60014 ( .a(n_1109), .o(n_1108) );
NAND2_Z01 g59933 ( .a(n_1116), .b(n_969), .o(n_1210) );
NAND2_Z01 g60495 ( .a(n_349), .b(U_0_), .o(n_651) );
NAND2_Z01 g57707 ( .a(n_3134), .b(n_2430), .o(n_3162) );
XOR2_X1 g59596 ( .a(n_1409), .b(PC_10_), .o(n_1533) );
BUF_X2 newInst_1706 ( .a(newNet_1705), .o(newNet_1706) );
BUF_X2 newInst_967 ( .a(newNet_322), .o(newNet_967) );
BUF_X2 newInst_906 ( .a(newNet_549), .o(newNet_906) );
BUF_X2 newInst_1586 ( .a(newNet_1585), .o(newNet_1586) );
NAND2_Z01 g34636 ( .a(n_3769), .b(pZ_6_), .o(n_3924) );
INV_X1 g35479 ( .a(pZ_3_), .o(n_3245) );
INV_X1 g58747 ( .a(n_2355), .o(n_2356) );
INV_X1 g34371 ( .a(n_4612), .o(n_4161) );
INV_X1 g34981 ( .a(n_3570), .o(n_3571) );
AND2_X1 g57897 ( .a(n_3009), .b(n_2208), .o(n_3041) );
AND3_X1 g59665 ( .a(SP_9_), .b(n_1352), .c(SP_10_), .o(n_1484) );
BUF_X2 newInst_1636 ( .a(newNet_1635), .o(newNet_1636) );
NOR2_Z1 g59974 ( .a(n_1106), .b(PC_6_), .o(n_1163) );
BUF_X2 newInst_1038 ( .a(newNet_794), .o(newNet_1038) );
BUF_X2 newInst_1659 ( .a(newNet_1658), .o(newNet_1659) );
NAND2_Z01 g58455 ( .a(n_2602), .b(n_1840), .o(n_2641) );
BUF_X2 newInst_116 ( .a(newNet_115), .o(newNet_116) );
NAND2_Z01 g35162 ( .a(n_3418), .b(n_3446), .o(n_4642) );
AND3_X1 g59201 ( .a(n_1114), .b(n_1893), .c(pY_6_), .o(n_1909) );
NAND2_Z01 g34116 ( .a(n_4331), .b(n_4345), .o(n_4434) );
NAND2_Z01 g58101 ( .a(n_2851), .b(n_2198), .o(n_2912) );
BUF_X2 newInst_1258 ( .a(newNet_1257), .o(newNet_1258) );
NAND2_Z01 g58467 ( .a(n_2404), .b(n_2590), .o(n_2629) );
INV_X1 g34975 ( .a(n_3588), .o(n_3589) );
NAND2_Z01 g34721 ( .a(n_3625), .b(GPR_0__5_), .o(n_3844) );
BUF_X2 newInst_186 ( .a(newNet_185), .o(newNet_186) );
NOR2_Z1 g59714 ( .a(n_1316), .b(n_1166), .o(n_1419) );
NAND4_Z1 g57762 ( .a(n_1909), .b(n_2514), .c(n_3102), .d(n_2038), .o(n_3113) );
NOR2_Z1 g58482 ( .a(n_2603), .b(n_1734), .o(n_2614) );
NOR2_Z1 g58951 ( .a(n_2116), .b(n_964), .o(n_2160) );
XOR2_X1 g34515 ( .a(n_3902), .b(pY_5_), .o(n_4030) );
INV_X1 g59283 ( .a(n_1828), .o(n_1829) );
NOR4_Z1 g59898 ( .a(n_4485), .b(n_355), .c(n_785), .d(state_0_), .o(n_1231) );
NAND2_Z02 g58961 ( .a(n_2115), .b(n_1209), .o(n_2156) );
NAND2_Z01 g35316 ( .a(n_3289), .b(pY_7_), .o(n_3362) );
NAND3_Z1 g58013 ( .a(n_1237), .b(n_2871), .c(n_1098), .o(n_2959) );
NAND2_Z01 g58040 ( .a(n_2904), .b(n_2182), .o(n_2945) );
AND2_X1 g60074 ( .a(n_861), .b(n_55), .o(n_1110) );
BUF_X2 newInst_1748 ( .a(newNet_1747), .o(newNet_1748) );
NAND2_Z02 g34380 ( .a(n_4125), .b(n_4087), .o(n_16064_BAR) );
NAND2_Z01 g35121 ( .a(n_3468), .b(n_4632), .o(n_4478) );
AND3_X1 g58981 ( .a(n_94), .b(n_1982), .c(pZ_9_), .o(n_2126) );
BUF_X2 newInst_1688 ( .a(newNet_1687), .o(newNet_1688) );
NAND2_Z02 g58908 ( .a(n_2161), .b(n_1172), .o(n_2214) );
NAND2_Z01 g35262 ( .a(U_8_), .b(n_3275), .o(n_3410) );
AND2_X1 g34987 ( .a(n_3546), .b(pZ_9_), .o(n_3595) );
NAND2_Z01 g57721 ( .a(n_3119), .b(n_2224), .o(n_3146) );
BUF_X2 newInst_1072 ( .a(newNet_1071), .o(newNet_1072) );
NAND2_Z01 g60201 ( .a(n_598), .b(GPR_15__2_), .o(n_944) );
BUF_X2 newInst_1150 ( .a(newNet_1149), .o(newNet_1150) );
INV_X1 g35387 ( .a(n_3306), .o(n_4521) );
AND2_X1 g60080 ( .a(n_848), .b(n_59), .o(n_1055) );
AND2_X1 g57742 ( .a(n_3115), .b(n_2209), .o(n_3129) );
BUF_X2 newInst_1763 ( .a(newNet_1314), .o(newNet_1763) );
BUF_X2 newInst_1122 ( .a(newNet_1121), .o(newNet_1122) );
NAND2_Z01 g34290 ( .a(n_4164), .b(pmem_d_11), .o(n_4243) );
AND2_X1 g58496 ( .a(n_2567), .b(n_2159), .o(n_2601) );
NOR4_Z1 g59730 ( .a(n_492), .b(n_1145), .c(n_1230), .d(n_516), .o(n_1400) );
BUF_X2 newInst_1283 ( .a(newNet_1282), .o(newNet_1283) );
BUF_X2 newInst_682 ( .a(newNet_644), .o(newNet_682) );
BUF_X2 newInst_1420 ( .a(newNet_1419), .o(newNet_1420) );
fflopd GPR_reg_21__1_ ( .CK(newNet_1157), .D(n_2763), .Q(GPR_21__1_) );
NAND2_Z01 g59834 ( .a(n_1206), .b(io_do_4), .o(n_1291) );
NAND2_Z01 g58753 ( .a(n_2204), .b(GPR_3__5_), .o(n_2347) );
BUF_X2 newInst_451 ( .a(newNet_207), .o(newNet_451) );
AND2_X1 g59166 ( .a(n_1036), .b(n_1880), .o(n_1936) );
BUF_X2 newInst_870 ( .a(newNet_869), .o(newNet_870) );
INV_X1 g61075 ( .a(pY_14_), .o(n_77) );
NAND2_Z01 g34539 ( .a(n_3925), .b(n_3913), .o(pmem_a_6) );
NAND2_Z01 g35393 ( .a(SP_5_), .b(SP_4_), .o(n_4535) );
AND2_X1 g60063 ( .a(n_845), .b(n_65), .o(n_1071) );
XOR2_X1 final_adder_mux_R16_278_6_g376 ( .a(final_adder_mux_R16_278_6_n_71), .b(final_adder_mux_R16_278_6_n_29), .o(R16_10_) );
AND2_X1 g58363 ( .a(n_2657), .b(n_2157), .o(n_2708) );
BUF_X2 newInst_83 ( .a(newNet_82), .o(newNet_83) );
NOR2_Z1 g60356 ( .a(n_604), .b(n_170), .o(n_852) );
fflopd GPR_reg_5__4_ ( .CK(newNet_853), .D(n_2927), .Q(GPR_5__4_) );
BUF_X2 newInst_752 ( .a(newNet_751), .o(newNet_752) );
NAND2_Z01 g60654 ( .a(n_332), .b(n_181), .o(n_488) );
NOR2_Z1 g59426 ( .a(n_1646), .b(n_1533), .o(n_1693) );
NAND2_Z01 g60556 ( .a(n_389), .b(n_405), .o(n_550) );
BUF_X2 newInst_1823 ( .a(newNet_1822), .o(newNet_1823) );
BUF_X2 newInst_259 ( .a(newNet_258), .o(newNet_259) );
NAND2_Z01 g59060 ( .a(n_1871), .b(n_4607), .o(n_2047) );
BUF_X2 newInst_568 ( .a(newNet_567), .o(newNet_568) );
NOR2_Z1 g60111 ( .a(n_849), .b(n_25), .o(n_1041) );
BUF_X2 newInst_1295 ( .a(newNet_1294), .o(newNet_1295) );
AND2_X1 g58262 ( .a(n_2752), .b(n_2208), .o(n_2805) );
INV_X1 g59962 ( .a(n_1164), .o(n_1165) );
AND3_X1 g60373 ( .a(n_4535), .b(n_609), .c(SP_6_), .o(n_770) );
NOR4_Z1 g34215 ( .a(n_4193), .b(n_4194), .c(n_4261), .d(n_4108), .o(n_4311) );
fflopd pZ_reg_2_ ( .CK(newNet_78), .D(n_2873), .Q(pZ_2_) );
BUF_X2 newInst_1613 ( .a(newNet_1612), .o(newNet_1613) );
NAND4_Z1 g60156 ( .a(n_674), .b(n_649), .c(n_694), .d(n_661), .o(n_979) );
NAND2_Z01 g58698 ( .a(n_2210), .b(GPR_1__5_), .o(n_2408) );
NAND2_Z01 g58760 ( .a(n_2203), .b(GPR_4__4_), .o(n_2340) );
NAND2_Z01 g58849 ( .a(n_2158), .b(GPR_12__2_), .o(n_2258) );
NAND2_Z01 g60448 ( .a(n_361), .b(GPR_7__1_), .o(n_698) );
INV_X1 drc_bufs61229 ( .a(n_7), .o(n_8) );
NAND2_Z01 g59294 ( .a(n_61), .b(n_1764), .o(n_1817) );
NAND2_Z01 g58715 ( .a(n_2208), .b(GPR_21__4_), .o(n_2392) );
NAND2_Z01 g60719 ( .a(GPR_5__1_), .b(n_183), .o(n_419) );
BUF_X2 newInst_1059 ( .a(newNet_1058), .o(newNet_1059) );
INV_X1 g60872 ( .a(n_257), .o(n_256) );
NAND2_Z02 g58968 ( .a(n_2088), .b(n_1211), .o(n_2140) );
BUF_X2 newInst_1267 ( .a(newNet_1266), .o(newNet_1267) );
NAND2_Z01 g60571 ( .a(n_466), .b(pX_3_), .o(n_613) );
BUF_X2 newInst_634 ( .a(newNet_633), .o(newNet_634) );
BUF_X2 newInst_598 ( .a(newNet_597), .o(newNet_598) );
NOR2_Z1 g34775 ( .a(n_3576), .b(n_4404), .o(n_3790) );
BUF_X2 newInst_975 ( .a(newNet_974), .o(newNet_975) );
BUF_X2 newInst_484 ( .a(newNet_483), .o(newNet_484) );
fflopd Rd_r_reg_2_ ( .CK(newNet_585), .D(n_948), .Q(Rd_r_2_) );
NAND2_Z01 g58060 ( .a(n_2884), .b(n_2306), .o(n_2922) );
AND2_X1 g59766 ( .a(n_1229), .b(pmem_d_1), .o(n_1360) );
BUF_X2 newInst_1492 ( .a(newNet_941), .o(newNet_1492) );
XOR2_X1 g35105 ( .a(n_4616), .b(n_3232), .o(n_4464) );
INV_X1 g59020 ( .a(n_2086), .o(n_2085) );
fflopd GPR_Rd_r_reg_0_ ( .CK(newNet_1863), .D(io_do_0), .Q(GPR_Rd_r_0_) );
NAND2_Z01 g57879 ( .a(n_3010), .b(n_2194), .o(n_3060) );
NAND2_Z01 g35216 ( .a(n_4523), .b(pY_11_), .o(n_4524) );
AND3_X1 g58607 ( .a(n_1999), .b(n_2462), .c(n_1998), .o(n_2504) );
BUF_X2 newInst_170 ( .a(newNet_169), .o(newNet_170) );
NOR2_Z1 g35204 ( .a(n_3414), .b(n_3264), .o(n_4532) );
BUF_X2 newInst_1654 ( .a(newNet_1653), .o(newNet_1654) );
NAND2_Z01 g34890 ( .a(n_3630), .b(pX_10_), .o(n_3673) );
BUF_X2 newInst_1731 ( .a(newNet_1730), .o(newNet_1731) );
BUF_X2 newInst_1723 ( .a(newNet_1722), .o(newNet_1723) );
NAND2_Z01 g60921 ( .a(C), .b(n_45), .o(n_261) );
NOR2_Z1 g59524 ( .a(n_1526), .b(n_1552), .o(n_1605) );
NAND2_Z01 g59327 ( .a(n_1699), .b(dmem_di_0), .o(n_1786) );
BUF_X2 newInst_879 ( .a(newNet_878), .o(newNet_879) );
NOR4_Z1 g58531 ( .a(n_1323), .b(n_2532), .c(n_1577), .d(n_1264), .o(n_2566) );
NAND4_Z1 g60130 ( .a(n_655), .b(n_727), .c(n_726), .d(n_556), .o(n_1002) );
NAND2_Z01 g60229 ( .a(n_750), .b(n_22), .o(n_916) );
XNOR2_X1 g60674 ( .a(n_280), .b(pY_2_), .o(n_475) );
NAND2_Z01 g58475 ( .a(n_2328), .b(n_2581), .o(n_2619) );
AND4_X1 g59493 ( .a(n_4625), .b(n_4470), .c(n_1523), .d(n_4627), .o(n_1634) );
NAND2_Z01 final_adder_mux_R16_278_6_g365 ( .a(final_adder_mux_R16_278_6_n_83), .b(final_adder_mux_R16_278_6_n_6), .o(final_adder_mux_R16_278_6_n_84) );
NOR2_Z1 g59741 ( .a(n_1298), .b(n_4419), .o(n_1381) );
NAND2_Z01 g57689 ( .a(n_3157), .b(n_2198), .o(n_3177) );
BUF_X2 newInst_332 ( .a(newNet_331), .o(newNet_332) );
NAND2_Z01 g60705 ( .a(n_198), .b(GPR_23__7_), .o(n_433) );
BUF_X2 newInst_1372 ( .a(newNet_1371), .o(newNet_1372) );
BUF_X2 newInst_1067 ( .a(newNet_1066), .o(newNet_1067) );
BUF_X2 newInst_743 ( .a(newNet_742), .o(newNet_743) );
NAND2_Z01 g34680 ( .a(n_3629), .b(GPR_3__7_), .o(n_3885) );
INV_X1 drc_bufs61230 ( .a(n_460), .o(n_7) );
AND2_X1 g60594 ( .a(n_4556), .b(n_469), .o(n_604) );
NAND3_Z1 g35090 ( .a(n_3434), .b(n_3459), .c(n_3259), .o(n_3501) );
NOR3_Z1 g34493 ( .a(n_3990), .b(n_4008), .c(n_4021), .o(n_4051) );
AND2_X1 g58253 ( .a(n_2752), .b(n_2157), .o(n_2814) );
INV_X1 g61101 ( .a(n_4523), .o(n_51) );
NAND2_Z01 g34278 ( .a(n_4162), .b(pY_9_), .o(n_4255) );
NAND2_Z01 g60477 ( .a(n_357), .b(pZ_9_), .o(n_669) );
NOR2_Z1 g34225 ( .a(n_4281), .b(n_4178), .o(n_4305) );
NOR2_Z1 g59015 ( .a(n_1980), .b(n_83), .o(n_2093) );
BUF_X2 newInst_697 ( .a(newNet_696), .o(newNet_697) );
BUF_X2 newInst_1363 ( .a(newNet_736), .o(newNet_1363) );
BUF_X2 newInst_1229 ( .a(newNet_518), .o(newNet_1229) );
NAND2_Z01 g34954 ( .a(n_3549), .b(GPR_17__2_), .o(n_3608) );
AND2_X1 g59887 ( .a(n_1207), .b(n_271), .o(n_1240) );
BUF_X2 newInst_954 ( .a(newNet_417), .o(newNet_954) );
NOR2_Z1 g34510 ( .a(n_4012), .b(n_3516), .o(n_4035) );
INV_X1 drc_bufs61121 ( .a(n_31), .o(n_19) );
NAND2_Z01 g57771 ( .a(n_3100), .b(n_2292), .o(n_3110) );
BUF_X2 newInst_105 ( .a(newNet_104), .o(newNet_105) );
NAND3_Z1 g59183 ( .a(S), .b(n_1826), .c(n_41), .o(n_1924) );
NAND2_Z01 g59680 ( .a(n_1378), .b(n_231), .o(n_1453) );
NAND2_Z01 g34612 ( .a(n_3900), .b(n_3489), .o(n_3948) );
NAND2_Z01 g57804 ( .a(n_3080), .b(n_2215), .o(n_3103) );
INV_X1 g61057 ( .a(pX_5_), .o(n_95) );
NAND2_Z01 g60723 ( .a(n_198), .b(GPR_20__4_), .o(n_415) );
BUF_X2 newInst_1105 ( .a(newNet_1104), .o(newNet_1105) );
BUF_X2 newInst_804 ( .a(newNet_803), .o(newNet_804) );
fflopd GPR_reg_3__7_ ( .CK(newNet_934), .D(n_3152), .Q(GPR_3__7_) );
INV_X1 g34560 ( .a(n_3976), .o(n_3999) );
XOR2_X1 g35075 ( .a(n_3471), .b(pZ_2_), .o(n_3515) );
NAND2_Z01 g60395 ( .a(n_433), .b(n_423), .o(n_751) );
NAND2_Z02 g58929 ( .a(n_2131), .b(n_1979), .o(n_2196) );
NAND2_Z01 g60835 ( .a(n_176), .b(n_59), .o(n_297) );
INV_X1 g34355 ( .a(n_4179), .o(n_4180) );
AND2_X1 g59774 ( .a(n_161), .b(io_sel_0_), .o(n_1355) );
fflopd T_reg ( .CK(newNet_450), .D(n_1659), .Q(T) );
NOR2_Z1 g60817 ( .a(n_199), .b(n_160), .o(n_353) );
NAND3_Z1 g35182 ( .a(n_3384), .b(n_3439), .c(n_3405), .o(n_4682) );
INV_X1 g61026 ( .a(pZ_4_), .o(n_126) );
NAND2_Z01 g60291 ( .a(n_596), .b(GPR_3__6_), .o(n_833) );
NAND4_Z1 g59843 ( .a(n_293), .b(n_781), .c(n_974), .d(n_462), .o(n_1283) );
BUF_X2 newInst_1568 ( .a(newNet_1567), .o(newNet_1568) );
BUF_X2 newInst_1214 ( .a(newNet_1213), .o(newNet_1214) );
NAND2_Z01 g59871 ( .a(n_837), .b(n_1170), .o(n_1256) );
NAND2_Z01 g60040 ( .a(n_856), .b(n_4607), .o(n_1090) );
BUF_X2 newInst_394 ( .a(newNet_393), .o(newNet_394) );
NAND2_Z01 g59723 ( .a(n_1345), .b(n_1170), .o(n_1404) );
BUF_X2 newInst_222 ( .a(newNet_221), .o(newNet_222) );
BUF_X2 newInst_777 ( .a(newNet_776), .o(newNet_777) );
NAND2_Z01 g58442 ( .a(n_2621), .b(n_2215), .o(n_2651) );
NAND2_Z01 g58778 ( .a(n_2201), .b(GPR_6__6_), .o(n_2322) );
AND2_X1 g59284 ( .a(n_1800), .b(n_274), .o(n_1824) );
NOR2_Z1 g60897 ( .a(n_91), .b(n_122), .o(n_235) );
NAND2_Z01 g60466 ( .a(n_368), .b(GPR_13__0_), .o(n_680) );
NAND2_Z01 g58557 ( .a(n_2510), .b(n_1711), .o(n_2550) );
BUF_X2 newInst_178 ( .a(newNet_177), .o(newNet_178) );
NAND4_Z1 g58347 ( .a(n_2078), .b(n_2499), .c(n_2653), .d(n_2026), .o(n_2723) );
NAND2_Z01 g34751 ( .a(n_3638), .b(n_3284), .o(n_3814) );
BUF_X2 newInst_164 ( .a(newNet_163), .o(newNet_164) );
NAND2_Z01 g34860 ( .a(n_3636), .b(GPR_10__0_), .o(n_3703) );
NAND2_Z01 g60418 ( .a(n_349), .b(U_6_), .o(n_728) );
fflopd pZ_reg_11_ ( .CK(newNet_102), .D(n_2955), .Q(pZ_11_) );
NAND2_Z01 g60249 ( .a(n_751), .b(n_22), .o(n_896) );
BUF_X2 newInst_1499 ( .a(newNet_1498), .o(newNet_1499) );
INV_X1 g35126 ( .a(n_3484), .o(n_3483) );
NAND2_Z01 g60692 ( .a(GPR_0__4_), .b(n_183), .o(n_446) );
AND3_X1 g59196 ( .a(n_1806), .b(n_1827), .c(pmem_d_7), .o(n_1913) );
AND2_X1 g57992 ( .a(n_2940), .b(n_2155), .o(n_2979) );
BUF_X2 newInst_521 ( .a(newNet_520), .o(newNet_521) );
BUF_X2 newInst_262 ( .a(newNet_261), .o(newNet_262) );
AND2_X1 g34415 ( .a(n_4063), .b(n_4088), .o(n_4122) );
NAND2_Z01 g34877 ( .a(n_3587), .b(GPR_2__7_), .o(n_3686) );
NAND2_Z01 g60316 ( .a(n_597), .b(pX_10_), .o(n_810) );
NAND2_Z01 g59132 ( .a(n_1872), .b(n_477), .o(n_1966) );
BUF_X2 newInst_1518 ( .a(newNet_1517), .o(newNet_1518) );
NAND3_Z1 g58827 ( .a(n_1721), .b(n_2135), .c(n_1753), .o(n_2280) );
NAND2_Z01 g59105 ( .a(n_1896), .b(n_1112), .o(n_2004) );
NAND2_Z01 g60219 ( .a(n_580), .b(GPR_14__3_), .o(n_926) );
INV_X1 g34440 ( .a(n_4610), .o(n_4098) );
fflopd U_reg_14_ ( .CK(newNet_404), .D(n_3111), .Q(U_14_) );
NAND2_Z01 g58582 ( .a(n_2464), .b(pY_4_), .o(n_2516) );
AND2_X1 g58505 ( .a(n_2567), .b(n_2211), .o(n_2592) );
AND2_X1 g59411 ( .a(io_do_1), .b(n_1664), .o(n_1707) );
INV_X1 g60537 ( .a(n_587), .o(n_586) );
BUF_X2 newInst_285 ( .a(newNet_284), .o(newNet_285) );
NAND2_Z01 final_adder_mux_R16_278_6_g392 ( .a(final_adder_mux_R16_278_6_n_56), .b(final_adder_mux_R16_278_6_n_13), .o(final_adder_mux_R16_278_6_n_57) );
NAND2_Z01 g35056 ( .a(n_3512), .b(PC_7_), .o(n_3527) );
BUF_X2 newInst_476 ( .a(newNet_475), .o(newNet_476) );
AND2_X1 g60805 ( .a(n_171), .b(PC_2_), .o(n_362) );
BUF_X2 newInst_98 ( .a(newNet_97), .o(newNet_98) );
BUF_X2 newInst_27 ( .a(newNet_18), .o(newNet_27) );
NAND2_Z01 g34733 ( .a(n_3631), .b(GPR_11__5_), .o(n_3832) );
NAND2_Z01 g57847 ( .a(n_3056), .b(n_904), .o(n_3079) );
NAND4_Z1 g59589 ( .a(n_1041), .b(n_1347), .c(n_1346), .d(V), .o(n_1539) );
BUF_X2 newInst_1740 ( .a(newNet_1739), .o(newNet_1740) );
NAND2_Z01 g34730 ( .a(n_3585), .b(GPR_12__5_), .o(n_3835) );
NOR4_Z1 g59303 ( .a(n_852), .b(n_1037), .c(n_1635), .d(n_566), .o(n_1811) );
NOR4_Z1 g34070 ( .a(n_4278), .b(n_4156), .c(n_4388), .d(n_4257), .o(n_4398) );
NAND2_Z01 g34111 ( .a(n_4334), .b(n_4349), .o(n_4431) );
NOR4_Z1 g34087 ( .a(n_4249), .b(n_4266), .c(n_4327), .d(n_4123), .o(n_4389) );
NOR3_Z1 g35251 ( .a(n_3231), .b(n_4482), .c(pmem_d_0), .o(n_3424) );
BUF_X2 newInst_1784 ( .a(newNet_1783), .o(newNet_1784) );
BUF_X2 newInst_136 ( .a(newNet_135), .o(newNet_136) );
AND2_X1 g59639 ( .a(n_1334), .b(n_1445), .o(n_1482) );
BUF_X2 newInst_1136 ( .a(newNet_1135), .o(newNet_1136) );
NAND2_Z01 g59679 ( .a(n_1385), .b(pmem_d_6), .o(n_1444) );
BUF_X2 newInst_327 ( .a(newNet_326), .o(newNet_327) );
NOR4_Z1 g58489 ( .a(n_2451), .b(n_2565), .c(n_2098), .d(n_1259), .o(n_2607) );
BUF_X2 newInst_1793 ( .a(newNet_1792), .o(newNet_1793) );
NAND2_Z01 g34150 ( .a(n_4317), .b(n_4614), .o(n_4358) );
NOR2_Z1 g60825 ( .a(n_160), .b(n_250), .o(n_349) );
NAND2_Z01 g59927 ( .a(n_1115), .b(n_127), .o(n_1190) );
NAND2_Z01 g34943 ( .a(n_3551), .b(GPR_4__2_), .o(n_3619) );
NAND2_Z01 g59086 ( .a(n_1871), .b(n_4608), .o(n_2021) );
AND2_X1 g59153 ( .a(n_1870), .b(n_4609), .o(n_1946) );
NAND2_Z01 final_adder_mux_R16_278_6_g423 ( .a(n_4448), .b(n_4432), .o(final_adder_mux_R16_278_6_n_25) );
NAND2_Z01 g60405 ( .a(Rd_0_), .b(n_345), .o(n_741) );
AND4_X1 g34597 ( .a(n_3423), .b(n_4665), .c(n_3569), .d(n_4666), .o(n_3963) );
fflopd GPR_reg_1__3_ ( .CK(newNet_1244), .D(n_2855), .Q(GPR_1__3_) );
fflopd pX_reg_2_ ( .CK(newNet_236), .D(n_2881), .Q(pX_2_) );
INV_X1 g35512 ( .a(PC_8_), .o(n_3216) );
NAND2_Z01 g35285 ( .a(n_3289), .b(pY_15_), .o(n_3390) );
INV_X1 g35022 ( .a(n_3553), .o(n_3552) );
BUF_X2 newInst_1358 ( .a(newNet_1357), .o(newNet_1358) );
INV_X1 g34935 ( .a(n_3626), .o(n_3627) );
BUF_X2 newInst_436 ( .a(newNet_435), .o(newNet_436) );
INV_X1 g35459 ( .a(pY_2_), .o(n_3265) );
BUF_X2 newInst_887 ( .a(newNet_886), .o(newNet_887) );
NAND2_Z01 g34684 ( .a(n_3625), .b(GPR_1__7_), .o(n_3881) );
NAND2_Z01 g35364 ( .a(n_3283), .b(n_3304), .o(n_3325) );
fflopd GPR_reg_0__0_ ( .CK(newNet_1816), .D(n_2617), .Q(GPR_0__0_) );
NAND2_Z01 g58719 ( .a(n_2207), .b(GPR_22__0_), .o(n_2388) );
BUF_X2 newInst_250 ( .a(newNet_249), .o(newNet_250) );
NAND2_Z01 g60697 ( .a(n_198), .b(GPR_23__6_), .o(n_441) );
BUF_X2 newInst_1590 ( .a(newNet_819), .o(newNet_1590) );
NAND3_Z1 g59518 ( .a(n_1444), .b(n_1522), .c(n_244), .o(n_1608) );
NOR3_Z1 g58941 ( .a(n_1849), .b(n_2101), .c(n_1937), .o(n_2166) );
AND2_X1 final_adder_mux_R16_278_6_g442 ( .a(n_4445), .b(n_4429), .o(final_adder_mux_R16_278_6_n_7) );
NOR2_Z1 g35413 ( .a(n_3254), .b(n_3233), .o(n_3292) );
NAND2_Z01 g58644 ( .a(n_2358), .b(pZ_5_), .o(n_2453) );
AND3_X1 g59038 ( .a(n_4524), .b(n_1983), .c(pY_12_), .o(n_2070) );
XNOR2_X1 g60597 ( .a(io_do_0), .b(n_261), .o(n_520) );
NAND2_Z01 g59264 ( .a(n_1802), .b(n_1728), .o(n_1846) );
BUF_X2 newInst_280 ( .a(newNet_279), .o(newNet_280) );
INV_X1 g59578 ( .a(n_1546), .o(n_1547) );
fflopd GPR_reg_20__6_ ( .CK(newNet_1178), .D(n_3076), .Q(GPR_20__6_) );
NAND2_Z01 g58765 ( .a(n_2202), .b(GPR_5__1_), .o(n_2335) );
NAND2_Z01 g59268 ( .a(n_1223), .b(n_1766), .o(n_1843) );
NAND2_Z01 g58837 ( .a(n_2159), .b(GPR_10__3_), .o(n_2270) );
NAND2_Z01 g59622 ( .a(n_1445), .b(T), .o(n_1505) );
NAND2_Z01 g60240 ( .a(R16_13_), .b(n_571), .o(n_905) );
NAND3_Z1 g58611 ( .a(n_1274), .b(n_2281), .c(n_1148), .o(n_2487) );
AND2_X1 g60108 ( .a(n_848), .b(n_135), .o(n_1015) );
NAND2_Z01 g58318 ( .a(n_2677), .b(n_2350), .o(n_2747) );
fflopd GPR_reg_23__2_ ( .CK(newNet_1049), .D(n_2758), .Q(GPR_23__2_) );
NAND2_Z01 g57840 ( .a(n_3036), .b(n_2338), .o(n_3070) );
NOR2_Z1 g60798 ( .a(n_272), .b(state_1_), .o(n_315) );
NAND2_Z01 g59702 ( .a(n_1353), .b(io_do_5), .o(n_1428) );
NAND2_Z01 g58842 ( .a(n_2139), .b(GPR_11__0_), .o(n_2265) );
BUF_X2 newInst_61 ( .a(newNet_60), .o(newNet_61) );
NAND2_Z01 g57936 ( .a(n_2971), .b(n_2391), .o(n_3006) );
NAND2_Z01 g35409 ( .a(pZ_5_), .b(pmem_d_13), .o(n_3303) );
NAND2_Z01 g60884 ( .a(pZ_0_), .b(pZ_1_), .o(n_278) );
NAND3_Z1 g60664 ( .a(n_336), .b(n_38), .c(n_163), .o(n_482) );
INV_X1 g35484 ( .a(pZ_8_), .o(n_3240) );
NAND2_Z01 g60518 ( .a(n_361), .b(GPR_5__3_), .o(n_628) );
fflopd U_reg_1_ ( .CK(newNet_392), .D(n_2868), .Q(U_1_) );
fflopd GPR_reg_0__7_ ( .CK(newNet_1771), .D(n_3170), .Q(GPR_0__7_) );
NAND2_Z01 g34906 ( .a(n_3590), .b(pY_8_), .o(n_3657) );
NAND2_Z01 g34540 ( .a(n_3924), .b(n_3912), .o(pmem_a_5) );
INV_X2 g35496 ( .a(pmem_d_1), .o(n_3231) );
NOR2_Z1 g60655 ( .a(n_459), .b(n_250), .o(n_570) );
AND2_X1 g59437 ( .a(n_1662), .b(SP_14_), .o(n_1697) );
BUF_X2 newInst_1094 ( .a(newNet_1093), .o(newNet_1094) );
NAND2_Z01 g60328 ( .a(n_25), .b(pmem_d_11), .o(n_800) );
NOR3_Z1 g60846 ( .a(state_1_), .b(n_4648), .c(state_0_), .o(n_292) );
INV_X1 drc_bufs35528 ( .a(n_4622), .o(n_3205) );
NAND2_Z01 g34994 ( .a(n_3544), .b(n_3262), .o(n_3588) );
BUF_X2 newInst_1013 ( .a(newNet_850), .o(newNet_1013) );
AND2_X1 g34549 ( .a(n_3917), .b(state_3_), .o(n_4646) );
NAND4_Z1 g57811 ( .a(n_1955), .b(n_2515), .c(n_3058), .d(n_2045), .o(n_3096) );
NOR2_Z1 g60337 ( .a(n_23), .b(n_44), .o(n_793) );
NAND2_Z01 g60266 ( .a(n_578), .b(GPR_19__0_), .o(n_880) );
NOR2_Z1 g34532 ( .a(n_3937), .b(state_3_), .o(n_4013) );
NOR2_Z1 g58448 ( .a(n_2605), .b(rst), .o(n_2645) );
AND2_X1 g60737 ( .a(n_98), .b(n_204), .o(n_402) );
BUF_X2 newInst_1271 ( .a(newNet_1270), .o(newNet_1271) );
NAND2_Z01 g58157 ( .a(n_2808), .b(n_2419), .o(n_2856) );
NAND2_Z01 g59920 ( .a(n_1113), .b(n_4522), .o(n_1220) );
XNOR2_X1 g58524 ( .a(n_2563), .b(n_1876), .o(n_2573) );
NAND4_Z1 g58546 ( .a(n_2276), .b(n_1607), .c(n_2150), .d(n_2490), .o(n_2552) );
BUF_X2 newInst_358 ( .a(newNet_357), .o(newNet_358) );
NAND2_Z01 g60462 ( .a(n_353), .b(GPR_8__0_), .o(n_684) );
INV_Z1 g35493 ( .a(pZ_0_), .o(n_4635) );
BUF_X2 newInst_1809 ( .a(newNet_1808), .o(newNet_1809) );
AND2_X1 g58113 ( .a(n_2850), .b(n_2211), .o(n_2899) );
BUF_X2 newInst_547 ( .a(newNet_546), .o(newNet_547) );
NAND3_Z1 g59491 ( .a(n_1436), .b(n_1610), .c(n_1560), .o(n_1636) );
NOR2_Z1 g60054 ( .a(n_858), .b(n_90), .o(n_1080) );
NAND2_Z01 g34753 ( .a(n_3567), .b(GPR_6__4_), .o(n_3812) );
BUF_X2 newInst_442 ( .a(newNet_441), .o(newNet_442) );
NAND2_Z01 g57938 ( .a(n_2969), .b(n_2375), .o(n_3004) );
BUF_X2 newInst_447 ( .a(newNet_446), .o(newNet_447) );
NAND2_Z01 g34858 ( .a(n_3566), .b(GPR_18__0_), .o(n_3705) );
NAND2_Z01 g58034 ( .a(n_2913), .b(n_2302), .o(n_2951) );
NAND2_Z01 g58098 ( .a(n_2852), .b(n_2215), .o(n_2915) );
AND2_X1 g57750 ( .a(n_3115), .b(n_2201), .o(n_3121) );
BUF_X2 newInst_458 ( .a(newNet_457), .o(newNet_458) );
NOR2_Z1 g34310 ( .a(n_4612), .b(n_3534), .o(n_4223) );
INV_X1 g35476 ( .a(pmem_d_11), .o(n_3248) );
INV_X1 g61079 ( .a(SP_12_), .o(n_73) );
NOR2_Z1 g35356 ( .a(n_4482), .b(n_4490), .o(n_4662) );
NAND2_Z01 g59605 ( .a(n_1413), .b(io_sp_2_), .o(n_1521) );
NAND2_Z01 g34402 ( .a(n_3208), .b(pZ_2_), .o(n_4136) );
NAND2_Z01 g60974 ( .a(n_121), .b(n_65), .o(n_194) );
NOR2_Z1 g60606 ( .a(n_458), .b(n_182), .o(n_596) );
NAND2_Z01 g34094 ( .a(n_4375), .b(n_4374), .o(n_4436) );
AND2_X1 g35309 ( .a(n_3256), .b(n_3309), .o(n_3367) );
BUF_X2 newInst_425 ( .a(newNet_395), .o(newNet_425) );
NAND2_Z01 g57945 ( .a(n_2962), .b(n_2228), .o(n_2997) );
BUF_X2 newInst_1133 ( .a(newNet_1132), .o(newNet_1133) );
INV_X1 g34797 ( .a(n_3766), .o(n_4565) );
INV_X1 g59208 ( .a(n_1902), .o(n_1901) );
BUF_X2 newInst_1144 ( .a(newNet_1143), .o(newNet_1144) );
XOR2_X1 g59906 ( .a(n_1115), .b(PC_3_), .o(n_1225) );
NAND2_Z01 g34838 ( .a(n_3635), .b(GPR_14__1_), .o(n_3725) );
NAND2_Z01 g60330 ( .a(n_11), .b(pmem_d_8), .o(n_798) );
XOR2_X1 g34501 ( .a(n_4026), .b(pY_7_), .o(n_4043) );
NAND2_Z01 g59610 ( .a(n_1453), .b(n_146), .o(n_1517) );
BUF_X2 newInst_1165 ( .a(newNet_1164), .o(newNet_1165) );
NAND2_Z01 g60035 ( .a(n_766), .b(n_247), .o(n_1095) );
NAND2_Z01 g59027 ( .a(n_2061), .b(n_962), .o(n_2089) );
NAND2_Z01 g59334 ( .a(n_1714), .b(n_1252), .o(n_1780) );
NAND2_Z01 g34784 ( .a(n_3567), .b(GPR_6__3_), .o(n_3781) );
fflopd GPR_reg_8__0_ ( .CK(newNet_729), .D(n_2616), .Q(GPR_8__0_) );
BUF_X2 newInst_1846 ( .a(newNet_1845), .o(newNet_1846) );
AND2_X1 g58818 ( .a(n_2215), .b(n_2058), .o(n_2359) );
BUF_X2 newInst_724 ( .a(newNet_489), .o(newNet_724) );
BUF_X2 newInst_152 ( .a(newNet_107), .o(newNet_152) );
XOR2_X1 final_adder_mux_R16_278_6_g410 ( .a(n_4447), .b(n_4431), .o(final_adder_mux_R16_278_6_n_39) );
XOR2_X1 g34929 ( .a(n_3545), .b(pY_9_), .o(n_3765) );
BUF_X2 newInst_1675 ( .a(newNet_1674), .o(newNet_1675) );
NAND3_Z1 g60100 ( .a(n_4532), .b(n_567), .c(SP_12_), .o(n_1049) );
BUF_X2 newInst_1081 ( .a(newNet_1080), .o(newNet_1081) );
NOR2_Z1 g34182 ( .a(n_4324), .b(n_4617), .o(n_4422) );
INV_X1 drc_bufs61165 ( .a(n_579), .o(n_25) );
NAND2_Z01 g35292 ( .a(n_3299), .b(pX_12_), .o(n_3383) );
BUF_X2 newInst_539 ( .a(newNet_74), .o(newNet_539) );
NAND4_Z1 g34574 ( .a(n_3818), .b(n_3815), .c(n_3817), .d(n_3816), .o(n_3986) );
XOR2_X1 g34438 ( .a(n_4076), .b(SP_3_), .o(n_4101) );
NAND4_Z1 g58143 ( .a(n_1967), .b(n_2498), .c(n_2818), .d(n_2019), .o(n_2870) );
NAND2_Z01 g58462 ( .a(n_2596), .b(n_2245), .o(n_2634) );
INV_X1 g61087 ( .a(pmem_d_8), .o(n_65) );
NOR2_Z1 g60785 ( .a(n_202), .b(n_182), .o(n_380) );
NAND2_Z01 g34790 ( .a(n_3628), .b(GPR_19__3_), .o(n_3775) );
fflopd SP_reg_13_ ( .CK(newNet_543), .D(n_1858), .Q(SP_13_) );
BUF_X2 newInst_1574 ( .a(newNet_1573), .o(newNet_1574) );
BUF_X2 newInst_1558 ( .a(newNet_1557), .o(newNet_1558) );
BUF_X2 newInst_1685 ( .a(newNet_1684), .o(newNet_1685) );
AND2_X1 g35166 ( .a(n_4639), .b(n_4558), .o(n_4583) );
BUF_X2 newInst_54 ( .a(newNet_53), .o(newNet_54) );
INV_X1 g61109 ( .a(pmem_d_11), .o(n_43) );
NAND2_Z01 g34178 ( .a(n_4325), .b(n_4473), .o(n_4338) );
NAND2_Z01 g60711 ( .a(n_178), .b(n_4535), .o(n_427) );
XOR2_X1 final_adder_mux_R16_278_6_g414 ( .a(n_4451), .b(n_4435), .o(R16_0_) );
fflopd io_sp_reg_6_ ( .CK(newNet_304), .D(n_552), .Q(io_sp_6_) );
BUF_X2 newInst_1852 ( .a(newNet_1851), .o(newNet_1852) );
BUF_X2 newInst_1521 ( .a(newNet_1520), .o(newNet_1521) );
BUF_X2 newInst_1451 ( .a(newNet_1450), .o(newNet_1451) );
NAND2_Z01 g58044 ( .a(n_2901), .b(n_2406), .o(n_2938) );
BUF_X2 newInst_951 ( .a(newNet_950), .o(newNet_951) );
NAND4_Z1 g34247 ( .a(n_3676), .b(n_3725), .c(n_4174), .d(n_3724), .o(n_4286) );
BUF_X2 newInst_1241 ( .a(newNet_1240), .o(newNet_1241) );
BUF_X2 newInst_382 ( .a(newNet_381), .o(newNet_382) );
INV_X1 g61080 ( .a(n_4527), .o(n_72) );
BUF_X2 newInst_373 ( .a(newNet_372), .o(newNet_373) );
NOR2_Z1 g59716 ( .a(n_1308), .b(n_1388), .o(n_1418) );
NAND2_Z01 g60274 ( .a(R16_14_), .b(n_14), .o(n_872) );
NAND2_Z01 g58637 ( .a(n_2361), .b(n_2006), .o(n_2465) );
INV_X2 newInst_1033 ( .a(newNet_1032), .o(newNet_1033) );
NAND2_Z01 g60643 ( .a(n_287), .b(n_255), .o(n_495) );
NAND2_Z01 g58621 ( .a(n_2360), .b(pY_1_), .o(n_2476) );
AND3_X1 g60151 ( .a(state_2_), .b(n_498), .c(state_3_), .o(n_1027) );
BUF_X2 newInst_1753 ( .a(newNet_1752), .o(newNet_1753) );
NAND2_Z01 g60940 ( .a(n_61), .b(pmem_d_10), .o(n_211) );
NOR2_Z1 g34622 ( .a(n_3675), .b(n_3650), .o(n_3938) );
NAND2_Z01 g58799 ( .a(n_2195), .b(U_12_), .o(n_2301) );
NAND2_Z01 g60048 ( .a(n_792), .b(n_823), .o(n_1083) );
NOR2_Z1 g34344 ( .a(n_16064_BAR), .b(n_3762), .o(n_4190) );
AND2_X1 g60803 ( .a(n_177), .b(n_4532), .o(n_313) );
NOR4_Z1 g59795 ( .a(n_991), .b(n_983), .c(n_1150), .d(n_955), .o(n_1329) );
NOR2_Z1 g35009 ( .a(n_4650), .b(n_3429), .o(n_3559) );
NAND2_Z01 g59822 ( .a(n_1171), .b(dmem_di_1), .o(n_1302) );
NAND2_Z01 g59690 ( .a(n_1326), .b(io_do_0), .o(n_1439) );
BUF_X2 newInst_806 ( .a(newNet_521), .o(newNet_806) );
INV_X1 g61065 ( .a(PC_2_), .o(n_87) );
NAND2_Z01 g57841 ( .a(n_3035), .b(n_2330), .o(n_3069) );
NAND2_Z01 g60324 ( .a(n_577), .b(pZ_13_), .o(n_803) );
BUF_X2 newInst_1547 ( .a(newNet_1546), .o(newNet_1547) );
INV_Z1 g35508 ( .a(PC_0_), .o(n_4555) );
INV_X1 g60776 ( .a(n_344), .o(n_343) );
NAND2_Z01 g60211 ( .a(n_582), .b(GPR_11__7_), .o(n_934) );
NAND4_Z1 g59992 ( .a(n_922), .b(n_927), .c(n_943), .d(n_806), .o(n_1137) );
NOR2_Z1 g34967 ( .a(n_3553), .b(n_3492), .o(n_3631) );
INV_X2 newInst_845 ( .a(newNet_844), .o(newNet_845) );
BUF_X2 newInst_813 ( .a(newNet_812), .o(newNet_813) );
NAND4_Z1 g58935 ( .a(n_1689), .b(n_1792), .c(n_2120), .d(n_1641), .o(n_2172) );
NAND2_Z01 g60521 ( .a(n_353), .b(GPR_8__7_), .o(n_625) );
fflopd GPR_reg_7__2_ ( .CK(newNet_771), .D(n_2739), .Q(GPR_7__2_) );
INV_X1 g59860 ( .a(n_1270), .o(n_1271) );
NOR2_Z4 g58450 ( .a(n_2608), .b(n_1589), .o(n_2657) );
AND2_X1 g60060 ( .a(n_845), .b(n_43), .o(n_1074) );
NOR2_Z1 g58964 ( .a(n_2116), .b(n_965), .o(n_2154) );
NOR2_Z1 g60348 ( .a(n_514), .b(n_503), .o(n_783) );
NAND2_Z01 g58310 ( .a(n_2683), .b(n_2386), .o(n_2760) );
BUF_X2 newInst_1479 ( .a(newNet_1478), .o(newNet_1479) );
fflopd io_sp_reg_0_ ( .CK(newNet_335), .D(n_547), .Q(io_sp_0_) );
BUF_X2 newInst_1141 ( .a(newNet_1140), .o(newNet_1141) );
BUF_X2 newInst_73 ( .a(newNet_72), .o(newNet_73) );
NAND2_Z01 g34949 ( .a(n_3551), .b(GPR_14__5_), .o(n_3613) );
NAND2_Z01 g58776 ( .a(n_2201), .b(GPR_6__4_), .o(n_2324) );
BUF_X2 newInst_903 ( .a(newNet_902), .o(newNet_903) );
NAND2_Z01 g60938 ( .a(n_64), .b(pmem_d_8), .o(n_213) );
NAND2_Z01 g58144 ( .a(n_2822), .b(n_2303), .o(n_2869) );
NAND2_Z01 g34648 ( .a(n_3768), .b(n_4545), .o(n_3912) );
BUF_X2 newInst_1201 ( .a(newNet_446), .o(newNet_1201) );
NAND2_Z01 g34773 ( .a(n_3597), .b(GPR_17__4_), .o(n_3792) );
NAND2_Z01 g59077 ( .a(n_1871), .b(n_4604), .o(n_2030) );
NAND2_Z01 g59619 ( .a(n_1414), .b(io_di_4), .o(n_1508) );
BUF_X2 newInst_1189 ( .a(newNet_1188), .o(newNet_1189) );
NAND2_Z01 g34908 ( .a(n_3590), .b(pY_10_), .o(n_3655) );
NAND2_Z01 g59394 ( .a(n_1197), .b(n_1663), .o(n_1721) );
NAND2_Z01 g34521 ( .a(n_3850), .b(n_3947), .o(n_4022) );
BUF_X2 newInst_494 ( .a(newNet_493), .o(newNet_494) );
BUF_X2 newInst_431 ( .a(newNet_101), .o(newNet_431) );
NAND2_Z01 g60053 ( .a(n_865), .b(pX_5_), .o(n_1111) );
BUF_X2 newInst_1309 ( .a(newNet_1308), .o(newNet_1309) );
NAND3_Z1 g59489 ( .a(n_1399), .b(n_1554), .c(n_909), .o(n_1637) );
BUF_X2 newInst_1202 ( .a(newNet_1201), .o(newNet_1202) );
fflopd GPR_reg_5__3_ ( .CK(newNet_859), .D(n_2843), .Q(GPR_5__3_) );
NAND2_Z01 g34110 ( .a(n_4339), .b(n_4352), .o(n_4447) );
AND2_X1 g59367 ( .a(n_1694), .b(n_850), .o(n_1747) );
BUF_X2 newInst_1348 ( .a(newNet_1347), .o(newNet_1348) );
BUF_X2 newInst_12 ( .a(newNet_11), .o(newNet_12) );
AND2_X1 g58255 ( .a(n_2752), .b(n_2156), .o(n_2812) );
AND4_X1 g58937 ( .a(n_1755), .b(n_1860), .c(n_2097), .d(n_1640), .o(n_2170) );
NAND2_Z01 g59387 ( .a(n_1667), .b(PC_7_), .o(n_1728) );
NAND2_Z01 g58850 ( .a(n_2158), .b(GPR_12__3_), .o(n_2257) );
NAND2_Z01 g58901 ( .a(n_2162), .b(n_1772), .o(n_2181) );
BUF_X2 newInst_1698 ( .a(newNet_1697), .o(newNet_1698) );
NAND2_Z01 final_adder_mux_R16_278_6_g393 ( .a(final_adder_mux_R16_278_6_n_54), .b(final_adder_mux_R16_278_6_n_26), .o(final_adder_mux_R16_278_6_n_56) );
NOR2_Z1 g61014 ( .a(n_4657), .b(state_1_), .o(n_130) );
NAND2_Z01 g34688 ( .a(n_3594), .b(GPR_7__7_), .o(n_3877) );
BUF_X2 newInst_1099 ( .a(newNet_1098), .o(newNet_1099) );
BUF_X2 newInst_317 ( .a(newNet_316), .o(newNet_317) );
NAND2_Z01 g58807 ( .a(n_2197), .b(U_5_), .o(n_2293) );
BUF_X2 newInst_260 ( .a(newNet_259), .o(newNet_260) );
BUF_X2 newInst_111 ( .a(newNet_11), .o(newNet_111) );
BUF_X2 newInst_49 ( .a(newNet_48), .o(newNet_49) );
NOR2_Z1 g35313 ( .a(n_3235), .b(n_3288), .o(n_3364) );
NAND2_Z01 g58896 ( .a(n_2156), .b(GPR_15__7_), .o(n_2186) );
BUF_X2 newInst_1182 ( .a(newNet_1181), .o(newNet_1182) );
fflopd io_sel_reg_0_ ( .CK(newNet_342), .D(n_1144), .Q(io_sel_0_) );
NAND4_Z1 g34568 ( .a(n_3851), .b(n_3854), .c(n_3853), .d(n_3852), .o(n_3992) );
NAND2_Z01 g60732 ( .a(n_178), .b(n_275), .o(n_407) );
NAND2_Z01 g34160 ( .a(n_4317), .b(pmem_d_7), .o(n_4348) );
BUF_X2 newInst_1504 ( .a(newNet_1503), .o(newNet_1504) );
NAND2_Z01 g35206 ( .a(n_3415), .b(PC_3_), .o(n_3452) );
INV_X1 g61039 ( .a(pY_6_), .o(n_113) );
AND2_X1 g60345 ( .a(n_613), .b(pX_4_), .o(n_786) );
NAND2_Z01 g58735 ( .a(n_2205), .b(GPR_2__0_), .o(n_2372) );
NAND2_Z01 g60568 ( .a(n_357), .b(pY_8_), .o(n_541) );
NAND2_Z01 g58336 ( .a(n_827), .b(n_2689), .o(n_2753) );
NOR4_Z1 g59538 ( .a(n_307), .b(n_1231), .c(n_1548), .d(n_215), .o(n_1601) );
AND2_X1 g59945 ( .a(n_1111), .b(pX_6_), .o(n_1181) );
NAND2_Z01 g60298 ( .a(n_580), .b(GPR_14__7_), .o(n_826) );
NAND2_Z01 g58685 ( .a(n_2211), .b(GPR_19__1_), .o(n_2421) );
BUF_X2 newInst_97 ( .a(newNet_96), .o(newNet_97) );
NAND2_Z01 g58284 ( .a(n_2714), .b(n_2271), .o(n_2786) );
INV_X1 drc_bufs61202 ( .a(n_2193), .o(n_12) );
BUF_X2 newInst_306 ( .a(newNet_305), .o(newNet_306) );
NAND2_Z01 g60315 ( .a(n_570), .b(pZ_3_), .o(n_811) );
NAND2_Z01 g34846 ( .a(n_3631), .b(GPR_11__1_), .o(n_3717) );
NAND4_Z1 g58017 ( .a(n_2068), .b(n_2543), .c(n_2918), .d(n_2034), .o(n_2955) );
NAND2_Z03 g34226 ( .a(n_4288), .b(n_3999), .o(io_do_2) );
BUF_X2 newInst_524 ( .a(newNet_523), .o(newNet_524) );
NOR2_Z1 g35011 ( .a(n_3510), .b(n_3548), .o(n_3566) );
BUF_X2 newInst_1500 ( .a(newNet_1499), .o(newNet_1500) );
NAND2_Z01 g57659 ( .a(n_3177), .b(n_2291), .o(n_3183) );
BUF_X2 newInst_1230 ( .a(newNet_1229), .o(newNet_1230) );
BUF_X2 newInst_1439 ( .a(newNet_1438), .o(newNet_1439) );
NAND2_Z01 g59222 ( .a(n_1853), .b(n_25), .o(n_1884) );
NAND3_Z1 g59892 ( .a(io_do_6), .b(n_1026), .c(n_459), .o(n_1237) );
NOR2_Z1 g34255 ( .a(n_4175), .b(n_3241), .o(n_4278) );
NAND3_Z1 g60849 ( .a(n_52), .b(n_47), .c(n_48), .o(n_337) );
BUF_X2 newInst_59 ( .a(newNet_58), .o(newNet_59) );
AND2_X1 g58114 ( .a(n_2850), .b(n_2210), .o(n_2898) );
NAND4_Z1 g59256 ( .a(n_1183), .b(n_1751), .c(n_1555), .d(n_791), .o(n_1856) );
BUF_X2 newInst_69 ( .a(newNet_68), .o(newNet_69) );
AND2_X1 g34989 ( .a(n_3545), .b(pY_9_), .o(n_3593) );
fflopd io_sp_reg_7_ ( .CK(newNet_296), .D(n_745), .Q(io_sp_7_) );
AND2_X1 g59476 ( .a(n_1595), .b(n_1128), .o(n_1661) );
BUF_X2 newInst_424 ( .a(newNet_423), .o(newNet_424) );
NOR2_Z1 g35079 ( .a(n_3493), .b(n_3221), .o(n_3512) );
NAND2_Z01 g58703 ( .a(n_2209), .b(GPR_20__0_), .o(n_2404) );
NAND2_Z01 final_adder_mux_R16_278_6_g398 ( .a(final_adder_mux_R16_278_6_n_50), .b(final_adder_mux_R16_278_6_n_9), .o(final_adder_mux_R16_278_6_n_51) );
NAND2_Z01 g60334 ( .a(n_566), .b(pmem_d_10), .o(n_795) );
NAND2_Z01 g59466 ( .a(n_1627), .b(n_154), .o(n_1657) );
BUF_X2 newInst_860 ( .a(newNet_523), .o(newNet_860) );
BUF_X2 newInst_778 ( .a(newNet_777), .o(newNet_778) );
NAND2_Z01 g60189 ( .a(n_659), .b(n_660), .o(n_963) );
NAND2_Z01 g35001 ( .a(n_3509), .b(n_3551), .o(n_3580) );
NOR2_Z1 g59469 ( .a(n_1626), .b(n_106), .o(n_1665) );
BUF_X2 newInst_984 ( .a(newNet_853), .o(newNet_984) );
BUF_X2 newInst_771 ( .a(newNet_312), .o(newNet_771) );
INV_X2 g61120 ( .a(pmem_d_13), .o(n_32) );
BUF_X2 newInst_841 ( .a(newNet_840), .o(newNet_841) );
AND3_X1 g59771 ( .a(pmem_d_8), .b(n_1129), .c(pmem_d_7), .o(n_1383) );
BUF_X2 newInst_686 ( .a(newNet_685), .o(newNet_686) );
NAND2_Z01 g57877 ( .a(n_3011), .b(n_2217), .o(n_3062) );
BUF_X2 newInst_1835 ( .a(newNet_1834), .o(newNet_1835) );
NAND3_Z1 g60364 ( .a(n_434), .b(n_413), .c(n_446), .o(n_776) );
NOR2_Z1 g59011 ( .a(n_1981), .b(n_91), .o(n_2097) );
BUF_X2 newInst_1666 ( .a(newNet_1665), .o(newNet_1666) );
INV_X1 g34979 ( .a(n_3576), .o(n_3575) );
AND3_X1 g59656 ( .a(n_994), .b(n_1324), .c(n_957), .o(n_1470) );
INV_X1 g59777 ( .a(n_1351), .o(n_1352) );
NAND2_Z01 g60824 ( .a(n_185), .b(n_263), .o(n_304) );
BUF_X2 newInst_1208 ( .a(newNet_1207), .o(newNet_1208) );
BUF_X2 newInst_1088 ( .a(newNet_1087), .o(newNet_1088) );
INV_X2 newInst_986 ( .a(newNet_985), .o(newNet_986) );
NAND2_Z01 g58756 ( .a(n_2203), .b(GPR_4__0_), .o(n_2344) );
NAND2_Z01 g59632 ( .a(n_17), .b(C), .o(n_1497) );
BUF_X2 newInst_947 ( .a(newNet_96), .o(newNet_947) );
BUF_X2 newInst_867 ( .a(newNet_866), .o(newNet_867) );
NAND2_Z01 g35282 ( .a(U_10_), .b(n_3275), .o(n_3393) );
NOR2_Z1 g34788 ( .a(n_3626), .b(n_4408), .o(n_3777) );
BUF_X2 newInst_1645 ( .a(newNet_1644), .o(newNet_1645) );
NOR2_Z1 g35114 ( .a(n_3204), .b(pmem_d_6), .o(n_4471) );
NAND2_Z01 g60218 ( .a(n_585), .b(GPR_23__3_), .o(n_927) );
NAND2_Z01 g60903 ( .a(state_1_), .b(state_3_), .o(n_268) );
NAND2_Z01 g59762 ( .a(n_1268), .b(n_1161), .o(n_1363) );
fflopd GPR_reg_1__0_ ( .CK(newNet_1267), .D(n_2630), .Q(GPR_1__0_) );
INV_X1 g35467 ( .a(PC_2_), .o(n_3257) );
NOR2_Z1 g59357 ( .a(n_19), .b(n_1394), .o(n_1756) );
NAND2_Z01 g34823 ( .a(n_3585), .b(GPR_13__2_), .o(n_3740) );
NAND4_Z1 g58119 ( .a(n_1545), .b(n_2124), .c(n_2757), .d(n_1538), .o(n_2893) );
BUF_X2 newInst_135 ( .a(newNet_134), .o(newNet_135) );
NAND2_Z01 g34608 ( .a(n_3713), .b(n_3652), .o(n_3952) );
AND3_X1 g59191 ( .a(n_1390), .b(n_1873), .c(pX_9_), .o(n_1916) );
BUF_X2 newInst_64 ( .a(newNet_45), .o(newNet_64) );
NAND2_Z01 g60268 ( .a(n_582), .b(GPR_11__5_), .o(n_878) );
NAND2_Z01 g59484 ( .a(n_27), .b(n_1227), .o(n_1641) );
BUF_X2 newInst_1026 ( .a(newNet_1025), .o(newNet_1026) );
BUF_X2 newInst_604 ( .a(newNet_603), .o(newNet_604) );
BUF_X2 newInst_738 ( .a(newNet_737), .o(newNet_738) );
fflopd GPR_reg_11__1_ ( .CK(newNet_1702), .D(n_2784), .Q(GPR_11__1_) );
NAND2_Z01 g57926 ( .a(n_2981), .b(n_2255), .o(n_3019) );
BUF_X2 newInst_1842 ( .a(newNet_1841), .o(newNet_1842) );
NAND2_Z01 g60070 ( .a(io_do_3), .b(n_841), .o(n_1064) );
BUF_X2 newInst_1256 ( .a(newNet_1255), .o(newNet_1256) );
NAND2_Z02 g34378 ( .a(n_4643), .b(n_4093), .o(n_4613) );
NOR2_Z1 g59163 ( .a(n_1890), .b(n_1688), .o(n_1981) );
NAND2_Z01 g34189 ( .a(n_4325), .b(n_4465), .o(n_4334) );
BUF_X2 newInst_1329 ( .a(newNet_1328), .o(newNet_1329) );
NAND2_Z01 g60259 ( .a(n_590), .b(GPR_6__5_), .o(n_887) );
NAND2_Z01 g58539 ( .a(n_2550), .b(n_1940), .o(n_2559) );
NAND2_Z01 g60194 ( .a(n_637), .b(n_619), .o(n_951) );
XNOR2_X1 g60869 ( .a(n_4446), .b(n_4430), .o(n_325) );
AND2_X1 g57749 ( .a(n_3115), .b(n_2202), .o(n_3122) );
BUF_X2 newInst_1534 ( .a(newNet_1533), .o(newNet_1534) );
BUF_X2 newInst_1463 ( .a(newNet_1462), .o(newNet_1463) );
NAND2_Z01 g60458 ( .a(n_358), .b(GPR_0__0_), .o(n_688) );
NOR2_Z1 g35272 ( .a(n_4534), .b(n_3246), .o(n_4531) );
BUF_X2 newInst_768 ( .a(newNet_767), .o(newNet_768) );
AND2_X1 g59343 ( .a(io_do_3), .b(n_15), .o(n_1774) );
NAND2_Z01 g59882 ( .a(n_1164), .b(n_55), .o(n_1245) );
NOR3_Z1 g34655 ( .a(n_3601), .b(n_4650), .c(n_4637), .o(n_3905) );
NAND2_Z01 g59785 ( .a(n_1268), .b(n_359), .o(n_1339) );
NAND4_Z1 g57656 ( .a(n_1987), .b(n_2519), .c(n_3180), .d(n_2037), .o(n_3186) );
NAND2_Z01 g35041 ( .a(n_4515), .b(n_4516), .o(n_3539) );
NOR2_Z1 g60991 ( .a(rst), .b(pmem_d_0), .o(n_180) );
NOR2_Z1 g34269 ( .a(n_4613), .b(n_3214), .o(n_4264) );
NOR4_Z1 g34214 ( .a(n_4207), .b(n_4264), .c(n_4206), .d(n_4112), .o(n_4312) );
INV_X1 g35318 ( .a(n_3359), .o(n_3358) );
NAND2_Z01 g34395 ( .a(n_4599), .b(n_4098), .o(n_4143) );
BUF_X2 newInst_50 ( .a(newNet_49), .o(newNet_50) );
NOR2_Z1 g60049 ( .a(n_964), .b(n_26), .o(n_1082) );
NAND2_Z01 g34868 ( .a(n_3594), .b(GPR_7__0_), .o(n_3695) );
NAND2_Z01 final_adder_mux_R16_278_6_g386 ( .a(final_adder_mux_R16_278_6_n_62), .b(final_adder_mux_R16_278_6_n_11), .o(final_adder_mux_R16_278_6_n_63) );
NAND2_Z01 g34708 ( .a(n_3633), .b(pZ_14_), .o(n_3857) );
BUF_X2 newInst_552 ( .a(newNet_551), .o(newNet_552) );
INV_X1 g35203 ( .a(n_3443), .o(n_3444) );
XOR2_X1 final_adder_mux_R16_278_6_g406 ( .a(n_4443), .b(n_4427), .o(final_adder_mux_R16_278_6_n_43) );
NAND2_Z01 g60429 ( .a(n_349), .b(U_2_), .o(n_717) );
AND2_X1 g57887 ( .a(n_3009), .b(n_2158), .o(n_3051) );
NAND2_Z01 g58676 ( .a(n_2213), .b(GPR_17__7_), .o(n_2430) );
NAND4_Z1 g59036 ( .a(n_24), .b(n_1169), .c(n_1811), .d(n_587), .o(n_2072) );
BUF_X2 newInst_1715 ( .a(newNet_1714), .o(newNet_1715) );
BUF_X2 newInst_121 ( .a(newNet_120), .o(newNet_121) );
BUF_X2 newInst_1595 ( .a(newNet_539), .o(newNet_1595) );
NAND3_Z1 g57651 ( .a(n_2561), .b(n_3174), .c(n_2146), .o(n_3191) );
NAND2_Z01 g60681 ( .a(GPR_5__4_), .b(n_183), .o(n_456) );
NOR2_Z1 g59119 ( .a(n_1867), .b(n_48), .o(n_2059) );
NAND4_Z1 g34563 ( .a(n_3878), .b(n_3881), .c(n_3880), .d(n_3879), .o(n_3997) );
NAND2_Z01 g60501 ( .a(n_53), .b(n_410), .o(n_645) );
fflopd GPR_reg_21__3_ ( .CK(newNet_1141), .D(n_2853), .Q(GPR_21__3_) );
BUF_X2 newInst_654 ( .a(newNet_653), .o(newNet_654) );
NAND2_Z01 g58248 ( .a(n_2753), .b(n_2196), .o(n_2819) );
BUF_X2 newInst_1350 ( .a(newNet_1349), .o(newNet_1350) );
NOR3_Z1 g35070 ( .a(n_3433), .b(n_3486), .c(n_3424), .o(n_3517) );
NAND2_Z01 g58587 ( .a(n_2478), .b(pY_8_), .o(n_2511) );
BUF_X2 newInst_1710 ( .a(newNet_1709), .o(newNet_1710) );
NAND2_Z01 g60067 ( .a(n_841), .b(io_do_1), .o(n_1067) );
XNOR2_X1 g58547 ( .a(n_2526), .b(n_2087), .o(n_2551) );
NAND2_Z01 g59068 ( .a(n_1896), .b(n_4609), .o(n_2039) );
NAND2_Z01 g59519 ( .a(n_1276), .b(n_1546), .o(n_1607) );
fflopd GPR_reg_12__6_ ( .CK(newNet_1621), .D(n_3088), .Q(GPR_12__6_) );
NAND2_Z01 g60208 ( .a(n_591), .b(GPR_22__6_), .o(n_937) );
XOR2_X1 g59381 ( .a(n_1669), .b(n_318), .o(n_1737) );
NAND2_Z01 g34158 ( .a(n_4317), .b(n_4624), .o(n_4350) );
NAND2_Z01 g34959 ( .a(n_3551), .b(GPR_15__0_), .o(n_3603) );
BUF_X2 newInst_999 ( .a(newNet_998), .o(newNet_999) );
BUF_X2 newInst_656 ( .a(newNet_655), .o(newNet_656) );
NAND2_Z01 g35405 ( .a(pZ_9_), .b(pZ_8_), .o(n_4514) );
XOR2_X1 g60854 ( .a(state_0_), .b(state_3_), .o(n_333) );
XOR2_X1 g34659 ( .a(n_3634), .b(pX_10_), .o(n_4564) );
NAND2_Z01 g59145 ( .a(n_1894), .b(n_120), .o(n_1954) );
NOR2_Z4 g57950 ( .a(n_2959), .b(n_1582), .o(n_3009) );
NAND2_Z01 g58723 ( .a(n_2207), .b(GPR_22__4_), .o(n_2384) );
NAND4_Z1 g58823 ( .a(n_1716), .b(n_1788), .c(n_2167), .d(n_1926), .o(n_2282) );
BUF_X2 newInst_179 ( .a(newNet_178), .o(newNet_179) );
INV_X1 g61114 ( .a(n_4487), .o(n_38) );
NAND2_Z01 g59091 ( .a(n_1871), .b(n_4606), .o(n_2016) );
BUF_X2 newInst_1345 ( .a(newNet_1344), .o(newNet_1345) );
AND3_X1 g59542 ( .a(n_1337), .b(n_1573), .c(n_306), .o(n_1586) );
BUF_X2 newInst_1389 ( .a(newNet_1388), .o(newNet_1389) );
fflopd pY_reg_10_ ( .CK(newNet_186), .D(n_2879), .Q(pY_10_) );
NAND2_Z01 g35068 ( .a(n_3496), .b(pmem_d_7), .o(n_3522) );
NAND2_Z01 g34432 ( .a(n_4098), .b(n_4635), .o(n_4105) );
NAND2_Z01 g60032 ( .a(n_768), .b(n_364), .o(n_1097) );
BUF_X2 newInst_1540 ( .a(newNet_1539), .o(newNet_1540) );
INV_Y1 g35320 ( .a(n_3352), .o(n_4559) );
XOR2_X1 g60167 ( .a(n_617), .b(n_87), .o(n_970) );
INV_X2 newInst_1409 ( .a(newNet_1408), .o(newNet_1409) );
fflopd pY_reg_3_ ( .CK(newNet_151), .D(n_2956), .Q(pY_3_) );
NAND2_Z01 g58666 ( .a(n_2213), .b(GPR_17__6_), .o(n_2440) );
NAND2_Z01 g59439 ( .a(n_852), .b(n_1650), .o(n_1681) );
INV_X2 newInst_939 ( .a(newNet_938), .o(newNet_939) );
BUF_X2 newInst_493 ( .a(newNet_300), .o(newNet_493) );
NAND2_Z01 g58239 ( .a(n_2754), .b(n_2194), .o(n_2828) );
BUF_X2 newInst_749 ( .a(newNet_435), .o(newNet_749) );
XOR2_X1 g35377 ( .a(pY_1_), .b(pY_0_), .o(n_3345) );
NAND2_Z01 g57983 ( .a(n_2942), .b(n_2215), .o(n_2989) );
NAND2_Z01 g59757 ( .a(n_1312), .b(io_do_6), .o(n_1367) );
INV_X2 newInst_704 ( .a(newNet_74), .o(newNet_704) );
AND2_X1 g35457 ( .a(pZ_4_), .b(pmem_d_11), .o(n_3267) );
BUF_X2 newInst_272 ( .a(newNet_271), .o(newNet_272) );
NAND3_Z1 g35248 ( .a(n_3252), .b(n_4560), .c(state_1_), .o(n_3426) );
NAND2_Z01 g59009 ( .a(n_1994), .b(n_1768), .o(n_2099) );
NOR2_Z1 g60625 ( .a(n_462), .b(n_197), .o(n_585) );
NAND2_Z01 g59440 ( .a(n_960), .b(n_1661), .o(n_1680) );
NOR2_Z1 g59934 ( .a(n_1121), .b(n_26), .o(n_1209) );
NOR2_Z1 g60033 ( .a(n_967), .b(n_966), .o(n_1116) );
BUF_X2 newInst_1318 ( .a(newNet_1295), .o(newNet_1318) );
BUF_X2 newInst_201 ( .a(newNet_150), .o(newNet_201) );
NAND2_Z01 g34946 ( .a(n_3552), .b(GPR_9__6_), .o(n_3616) );
XOR2_X1 g59672 ( .a(n_1382), .b(PC_9_), .o(n_1456) );
BUF_X2 newInst_1551 ( .a(newNet_1550), .o(newNet_1551) );
NOR4_Z1 g34234 ( .a(n_4191), .b(n_4192), .c(n_4240), .d(n_4107), .o(n_4297) );
XOR2_X1 g60386 ( .a(n_463), .b(io_do_3), .o(n_760) );
NAND4_Z1 g59541 ( .a(n_797), .b(n_1300), .c(n_1508), .d(n_1072), .o(n_1587) );
NOR2_Z1 g61005 ( .a(n_4654), .b(n_4655), .o(n_134) );
BUF_X2 newInst_1781 ( .a(newNet_1780), .o(newNet_1781) );
BUF_X2 newInst_400 ( .a(newNet_399), .o(newNet_400) );
XOR2_X1 g34464 ( .a(n_4059), .b(SP_2_), .o(n_4078) );
BUF_X2 newInst_1009 ( .a(newNet_1008), .o(newNet_1009) );
NOR2_Z1 g34304 ( .a(n_4612), .b(n_3766), .o(n_4229) );
NAND2_Z01 g58731 ( .a(n_2206), .b(GPR_23__4_), .o(n_2376) );
AND3_X1 g34495 ( .a(n_4006), .b(n_3977), .c(n_4018), .o(n_4049) );
NAND2_Z01 g34163 ( .a(n_4317), .b(pmem_d_1), .o(n_4345) );
BUF_X2 newInst_1041 ( .a(newNet_1040), .o(newNet_1041) );
AND2_X1 g60980 ( .a(n_4448), .b(n_4432), .o(n_188) );
NAND4_Z2 g35190 ( .a(n_3341), .b(n_3386), .c(n_3370), .d(n_3409), .o(n_4618) );
NAND2_Z01 g58294 ( .a(n_2702), .b(n_2248), .o(n_2776) );
NAND2_Z01 g34240 ( .a(io_do_5), .b(n_4177), .o(n_4293) );
NAND2_Z01 g34690 ( .a(n_3592), .b(GPR_23__7_), .o(n_3875) );
NAND2_Z01 g59179 ( .a(n_18), .b(n_606), .o(n_1928) );
NAND2_Z01 g60021 ( .a(n_968), .b(n_966), .o(n_1121) );
NAND2_Z01 g57835 ( .a(n_3041), .b(n_2390), .o(n_3075) );
NAND2_Z01 g58576 ( .a(n_2449), .b(n_1441), .o(n_2527) );
fflopd GPR_reg_12__5_ ( .CK(newNet_1629), .D(n_3019), .Q(GPR_12__5_) );
NAND2_Z01 g34624 ( .a(n_3646), .b(pX_11_), .o(n_3936) );
NAND2_Z02 g34451 ( .a(n_4068), .b(n_3930), .o(n_4610) );
NAND2_Z01 g60946 ( .a(n_44), .b(pmem_d_0), .o(n_248) );
NOR4_Z1 g34128 ( .a(n_4229), .b(n_4258), .c(n_4319), .d(n_4228), .o(n_4380) );
XOR2_X1 g35143 ( .a(n_3442), .b(pZ_4_), .o(n_3476) );
BUF_X2 newInst_500 ( .a(newNet_499), .o(newNet_500) );
NAND2_Z01 g59748 ( .a(n_1268), .b(SP_9_), .o(n_1374) );
BUF_X2 newInst_1354 ( .a(newNet_1353), .o(newNet_1354) );
NAND2_Z01 g58861 ( .a(n_2155), .b(GPR_14__7_), .o(n_2246) );
NOR2_Z3 g34202 ( .a(n_4556), .b(n_3259), .o(n_4325) );
NAND4_Z1 g34121 ( .a(n_4270), .b(n_4297), .c(n_4310), .d(n_4145), .o(dmem_a_1) );
BUF_X2 newInst_1620 ( .a(newNet_174), .o(newNet_1620) );
BUF_X2 newInst_557 ( .a(newNet_556), .o(newNet_557) );
XNOR2_X1 g35107 ( .a(n_4620), .b(pmem_d_3), .o(n_4466) );
NAND2_Z01 g34153 ( .a(n_4317), .b(n_4626), .o(n_4355) );
BUF_X2 newInst_990 ( .a(newNet_989), .o(newNet_990) );
BUF_X2 newInst_203 ( .a(newNet_202), .o(newNet_203) );
NOR2_Z1 g60959 ( .a(n_44), .b(pmem_d_1), .o(n_158) );
AND2_X1 g59373 ( .a(n_1678), .b(n_1140), .o(n_1764) );
BUF_X2 newInst_993 ( .a(newNet_696), .o(newNet_993) );
NOR2_Z1 g60795 ( .a(n_197), .b(n_258), .o(n_371) );
BUF_X2 newInst_921 ( .a(newNet_920), .o(newNet_921) );
BUF_X2 newInst_728 ( .a(newNet_727), .o(newNet_728) );
NAND2_Z01 g60787 ( .a(n_247), .b(n_35), .o(n_378) );
BUF_X2 newInst_1172 ( .a(newNet_1171), .o(newNet_1172) );
INV_X1 g60952 ( .a(n_188), .o(n_189) );
NAND2_Z01 g59054 ( .a(n_1902), .b(n_4587), .o(n_2053) );
fflopd pZ_reg_13_ ( .CK(newNet_98), .D(n_3095), .Q(pZ_13_) );
AND2_X1 g35288 ( .a(n_3239), .b(n_4640), .o(n_3387) );
NAND2_Z01 g34710 ( .a(n_3627), .b(GPR_15__6_), .o(n_3855) );
NAND2_Z01 g58762 ( .a(n_2203), .b(GPR_4__6_), .o(n_2338) );
NAND4_Z1 g59899 ( .a(n_490), .b(n_754), .c(n_996), .d(n_523), .o(n_1230) );
BUF_X2 newInst_155 ( .a(newNet_154), .o(newNet_155) );
BUF_X2 newInst_1334 ( .a(newNet_1333), .o(newNet_1334) );
NAND2_Z01 g60483 ( .a(Rd_1_), .b(n_340), .o(n_663) );
fflopd GPR_reg_15__3_ ( .CK(newNet_1504), .D(n_2860), .Q(GPR_15__3_) );
BUF_X2 newInst_1050 ( .a(newNet_522), .o(newNet_1050) );
fflopd GPR_reg_11__2_ ( .CK(newNet_1698), .D(n_2785), .Q(GPR_11__2_) );
NAND2_Z01 final_adder_mux_R16_278_6_g381 ( .a(final_adder_mux_R16_278_6_n_66), .b(final_adder_mux_R16_278_6_n_20), .o(final_adder_mux_R16_278_6_n_68) );
NAND2_Z01 g58153 ( .a(n_2812), .b(n_2243), .o(n_2860) );
NAND4_Z1 g60002 ( .a(n_895), .b(n_940), .c(n_914), .d(n_809), .o(n_1127) );
NAND4_Z1 g34595 ( .a(n_3700), .b(n_3845), .c(n_3754), .d(n_3701), .o(n_3965) );
AND2_X1 g58391 ( .a(n_2656), .b(n_2204), .o(n_2677) );
NOR2_Z1 g35335 ( .a(n_3222), .b(n_3288), .o(n_3335) );
BUF_X2 newInst_1090 ( .a(newNet_1089), .o(newNet_1090) );
NAND4_Z1 g59661 ( .a(n_1222), .b(n_1295), .c(n_66), .d(n_4636), .o(n_1485) );
XNOR2_X1 g58614 ( .a(n_2362), .b(n_1770), .o(n_2484) );
NOR3_Z1 g35095 ( .a(n_3249), .b(n_4656), .c(pmem_d_2), .o(n_4654) );
AND2_X1 g58386 ( .a(n_2657), .b(n_2206), .o(n_2682) );
NAND2_Z01 g59000 ( .a(n_2060), .b(n_1850), .o(n_2107) );
BUF_X2 newInst_1161 ( .a(newNet_1160), .o(newNet_1161) );
AND2_X1 g58265 ( .a(n_2752), .b(n_2205), .o(n_2802) );
NAND2_Z01 g57806 ( .a(n_3080), .b(n_2196), .o(n_3101) );
BUF_X2 newInst_859 ( .a(newNet_858), .o(newNet_859) );
NAND2_Z01 g35026 ( .a(n_3529), .b(n_3267), .o(n_3543) );
BUF_X2 newInst_756 ( .a(newNet_755), .o(newNet_756) );
NOR4_Z1 g58830 ( .a(n_4644), .b(n_69), .c(n_2082), .d(n_65), .o(n_2277) );
BUF_X2 newInst_890 ( .a(newNet_889), .o(newNet_890) );
BUF_X2 newInst_1557 ( .a(newNet_1556), .o(newNet_1557) );
BUF_X2 newInst_1000 ( .a(newNet_999), .o(newNet_1000) );
AND2_X1 g60358 ( .a(n_579), .b(n_261), .o(n_779) );
AND4_X1 g34208 ( .a(n_4642), .b(n_3540), .c(n_4480), .d(n_4664), .o(n_4318) );
INV_X1 g59212 ( .a(n_1891), .o(n_1890) );
NOR2_Z1 g60996 ( .a(n_4438), .b(n_4422), .o(n_140) );
NAND2_Z01 g35334 ( .a(n_3289), .b(pY_0_), .o(n_3336) );
NAND2_Z01 g60883 ( .a(n_4620), .b(pmem_d_3), .o(n_242) );
INV_X1 g58592 ( .a(n_2505), .o(n_2506) );
NAND2_Z01 final_adder_mux_R16_278_6_g428 ( .a(n_4443), .b(n_4427), .o(final_adder_mux_R16_278_6_n_20) );
INV_X2 drc_bufs61161 ( .a(n_24), .o(n_14) );
BUF_X2 newInst_1238 ( .a(newNet_1237), .o(newNet_1238) );
AND2_X1 g58398 ( .a(n_2656), .b(n_2201), .o(n_2670) );
BUF_X2 newInst_1406 ( .a(newNet_1405), .o(newNet_1406) );
NAND2_Z01 g34905 ( .a(n_3563), .b(pZ_4_), .o(n_3658) );
NAND2_Z01 g59869 ( .a(n_1201), .b(n_85), .o(n_1258) );
fflopd pZ_reg_0_ ( .CK(newNet_111), .D(n_2730), .Q(pZ_0_) );
BUF_X2 newInst_40 ( .a(newNet_39), .o(newNet_40) );
NAND4_Z1 g34578 ( .a(n_3680), .b(n_3800), .c(n_3801), .d(n_3799), .o(n_3982) );
NAND2_Z01 g58882 ( .a(n_2153), .b(GPR_8__6_), .o(n_2225) );
NAND2_Z01 g59415 ( .a(n_64), .b(n_1649), .o(n_1705) );
NAND2_Z01 g58168 ( .a(n_2798), .b(n_2325), .o(n_2842) );
NAND2_Z01 g60309 ( .a(n_570), .b(pZ_5_), .o(n_816) );
NAND2_Z01 g59557 ( .a(n_1517), .b(n_233), .o(n_1575) );
NOR4_Z1 g34079 ( .a(n_4196), .b(n_4244), .c(n_4383), .d(n_4190), .o(n_4394) );
AND2_X1 g60753 ( .a(n_118), .b(n_204), .o(n_389) );
BUF_X2 newInst_535 ( .a(newNet_344), .o(newNet_535) );
BUF_X2 newInst_342 ( .a(newNet_341), .o(newNet_342) );
INV_X1 drc_bufs61212 ( .a(n_340), .o(n_20) );
BUF_X2 newInst_783 ( .a(newNet_782), .o(newNet_783) );
BUF_X2 newInst_462 ( .a(newNet_461), .o(newNet_462) );
NOR2_Z1 g59350 ( .a(n_1700), .b(n_1647), .o(n_1763) );
NAND2_Z01 g59627 ( .a(n_1413), .b(io_sp_6_), .o(n_1500) );
BUF_X2 newInst_514 ( .a(newNet_513), .o(newNet_514) );
INV_X1 g61048 ( .a(state_2_), .o(n_104) );
NAND2_Z01 g59101 ( .a(n_1781), .b(n_1866), .o(n_2008) );
BUF_X2 newInst_189 ( .a(newNet_188), .o(newNet_189) );
fflopd GPR_reg_18__6_ ( .CK(newNet_1336), .D(n_3082), .Q(GPR_18__6_) );
BUF_X2 newInst_507 ( .a(newNet_506), .o(newNet_507) );
BUF_X2 newInst_182 ( .a(newNet_181), .o(newNet_182) );
BUF_X2 newInst_1672 ( .a(newNet_1671), .o(newNet_1672) );
BUF_X2 newInst_1082 ( .a(newNet_1081), .o(newNet_1082) );
INV_X1 g35322 ( .a(n_4660), .o(n_3348) );
NAND4_Z1 g57810 ( .a(n_1957), .b(n_2512), .c(n_3059), .d(n_1942), .o(n_3097) );
INV_X1 g34800 ( .a(n_4562), .o(n_3763) );
AND2_X1 g57748 ( .a(n_3115), .b(n_2203), .o(n_3123) );
NAND2_Z01 g60435 ( .a(n_20), .b(Rd_r_0_), .o(n_711) );
BUF_X2 newInst_633 ( .a(newNet_632), .o(newNet_633) );
BUF_X2 newInst_499 ( .a(newNet_498), .o(newNet_499) );
NAND2_Z01 g60698 ( .a(n_200), .b(GPR_12__1_), .o(n_440) );
NAND4_Z1 g60141 ( .a(n_546), .b(n_729), .c(n_665), .d(n_638), .o(n_991) );
BUF_X2 newInst_1495 ( .a(newNet_1494), .o(newNet_1495) );
AND2_X1 g34918 ( .a(n_3595), .b(pZ_10_), .o(n_3645) );
BUF_X2 newInst_942 ( .a(newNet_941), .o(newNet_942) );
fflopd SP_reg_10_ ( .CK(newNet_565), .D(n_1677), .Q(SP_10_) );
NAND2_Z01 g59611 ( .a(n_1452), .b(n_138), .o(n_1516) );
BUF_X2 newInst_1768 ( .a(newNet_1767), .o(newNet_1768) );
BUF_X2 newInst_1311 ( .a(newNet_1310), .o(newNet_1311) );
NAND2_Z01 g57710 ( .a(n_3130), .b(n_2405), .o(n_3159) );
INV_X1 g35471 ( .a(pX_8_), .o(n_3253) );
NAND2_Z01 g59084 ( .a(n_1903), .b(n_192), .o(n_2023) );
INV_X1 g35494 ( .a(pmem_d_7), .o(n_3232) );
AND2_X1 g59515 ( .a(n_1269), .b(n_1568), .o(n_1609) );
NAND2_Z01 g59573 ( .a(n_1483), .b(n_849), .o(n_1555) );
INV_X1 g35517 ( .a(PC_4_), .o(n_3211) );
NAND2_Z01 g58585 ( .a(n_2463), .b(pZ_6_), .o(n_2513) );
BUF_X2 newInst_32 ( .a(newNet_31), .o(newNet_32) );
NAND2_Z01 g34754 ( .a(n_3579), .b(GPR_12__4_), .o(n_3811) );
NAND2_Z01 g58444 ( .a(n_2641), .b(n_1732), .o(n_2649) );
XNOR2_X1 g35146 ( .a(n_3452), .b(PC_4_), .o(n_4547) );
NAND4_Z1 g59804 ( .a(n_715), .b(n_657), .c(n_1178), .d(n_545), .o(n_1324) );
BUF_X2 newInst_1303 ( .a(newNet_1302), .o(newNet_1303) );
AND2_X1 g59031 ( .a(n_1976), .b(n_1449), .o(n_2073) );
NAND2_Z01 g59821 ( .a(n_1171), .b(dmem_di_0), .o(n_1303) );
NAND2_Z01 g60919 ( .a(n_124), .b(pY_5_), .o(n_223) );
BUF_X2 newInst_826 ( .a(newNet_825), .o(newNet_826) );
NAND2_Z01 g60461 ( .a(n_342), .b(GPR_17__0_), .o(n_685) );
fflopd pX_reg_5_ ( .CK(newNet_214), .D(n_3098), .Q(pX_5_) );
NAND2_Z01 g58873 ( .a(n_2155), .b(GPR_14__2_), .o(n_2234) );
fflopd GPR_reg_19__3_ ( .CK(newNet_1299), .D(n_2856), .Q(GPR_19__3_) );
NAND2_Z01 g35408 ( .a(pZ_3_), .b(pmem_d_10), .o(n_3295) );
NAND4_Z1 g34569 ( .a(n_3841), .b(n_3842), .c(n_3844), .d(n_3840), .o(n_3991) );
NAND2_Z01 g34998 ( .a(n_3536), .b(n_3461), .o(n_3583) );
fflopd GPR_reg_20__4_ ( .CK(newNet_1197), .D(n_2934), .Q(GPR_20__4_) );
NAND4_Z1 g59988 ( .a(n_811), .b(n_941), .c(n_818), .d(n_906), .o(n_1141) );
BUF_X2 newInst_1078 ( .a(newNet_1077), .o(newNet_1078) );
AND2_X1 g35357 ( .a(n_3276), .b(pY_2_), .o(n_3349) );
AND2_X1 g35291 ( .a(n_3229), .b(n_3298), .o(n_3384) );
NOR2_Z1 g59295 ( .a(n_1036), .b(n_1770), .o(n_1816) );
NAND2_Z01 g60441 ( .a(n_358), .b(GPR_2__4_), .o(n_705) );
NAND2_Z01 g58495 ( .a(n_2572), .b(n_1836), .o(n_2602) );
BUF_X2 newInst_218 ( .a(newNet_217), .o(newNet_218) );
NAND2_Z01 g57772 ( .a(n_3099), .b(n_1433), .o(n_3109) );
NAND2_Z01 g58476 ( .a(n_2320), .b(n_2580), .o(n_2618) );
NAND2_Z01 g34865 ( .a(n_3592), .b(GPR_23__0_), .o(n_3698) );
NAND2_Z01 g59607 ( .a(n_1414), .b(io_di_0), .o(n_1519) );
AND2_X1 g57730 ( .a(n_3115), .b(n_2139), .o(n_3142) );
BUF_X2 newInst_744 ( .a(newNet_743), .o(newNet_744) );
BUF_X2 newInst_26 ( .a(newNet_25), .o(newNet_26) );
NAND2_Z01 g60704 ( .a(U_4_), .b(n_249), .o(n_434) );
NOR2_Z1 g34396 ( .a(n_4611), .b(n_3258), .o(n_4142) );
AND3_X1 g60665 ( .a(n_196), .b(n_4634), .c(n_4491), .o(n_481) );
AND2_X1 g57995 ( .a(n_2940), .b(n_2213), .o(n_2976) );
NAND2_Z01 g59640 ( .a(io_do_0), .b(n_1418), .o(n_1481) );
NOR4_Z1 g59731 ( .a(n_1105), .b(n_1131), .c(n_1132), .d(n_890), .o(n_1399) );
AND2_X1 g59981 ( .a(n_978), .b(n_977), .o(n_1159) );
NAND3_Z1 g58605 ( .a(n_2443), .b(n_1624), .c(n_4615), .o(n_2490) );
AND3_X1 g59037 ( .a(n_46), .b(n_1983), .c(pY_10_), .o(n_2071) );
NAND2_Z01 g60428 ( .a(n_361), .b(GPR_5__2_), .o(n_718) );
INV_Z1 g35485 ( .a(pY_0_), .o(n_4597) );
BUF_X2 newInst_441 ( .a(newNet_427), .o(newNet_441) );
BUF_X2 newInst_169 ( .a(newNet_168), .o(newNet_169) );
NAND2_Z01 g34336 ( .a(n_4165), .b(n_4539), .o(n_4198) );
BUF_X2 newInst_1162 ( .a(newNet_1161), .o(newNet_1162) );
INV_X1 g61078 ( .a(GPR_16__4_), .o(n_74) );
NAND2_Z01 g59859 ( .a(n_1156), .b(n_849), .o(n_1272) );
BUF_X2 newInst_549 ( .a(newNet_548), .o(newNet_549) );
INV_X1 g61100 ( .a(pmem_d_6), .o(n_52) );
BUF_X2 newInst_1527 ( .a(newNet_1526), .o(newNet_1527) );
fflopd Rd_r_reg_1_ ( .CK(newNet_589), .D(n_949), .Q(Rd_r_1_) );
NAND2_Z01 g58727 ( .a(n_2206), .b(GPR_23__0_), .o(n_2380) );
NAND2_Z01 g60898 ( .a(PC_6_), .b(PC_7_), .o(n_234) );
NAND2_Z01 g59337 ( .a(io_do_3), .b(n_30), .o(n_1803) );
NAND2_Z01 g57939 ( .a(n_2968), .b(n_2367), .o(n_3003) );
fflopd GPR_reg_15__7_ ( .CK(newNet_1486), .D(n_3164), .Q(GPR_15__7_) );
fflopd GPR_reg_0__2_ ( .CK(newNet_1801), .D(n_2734), .Q(GPR_0__2_) );
BUF_X2 newInst_1369 ( .a(newNet_1368), .o(newNet_1369) );
NAND2_Z01 g60517 ( .a(n_380), .b(GPR_6__1_), .o(n_629) );
NAND3_Z1 g58984 ( .a(n_1939), .b(n_1747), .c(n_789), .o(n_2123) );
NOR2_Z1 g59135 ( .a(n_1873), .b(n_865), .o(n_1963) );
NAND2_Z01 g57948 ( .a(n_905), .b(n_2985), .o(n_3011) );
NAND2_Z01 g60908 ( .a(PC_7_), .b(pmem_d_7), .o(n_264) );
AND2_X1 g58817 ( .a(n_2216), .b(n_2058), .o(n_2361) );
NAND2_Z01 g34095 ( .a(n_4373), .b(n_4372), .o(n_4437) );
NAND2_Z01 g60551 ( .a(n_360), .b(GPR_1__3_), .o(n_555) );
BUF_X2 newInst_627 ( .a(newNet_626), .o(newNet_627) );
NAND2_Z01 g58441 ( .a(n_2621), .b(n_13), .o(n_2652) );
NAND2_Z01 g59057 ( .a(n_1902), .b(n_4585), .o(n_2050) );
NAND2_Z01 g60573 ( .a(n_372), .b(pX_9_), .o(n_538) );
NAND2_Z01 g59330 ( .a(n_1690), .b(n_1724), .o(n_1783) );
BUF_X2 newInst_1829 ( .a(newNet_1828), .o(newNet_1829) );
BUF_X2 newInst_1548 ( .a(newNet_1547), .o(newNet_1548) );
NAND3_Z1 g34084 ( .a(n_4378), .b(n_4323), .c(n_4231), .o(dmem_do_6) );
INV_X1 g34473 ( .a(n_4068), .o(n_4069) );
NAND2_Z01 g59604 ( .a(n_1411), .b(n_4618), .o(n_1522) );
INV_X1 g35040 ( .a(n_4590), .o(n_3532) );
BUF_X2 newInst_1384 ( .a(newNet_1383), .o(newNet_1384) );
BUF_X2 newInst_918 ( .a(newNet_917), .o(newNet_918) );
INV_X1 g34630 ( .a(n_4645), .o(n_3930) );
BUF_X2 newInst_409 ( .a(newNet_408), .o(newNet_409) );
BUF_X2 newInst_364 ( .a(newNet_142), .o(newNet_364) );
NAND2_Z01 g58768 ( .a(n_2202), .b(GPR_5__4_), .o(n_2332) );
INV_X1 g60013 ( .a(n_1114), .o(n_1113) );
BUF_X2 newInst_669 ( .a(newNet_668), .o(newNet_669) );
NOR3_Z1 g59726 ( .a(n_1025), .b(n_1266), .c(n_1285), .o(n_1401) );
INV_X1 drc_bufs61222 ( .a(n_1489), .o(n_9) );
NAND2_Z01 g60516 ( .a(n_347), .b(GPR_9__0_), .o(n_630) );
XOR2_X1 g34931 ( .a(n_3554), .b(PC_9_), .o(n_4538) );
NOR4_Z1 g34229 ( .a(n_4208), .b(n_4209), .c(n_4265), .d(n_4114), .o(n_4302) );
INV_X1 g58746 ( .a(n_2357), .o(n_2358) );
NAND2_Z01 g59108 ( .a(n_1871), .b(pZ_14_), .o(n_2001) );
INV_X1 g60094 ( .a(n_995), .o(n_1030) );
BUF_X2 newInst_1593 ( .a(newNet_1592), .o(newNet_1593) );
NAND2_Z01 g60066 ( .a(n_852), .b(io_do_1), .o(n_1068) );
NAND2_Z01 g57884 ( .a(n_3011), .b(n_13), .o(n_3054) );
NAND2_Z01 g58897 ( .a(n_2158), .b(GPR_12__7_), .o(n_2185) );
NAND2_Z01 g60465 ( .a(n_372), .b(U_11_), .o(n_681) );
NAND2_Z01 g34441 ( .a(n_4077), .b(SP_3_), .o(n_4099) );
NOR3_Z1 g60136 ( .a(n_517), .b(n_761), .c(n_518), .o(n_996) );
NAND2_Z01 g57695 ( .a(n_3144), .b(n_1581), .o(n_3171) );
NAND2_Z01 g59784 ( .a(n_1268), .b(n_593), .o(n_1340) );
NAND2_Z01 g34787 ( .a(n_3636), .b(GPR_10__3_), .o(n_3778) );
NAND2_Z01 g34637 ( .a(n_3769), .b(pZ_4_), .o(n_3923) );
AND2_X1 g59361 ( .a(n_1671), .b(pmem_d_9), .o(n_1752) );
BUF_X2 newInst_770 ( .a(newNet_769), .o(newNet_770) );
NAND2_Z01 g58468 ( .a(n_2396), .b(n_2589), .o(n_2628) );
BUF_X2 newInst_1390 ( .a(newNet_50), .o(newNet_1390) );
BUF_X2 newInst_341 ( .a(newNet_340), .o(newNet_341) );
NAND2_Z01 g60977 ( .a(n_83), .b(n_52), .o(n_148) );
BUF_X2 newInst_291 ( .a(newNet_290), .o(newNet_291) );
NAND2_Z01 g60277 ( .a(n_574), .b(GPR_10__3_), .o(n_869) );
NAND2_Z01 g60912 ( .a(PC_5_), .b(pmem_d_8), .o(n_229) );
NAND2_Z01 g57807 ( .a(n_3079), .b(n_2198), .o(n_3100) );
INV_X1 g34798 ( .a(n_3765), .o(n_4588) );
NAND2_Z01 g35059 ( .a(n_3502), .b(n_3443), .o(n_3525) );
NAND2_Z01 g59102 ( .a(n_1223), .b(n_1878), .o(n_2007) );
XOR2_X1 g35197 ( .a(n_3356), .b(pX_3_), .o(n_4571) );
NAND2_Z01 g34855 ( .a(n_3587), .b(GPR_2__0_), .o(n_3708) );
BUF_X2 newInst_660 ( .a(newNet_659), .o(newNet_660) );
NAND2_Z01 g34881 ( .a(n_3630), .b(pX_5_), .o(n_3682) );
BUF_X2 newInst_1470 ( .a(newNet_1469), .o(newNet_1470) );
BUF_X2 newInst_171 ( .a(newNet_170), .o(newNet_171) );
INV_X1 g35478 ( .a(SP_10_), .o(n_3246) );
NOR2_Z1 g35431 ( .a(n_3217), .b(pmem_d_12), .o(n_3274) );
NAND2_Z01 g59026 ( .a(n_2059), .b(n_47), .o(n_2090) );
AND2_X1 g58366 ( .a(n_2657), .b(n_2155), .o(n_2705) );
BUF_X2 newInst_1716 ( .a(newNet_1715), .o(newNet_1716) );
NAND2_Z01 g59154 ( .a(n_1896), .b(n_94), .o(n_1945) );
AND2_X1 g59763 ( .a(n_1269), .b(n_1309), .o(n_1362) );
NAND4_Z1 g57763 ( .a(n_1915), .b(n_2513), .c(n_3106), .d(n_2030), .o(n_3112) );
BUF_X2 newInst_213 ( .a(newNet_212), .o(newNet_213) );
NAND2_Z01 g60734 ( .a(SP_10_), .b(n_180), .o(n_405) );
NAND2_Z01 g34752 ( .a(n_3587), .b(GPR_2__4_), .o(n_3813) );
NAND2_Z01 g58777 ( .a(n_2201), .b(GPR_6__5_), .o(n_2323) );
NAND2_Z01 g59844 ( .a(n_1181), .b(n_224), .o(n_1282) );
NOR2_Z1 g34902 ( .a(n_3562), .b(n_3230), .o(n_3661) );
BUF_X2 newInst_1629 ( .a(newNet_1628), .o(newNet_1629) );
NAND2_Z01 g34324 ( .a(n_4157), .b(n_4558), .o(n_4480) );
NAND2_Z01 g34822 ( .a(n_3628), .b(GPR_19__2_), .o(n_3741) );
NOR2_Z1 g34414 ( .a(n_4610), .b(n_3561), .o(n_4123) );
BUF_X2 newInst_581 ( .a(newNet_580), .o(newNet_581) );
NOR2_Z2 g60962 ( .a(n_71), .b(pmem_d_9), .o(n_200) );
AND2_X1 g60656 ( .a(n_339), .b(pmem_d_0), .o(n_487) );
AND2_X1 g57753 ( .a(n_3115), .b(n_2140), .o(n_3118) );
fflopd GPR_Rd_r_reg_6_ ( .CK(newNet_1837), .D(io_do_6), .Q(GPR_Rd_r_6_) );
NAND2_Z01 g58447 ( .a(n_2622), .b(n_2194), .o(n_2646) );
NAND2_Z01 g60413 ( .a(n_380), .b(GPR_4__5_), .o(n_733) );
AND2_X1 final_adder_mux_R16_278_6_g441 ( .a(n_4440), .b(n_4424), .o(final_adder_mux_R16_278_6_n_8) );
NAND4_Z1 g34382 ( .a(n_4630), .b(n_3522), .c(n_4064), .d(n_4558), .o(n_4157) );
AND2_X1 g60746 ( .a(n_88), .b(n_250), .o(n_396) );
NOR2_Z1 g60840 ( .a(n_202), .b(n_250), .o(n_341) );
NAND2_Z01 g59125 ( .a(n_1894), .b(n_1286), .o(n_1986) );
BUF_X2 newInst_643 ( .a(newNet_642), .o(newNet_643) );
NAND2_Z01 g35447 ( .a(n_3236), .b(n_3249), .o(n_4489) );
fflopd GPR_reg_16__0_ ( .CK(newNet_1479), .D(n_2633), .Q(GPR_16__0_) );
NAND2_Z01 g58640 ( .a(n_2358), .b(pZ_2_), .o(n_2456) );
BUF_X2 newInst_1213 ( .a(newNet_1212), .o(newNet_1213) );
fflopd U_reg_8_ ( .CK(newNet_363), .D(n_2718), .Q(U_8_) );
AND2_X1 g57903 ( .a(n_3009), .b(n_2202), .o(n_3035) );
BUF_X2 newInst_452 ( .a(newNet_451), .o(newNet_452) );
BUF_X2 newInst_145 ( .a(newNet_144), .o(newNet_145) );
BUF_X2 newInst_1132 ( .a(newNet_125), .o(newNet_1132) );
fflopd GPR_reg_4__4_ ( .CK(newNet_905), .D(n_2928), .Q(GPR_4__4_) );
AND3_X1 g59657 ( .a(n_80), .b(n_1390), .c(pX_10_), .o(n_1469) );
NAND2_Z01 g34909 ( .a(n_3633), .b(pZ_9_), .o(n_3654) );
BUF_X2 newInst_1498 ( .a(newNet_1497), .o(newNet_1498) );
NAND2_Z01 g59742 ( .a(n_1267), .b(Z), .o(n_1380) );
BUF_X2 newInst_1796 ( .a(newNet_1795), .o(newNet_1796) );
BUF_X2 newInst_1397 ( .a(newNet_1396), .o(newNet_1397) );
NAND2_Z01 g60720 ( .a(SP_15_), .b(n_180), .o(n_418) );
INV_X1 g35424 ( .a(n_3280), .o(n_3279) );
NOR2_Z1 g35440 ( .a(pmem_d_15), .b(pmem_d_14), .o(n_4486) );
NAND2_Z01 g59852 ( .a(n_1161), .b(n_97), .o(n_1309) );
BUF_X2 newInst_1541 ( .a(newNet_1540), .o(newNet_1541) );
fflopd pZ_reg_10_ ( .CK(newNet_110), .D(n_2875), .Q(pZ_10_) );
NOR2_Z1 g34318 ( .a(n_16064_BAR), .b(n_3500), .o(n_4215) );
AND2_X1 g57891 ( .a(n_3009), .b(n_2214), .o(n_3047) );
NAND2_Z01 g34819 ( .a(n_3591), .b(U_10_), .o(n_3744) );
BUF_X2 newInst_888 ( .a(newNet_887), .o(newNet_888) );
fflopd pY_reg_11_ ( .CK(newNet_176), .D(n_2957), .Q(pY_11_) );
INV_X1 g34557 ( .a(n_4649), .o(n_4002) );
NAND2_Z01 g58836 ( .a(n_2159), .b(GPR_10__2_), .o(n_2271) );
NAND2_Z01 g59817 ( .a(n_1190), .b(n_220), .o(n_1315) );
BUF_X2 newInst_732 ( .a(newNet_731), .o(newNet_732) );
XOR2_X1 g58658 ( .a(n_2219), .b(n_1831), .o(n_2444) );
NAND2_Z01 g35456 ( .a(n_3251), .b(n_3225), .o(n_4584) );
BUF_X2 newInst_853 ( .a(newNet_852), .o(newNet_853) );
NAND2_Z01 g57720 ( .a(n_3120), .b(n_2312), .o(n_3147) );
BUF_X2 newInst_1233 ( .a(newNet_1232), .o(newNet_1233) );
fflopd GPR_reg_14__4_ ( .CK(newNet_1549), .D(n_2945), .Q(GPR_14__4_) );
NAND2_Z01 g34939 ( .a(n_3552), .b(GPR_9__7_), .o(n_3623) );
BUF_X2 newInst_833 ( .a(newNet_832), .o(newNet_833) );
NAND2_Z01 g59643 ( .a(n_1418), .b(io_do_5), .o(n_1478) );
BUF_X2 newInst_1226 ( .a(newNet_1225), .o(newNet_1226) );
NOR2_Z1 g35138 ( .a(n_4651), .b(n_4479), .o(n_3473) );
XOR2_X1 g59673 ( .a(n_1349), .b(n_112), .o(n_1455) );
BUF_X2 newInst_1426 ( .a(newNet_1425), .o(newNet_1426) );
fflopd SP_reg_14_ ( .CK(newNet_538), .D(n_1906), .Q(SP_14_) );
BUF_X2 newInst_1438 ( .a(newNet_1437), .o(newNet_1438) );
BUF_X2 newInst_1152 ( .a(newNet_1151), .o(newNet_1152) );
NAND2_Z01 g60193 ( .a(n_709), .b(n_639), .o(n_952) );
XOR2_X1 final_adder_mux_R16_278_6_g409 ( .a(n_4446), .b(n_4430), .o(final_adder_mux_R16_278_6_n_40) );
fflopd V_reg ( .CK(newNet_353), .D(n_3109), .Q(V) );
NAND2_Z01 g34723 ( .a(n_3584), .b(GPR_20__5_), .o(n_3842) );
INV_X2 g34198 ( .a(n_4325), .o(n_4324) );
BUF_X2 newInst_247 ( .a(newNet_246), .o(newNet_247) );
NAND2_Z01 g59061 ( .a(n_1902), .b(n_4593), .o(n_2046) );
NOR2_Z1 g58650 ( .a(n_2275), .b(n_579), .o(n_2451) );
fflopd pY_reg_7_ ( .CK(newNet_133), .D(n_3187), .Q(pY_7_) );
NAND4_Z1 g59496 ( .a(n_1341), .b(n_1476), .c(n_1567), .d(n_499), .o(n_1632) );
NAND2_Z01 g58770 ( .a(n_2202), .b(GPR_5__6_), .o(n_2330) );
NOR2_Z1 g35207 ( .a(n_3369), .b(n_3373), .o(n_3441) );
NOR2_Z1 g34376 ( .a(n_4125), .b(n_4069), .o(n_4165) );
BUF_X2 newInst_11 ( .a(newNet_10), .o(newNet_11) );
NAND2_Z01 g58714 ( .a(n_2208), .b(GPR_21__3_), .o(n_2393) );
NOR2_Z1 g34366 ( .a(n_4129), .b(n_3469), .o(n_4169) );
BUF_X2 newInst_1037 ( .a(newNet_1036), .o(newNet_1037) );
NAND2_Z01 g34641 ( .a(n_3769), .b(pZ_8_), .o(n_3919) );
AND3_X1 g35249 ( .a(n_3227), .b(n_4560), .c(state_2_), .o(n_3416) );
NOR2_Z1 g59164 ( .a(n_1890), .b(n_1686), .o(n_1980) );
INV_X2 newInst_751 ( .a(newNet_750), .o(newNet_751) );
NAND2_Z03 g34222 ( .a(n_4292), .b(n_3996), .o(io_do_6) );
BUF_X2 newInst_1604 ( .a(newNet_1603), .o(newNet_1604) );
NAND3_Z1 g59893 ( .a(io_do_1), .b(n_1026), .c(n_378), .o(n_1236) );
NAND2_Z01 g58309 ( .a(n_2684), .b(n_2387), .o(n_2761) );
NAND2_Z01 g59618 ( .a(n_1413), .b(io_sp_3_), .o(n_1509) );
NAND2_Z01 g34101 ( .a(n_4361), .b(n_4360), .o(n_4443) );
NAND2_Z01 g34876 ( .a(n_3568), .b(GPR_22__7_), .o(n_3687) );
NOR2_Z1 g59012 ( .a(n_1981), .b(n_122), .o(n_2096) );
NOR2_Z1 g35302 ( .a(n_3226), .b(n_3309), .o(n_3373) );
BUF_X2 newInst_1653 ( .a(newNet_1652), .o(newNet_1653) );
BUF_X2 newInst_972 ( .a(newNet_971), .o(newNet_972) );
NAND4_Z1 g58488 ( .a(n_1302), .b(n_1513), .c(n_2566), .d(n_1056), .o(n_2608) );
BUF_X2 newInst_1614 ( .a(newNet_976), .o(newNet_1614) );
BUF_X2 newInst_1110 ( .a(newNet_1109), .o(newNet_1110) );
AND2_X1 g58377 ( .a(n_2657), .b(n_2210), .o(n_2694) );
XOR2_X1 g59257 ( .a(n_1807), .b(n_316), .o(n_1855) );
NAND2_Z01 final_adder_mux_R16_278_6_g434 ( .a(n_4438), .b(n_4422), .o(final_adder_mux_R16_278_6_n_15) );
XOR2_X1 final_adder_mux_R16_278_6_g400 ( .a(final_adder_mux_R16_278_6_n_46), .b(final_adder_mux_R16_278_6_n_37), .o(R16_2_) );
NAND2_Z01 g60718 ( .a(U_12_), .b(n_249), .o(n_420) );
NAND2_Z01 g60724 ( .a(n_200), .b(GPR_12__5_), .o(n_414) );
NAND4_Z1 g34575 ( .a(n_3812), .b(n_3813), .c(n_3811), .d(n_3810), .o(n_3985) );
NOR2_Z1 g58926 ( .a(n_2117), .b(n_1619), .o(n_2177) );
NAND2_Z01 g59328 ( .a(n_1700), .b(n_4538), .o(n_1785) );
NOR2_Z1 g35307 ( .a(n_3219), .b(n_3288), .o(n_3369) );
NAND4_Z2 g35180 ( .a(n_3395), .b(n_3391), .c(n_3390), .d(n_3394), .o(n_4615) );
NAND2_Z01 g58976 ( .a(n_2084), .b(n_1211), .o(n_2131) );
NAND2_Z01 g60450 ( .a(n_374), .b(GPR_14__1_), .o(n_696) );
fflopd GPR_reg_16__2_ ( .CK(newNet_1471), .D(n_2773), .Q(GPR_16__2_) );
AND2_X1 g60624 ( .a(n_329), .b(n_4451), .o(n_505) );
AND2_X1 g60595 ( .a(n_362), .b(PC_3_), .o(n_602) );
NAND2_Z01 g34772 ( .a(n_3585), .b(GPR_13__4_), .o(n_3793) );
NAND2_Z01 g34717 ( .a(n_3591), .b(U_14_), .o(n_3848) );
AND2_X1 g59977 ( .a(n_563), .b(n_1031), .o(n_1148) );
NAND2_Z01 g58730 ( .a(n_2206), .b(GPR_23__3_), .o(n_2377) );
NAND2_Z01 g59272 ( .a(io_do_2), .b(n_1765), .o(n_1852) );
BUF_X2 newInst_695 ( .a(newNet_694), .o(newNet_695) );
NOR2_Z1 g34346 ( .a(n_4157), .b(n_4559), .o(n_4188) );
NAND2_Z01 g58458 ( .a(n_2600), .b(n_2265), .o(n_2638) );
NAND2_Z01 g59521 ( .a(n_1550), .b(n_335), .o(n_1620) );
NOR2_Z1 g34607 ( .a(n_3715), .b(n_3714), .o(n_3953) );
INV_X1 drc_bufs61234 ( .a(n_1764), .o(n_5) );
AND2_X1 g57736 ( .a(n_3115), .b(n_2156), .o(n_3136) );
NOR2_Z1 g58540 ( .a(n_2537), .b(n_24), .o(n_2558) );
AND2_X1 g35012 ( .a(n_3511), .b(n_3548), .o(n_3565) );
BUF_X2 newInst_831 ( .a(newNet_830), .o(newNet_831) );
NAND2_Z01 g60582 ( .a(io_do_5), .b(n_343), .o(n_530) );
INV_X1 drc_bufs61238 ( .a(n_345), .o(n_21) );
AND2_X1 g59965 ( .a(n_1025), .b(n_1031), .o(n_1154) );
BUF_X2 newInst_90 ( .a(newNet_89), .o(newNet_90) );
NAND2_Z02 g58915 ( .a(n_2160), .b(n_1203), .o(n_2207) );
NAND2_Z01 g57704 ( .a(n_3138), .b(n_2246), .o(n_3165) );
BUF_X2 newInst_687 ( .a(newNet_686), .o(newNet_687) );
NAND2_Z01 g34891 ( .a(n_3630), .b(pX_9_), .o(n_3672) );
BUF_X2 newInst_357 ( .a(newNet_356), .o(newNet_357) );
NOR2_Z1 g34274 ( .a(n_4175), .b(n_4574), .o(n_4259) );
XOR2_X1 g35072 ( .a(n_3480), .b(pY_6_), .o(n_3521) );
NAND2_Z01 g35034 ( .a(n_4520), .b(n_3240), .o(n_3546) );
NAND2_Z01 g34627 ( .a(n_3769), .b(pZ_1_), .o(n_3933) );
AND2_X1 g59794 ( .a(n_1266), .b(n_1031), .o(n_1330) );
NAND2_Z01 g59888 ( .a(n_1169), .b(n_1166), .o(n_1239) );
NAND2_Z01 final_adder_mux_R16_278_6_g399 ( .a(final_adder_mux_R16_278_6_n_48), .b(final_adder_mux_R16_278_6_n_22), .o(final_adder_mux_R16_278_6_n_50) );
NOR2_Z1 g34871 ( .a(n_3580), .b(n_4407), .o(n_3692) );
NAND2_Z01 g58323 ( .a(n_2671), .b(n_2327), .o(n_2742) );
NAND2_Z01 g58407 ( .a(n_2655), .b(n_1702), .o(n_2661) );
AND2_X1 g59848 ( .a(n_1219), .b(n_462), .o(n_1278) );
INV_X1 g35229 ( .a(n_4651), .o(n_3429) );
NAND2_Z01 g59321 ( .a(n_1700), .b(n_4549), .o(n_1792) );
BUF_X2 newInst_229 ( .a(newNet_228), .o(newNet_229) );
BUF_X2 newInst_192 ( .a(newNet_191), .o(newNet_192) );
NAND2_Z01 g60269 ( .a(n_584), .b(GPR_18__5_), .o(n_877) );
NOR2_Z1 g59471 ( .a(n_1619), .b(n_71), .o(n_1653) );
BUF_X2 newInst_352 ( .a(newNet_351), .o(newNet_352) );
fflopd PC_reg_8_ ( .CK(newNet_608), .D(n_2279), .Q(PC_8_) );
BUF_X2 newInst_1104 ( .a(newNet_1103), .o(newNet_1104) );
AND2_X1 g57739 ( .a(n_3115), .b(n_2212), .o(n_3133) );
NAND2_Z01 g58996 ( .a(n_2061), .b(n_963), .o(n_2116) );
NAND2_Z01 g34531 ( .a(n_3657), .b(n_3939), .o(n_4014) );
BUF_X2 newInst_1292 ( .a(newNet_1291), .o(newNet_1292) );
NAND2_Z01 g35210 ( .a(n_3326), .b(n_3291), .o(n_3450) );
XOR2_X1 g34500 ( .a(n_4027), .b(pZ_7_), .o(n_4044) );
AND2_X1 g58376 ( .a(n_2657), .b(n_2211), .o(n_2695) );
INV_X1 g61045 ( .a(pZ_2_), .o(n_107) );
AND2_X1 g60838 ( .a(n_258), .b(pmem_d_1), .o(n_344) );
BUF_X2 newInst_251 ( .a(newNet_222), .o(newNet_251) );
INV_X1 g58043 ( .a(n_2940), .o(n_2939) );
BUF_X2 newInst_194 ( .a(newNet_191), .o(newNet_194) );
NAND2_Z01 g58630 ( .a(n_2356), .b(n_2010), .o(n_2480) );
NAND2_X2 g58907 ( .a(n_2144), .b(n_2090), .o(n_2215) );
BUF_X2 newInst_1762 ( .a(newNet_1761), .o(newNet_1762) );
NOR2_Z1 g60968 ( .a(n_35), .b(pmem_d_2), .o(n_152) );
BUF_X2 newInst_1853 ( .a(newNet_1852), .o(newNet_1853) );
INV_X1 drc_bufs61233 ( .a(n_5), .o(n_6) );
NAND2_Z01 g57848 ( .a(n_3030), .b(n_2288), .o(n_3064) );
NOR2_Z1 g35005 ( .a(n_3550), .b(n_3490), .o(n_3572) );
NAND3_Z1 g58176 ( .a(n_104), .b(n_2788), .c(n_41), .o(n_2836) );
XNOR2_X1 g34437 ( .a(n_4073), .b(pZ_11_), .o(n_4102) );
AND4_X1 g58529 ( .a(n_1606), .b(n_1605), .c(n_2553), .d(n_1743), .o(n_2568) );
NAND2_Z01 g58556 ( .a(n_2526), .b(n_1933), .o(n_2541) );
INV_X1 g59282 ( .a(n_1830), .o(n_1831) );
NOR2_Z1 g60613 ( .a(n_337), .b(n_160), .o(n_511) );
AND2_X1 g57896 ( .a(n_3009), .b(n_2209), .o(n_3042) );
NAND2_Z01 g34829 ( .a(n_3573), .b(U_1_), .o(n_3734) );
NAND4_Z1 g58135 ( .a(n_1944), .b(n_2476), .c(n_2825), .d(n_2049), .o(n_2878) );
NAND3_Z1 g60086 ( .a(n_544), .b(n_723), .c(n_628), .o(n_1051) );
BUF_X2 newInst_1589 ( .a(newNet_1588), .o(newNet_1589) );
INV_X1 g61074 ( .a(pX_12_), .o(n_78) );
BUF_X2 newInst_1109 ( .a(newNet_303), .o(newNet_1109) );
NOR2_Z1 g34448 ( .a(n_4072), .b(n_3930), .o(n_4092) );
BUF_X2 newInst_790 ( .a(newNet_789), .o(newNet_790) );
NOR2_Z1 g35167 ( .a(n_3445), .b(pmem_d_9), .o(n_4479) );
AND2_X1 g58400 ( .a(n_2656), .b(n_2200), .o(n_2668) );
NAND2_Z01 g60037 ( .a(n_849), .b(pmem_d_14), .o(n_1093) );
NAND2_X2 g58904 ( .a(n_2137), .b(n_2113), .o(n_2218) );
NOR3_Z1 g59188 ( .a(n_1449), .b(n_1895), .c(n_89), .o(n_1919) );
NAND2_Z01 final_adder_mux_R16_278_6_g421 ( .a(n_4441), .b(n_4425), .o(final_adder_mux_R16_278_6_n_27) );
BUF_X2 newInst_1512 ( .a(newNet_637), .o(newNet_1512) );
AND2_X1 g58519 ( .a(n_2567), .b(n_2199), .o(n_2577) );
NOR4_Z1 g58973 ( .a(n_1257), .b(n_2008), .c(n_1457), .d(n_1263), .o(n_2133) );
AND2_X1 g57908 ( .a(n_3009), .b(n_14), .o(n_3056) );
fflopd pX_reg_15_ ( .CK(newNet_250), .D(n_3192), .Q(pX_15_) );
NOR2_Z1 g34423 ( .a(n_4610), .b(n_3476), .o(n_4114) );
NOR2_Z1 g35438 ( .a(pY_1_), .b(pmem_d_1), .o(n_3272) );
BUF_X2 newInst_1139 ( .a(newNet_1138), .o(newNet_1139) );
BUF_X2 newInst_928 ( .a(newNet_927), .o(newNet_928) );
NOR2_Z1 g35343 ( .a(n_4684), .b(n_3233), .o(n_3359) );
BUF_X2 newInst_1457 ( .a(newNet_1456), .o(newNet_1457) );
AND2_X1 g58121 ( .a(n_2850), .b(n_2204), .o(n_2891) );
NOR2_Z1 g59715 ( .a(n_1269), .b(n_1351), .o(n_1410) );
BUF_X2 newInst_1066 ( .a(newNet_1065), .o(newNet_1066) );
BUF_X2 newInst_475 ( .a(newNet_159), .o(newNet_475) );
NAND2_Z01 g34119 ( .a(io_do_0), .b(n_4177), .o(n_4384) );
AND2_X1 g59412 ( .a(io_do_7), .b(n_1661), .o(n_1732) );
NOR2_Z1 g59262 ( .a(n_1763), .b(n_4417), .o(n_1848) );
fflopd GPR_reg_21__4_ ( .CK(newNet_1131), .D(n_2933), .Q(GPR_21__4_) );
NAND2_Z01 g58790 ( .a(n_2213), .b(GPR_17__1_), .o(n_2310) );
NAND2_Z01 g35392 ( .a(PC_1_), .b(PC_0_), .o(n_3312) );
NAND2_Z01 g60251 ( .a(n_574), .b(GPR_10__7_), .o(n_894) );
BUF_X2 newInst_239 ( .a(newNet_238), .o(newNet_239) );
NAND2_Z01 g60228 ( .a(n_575), .b(GPR_2__0_), .o(n_917) );
NAND2_Z01 g35396 ( .a(pmem_d_15), .b(pmem_d_14), .o(n_3311) );
NOR2_Z1 g59174 ( .a(n_1036), .b(n_1876), .o(n_1932) );
BUF_X2 newInst_372 ( .a(newNet_169), .o(newNet_372) );
BUF_X2 newInst_275 ( .a(newNet_274), .o(newNet_275) );
INV_X1 g34982 ( .a(n_3565), .o(n_3564) );
NAND2_Z01 g59071 ( .a(n_1871), .b(n_4598), .o(n_2036) );
NAND2_Z01 g60802 ( .a(n_201), .b(n_35), .o(n_365) );
BUF_X2 newInst_1858 ( .a(newNet_1857), .o(newNet_1858) );
NAND2_Z01 g34734 ( .a(n_3627), .b(GPR_15__5_), .o(n_3831) );
NAND2_Z01 g60639 ( .a(n_326), .b(n_179), .o(n_497) );
fflopd SP_reg_7_ ( .CK(newNet_479), .D(n_1741), .Q(SP_7_) );
NAND2_Z01 g60302 ( .a(n_618), .b(n_167), .o(n_822) );
NAND2_Z01 g59833 ( .a(n_1206), .b(io_do_2), .o(n_1292) );
NAND2_Z01 g60398 ( .a(n_472), .b(state_2_), .o(n_748) );
NOR2_Z1 g34293 ( .a(n_4163), .b(n_3231), .o(n_4240) );
NAND2_Z01 g35239 ( .a(n_3360), .b(n_3248), .o(n_3419) );
NAND4_Z1 g34086 ( .a(n_4277), .b(n_4299), .c(n_4329), .d(n_4141), .o(dmem_a_7) );
INV_X1 g60875 ( .a(n_250), .o(n_249) );
AND2_X1 g59588 ( .a(n_1462), .b(n_612), .o(n_1540) );
AND2_X1 g35247 ( .a(n_3349), .b(pY_3_), .o(n_3427) );
NAND2_Z01 g58102 ( .a(n_2852), .b(n_13), .o(n_2911) );
INV_X1 g35232 ( .a(n_4608), .o(n_3422) );
NAND2_Z01 g34668 ( .a(n_3602), .b(n_3611), .o(n_3897) );
BUF_X2 newInst_571 ( .a(newNet_570), .o(newNet_571) );
AND4_X1 g59304 ( .a(n_4621), .b(n_4619), .c(n_1634), .d(n_4623), .o(n_1810) );
NAND2_Z01 g34911 ( .a(n_3577), .b(pY_0_), .o(n_3652) );
NAND2_Z01 g59325 ( .a(n_1700), .b(n_4541), .o(n_1788) );
AND2_X1 g57746 ( .a(n_3115), .b(n_2205), .o(n_3125) );
NAND2_Z01 g58057 ( .a(n_2887), .b(n_2315), .o(n_2925) );
NAND2_Z01 g60075 ( .a(n_841), .b(io_do_2), .o(n_1060) );
NAND4_Z1 g59045 ( .a(n_1822), .b(n_1882), .c(n_1151), .d(n_1821), .o(n_2064) );
NOR3_Z1 g59301 ( .a(n_1704), .b(n_1147), .c(n_1311), .o(n_1826) );
NAND2_Z01 g60922 ( .a(n_82), .b(pX_4_), .o(n_221) );
NAND2_Z01 g59686 ( .a(n_1380), .b(n_1332), .o(n_1450) );
BUF_X2 newInst_1225 ( .a(newNet_1224), .o(newNet_1225) );
BUF_X2 newInst_392 ( .a(newNet_391), .o(newNet_392) );
NAND2_Z01 g59502 ( .a(n_1543), .b(SP_10_), .o(n_1618) );
BUF_X2 newInst_199 ( .a(newNet_198), .o(newNet_199) );
fflopd pX_reg_0_ ( .CK(newNet_286), .D(n_2726), .Q(pX_0_) );
AND2_X1 g35363 ( .a(n_4488), .b(n_3286), .o(n_4631) );
BUF_X2 newInst_483 ( .a(newNet_141), .o(newNet_483) );
AND2_X1 g58256 ( .a(n_2752), .b(n_2214), .o(n_2811) );
NAND2_Z01 g34266 ( .a(n_4164), .b(pmem_d_8), .o(n_4267) );
BUF_X2 newInst_797 ( .a(newNet_796), .o(newNet_797) );
BUF_X2 newInst_299 ( .a(newNet_298), .o(newNet_299) );
BUF_X2 newInst_871 ( .a(newNet_870), .o(newNet_871) );
AND2_X1 g35087 ( .a(n_3488), .b(pZ_6_), .o(n_3508) );
NOR2_Z1 g34429 ( .a(n_4088), .b(n_3472), .o(n_4108) );
INV_X1 g35464 ( .a(pX_7_), .o(n_3260) );
XOR2_X1 g59595 ( .a(n_1452), .b(n_300), .o(n_1534) );
BUF_X2 newInst_1726 ( .a(newNet_1725), .o(newNet_1726) );
XOR2_X1 g58944 ( .a(n_2114), .b(n_1880), .o(n_2163) );
BUF_X2 newInst_725 ( .a(newNet_724), .o(newNet_725) );
NAND2_Z01 g34957 ( .a(n_3551), .b(GPR_7__1_), .o(n_3605) );
NAND3_Z1 g59248 ( .a(n_571), .b(n_1773), .c(n_41), .o(n_1867) );
XOR2_X1 g60392 ( .a(n_284), .b(n_149), .o(n_754) );
BUF_X2 newInst_1639 ( .a(newNet_1638), .o(newNet_1639) );
fflopd U_reg_5_ ( .CK(newNet_371), .D(n_3091), .Q(U_5_) );
INV_X1 g61099 ( .a(n_4634), .o(n_53) );
AND2_X1 g60331 ( .a(n_589), .b(n_65), .o(n_797) );
BUF_X2 newInst_1452 ( .a(newNet_585), .o(newNet_1452) );
NAND2_Z01 g35082 ( .a(n_3478), .b(n_4478), .o(n_3503) );
NOR2_Z1 g60987 ( .a(n_4449), .b(n_4433), .o(n_143) );
AND2_X1 g60069 ( .a(n_848), .b(n_36), .o(n_1065) );
NAND2_Z01 g60402 ( .a(n_457), .b(GPR_16__6_), .o(n_744) );
BUF_X2 newInst_714 ( .a(newNet_452), .o(newNet_714) );
BUF_X2 newInst_252 ( .a(newNet_251), .o(newNet_252) );
INV_X1 g61047 ( .a(PC_10_), .o(n_105) );
NOR4_Z1 g34129 ( .a(n_4235), .b(n_4233), .c(n_4320), .d(n_4130), .o(n_4379) );
NOR2_Z1 g35010 ( .a(n_3510), .b(n_3550), .o(n_3567) );
NAND2_Z01 g57715 ( .a(n_3124), .b(n_2345), .o(n_3152) );
fflopd GPR_reg_13__6_ ( .CK(newNet_1591), .D(n_3087), .Q(GPR_13__6_) );
NAND2_Z01 g59698 ( .a(io_do_5), .b(n_1384), .o(n_1432) );
BUF_X2 newInst_1340 ( .a(newNet_1339), .o(newNet_1340) );
BUF_X2 newInst_589 ( .a(newNet_588), .o(newNet_589) );
NOR2_Z1 g60609 ( .a(n_325), .b(n_169), .o(n_514) );
NAND2_Z01 g60902 ( .a(PC_5_), .b(pmem_d_5), .o(n_233) );
NOR2_Z1 g34913 ( .a(n_3562), .b(n_3215), .o(n_3650) );
NAND4_Z1 g58345 ( .a(n_1960), .b(n_2468), .c(n_2652), .d(n_2032), .o(n_2725) );
BUF_X2 newInst_1511 ( .a(newNet_1510), .o(newNet_1511) );
NAND2_Z01 final_adder_mux_R16_278_6_g390 ( .a(final_adder_mux_R16_278_6_n_57), .b(final_adder_mux_R16_278_6_n_14), .o(final_adder_mux_R16_278_6_n_59) );
NAND2_Z01 g60247 ( .a(n_508), .b(n_4478), .o(n_898) );
BUF_X2 newInst_305 ( .a(newNet_28), .o(newNet_305) );
fflopd io_sp_reg_1_ ( .CK(newNet_334), .D(n_549), .Q(io_sp_1_) );
XOR2_X1 g35378 ( .a(pX_1_), .b(pX_0_), .o(n_3344) );
NAND2_Z01 g58313 ( .a(n_2720), .b(n_1621), .o(n_2757) );
NOR2_Z1 g59358 ( .a(n_19), .b(n_1532), .o(n_1755) );
BUF_X2 newInst_1247 ( .a(newNet_1246), .o(newNet_1247) );
NOR2_Z1 g60365 ( .a(n_527), .b(n_509), .o(n_775) );
BUF_X2 newInst_842 ( .a(newNet_841), .o(newNet_842) );
fflopd Rd_r_reg_3_ ( .CK(newNet_584), .D(n_952), .Q(Rd_r_3_) );
NOR4_Z1 g34211 ( .a(n_3966), .b(n_3967), .c(n_4285), .d(n_3952), .o(n_4315) );
NAND2_Z01 g59779 ( .a(n_350), .b(n_1239), .o(n_1342) );
NAND2_Z01 g59468 ( .a(n_1585), .b(SP_7_), .o(n_1655) );
BUF_X2 newInst_268 ( .a(newNet_267), .o(newNet_268) );
BUF_X2 newInst_74 ( .a(newNet_73), .o(newNet_74) );
NOR2_Z1 g59560 ( .a(n_1472), .b(pmem_d_1), .o(n_1566) );
NOR2_Z1 g59951 ( .a(n_1121), .b(n_969), .o(n_1202) );
BUF_X2 newInst_791 ( .a(newNet_790), .o(newNet_791) );
BUF_X2 newInst_68 ( .a(newNet_67), .o(newNet_68) );
NAND2_Z01 g34884 ( .a(n_3564), .b(pX_3_), .o(n_3679) );
BUF_X2 newInst_938 ( .a(newNet_937), .o(newNet_938) );
BUF_X2 newInst_998 ( .a(newNet_997), .o(newNet_998) );
NOR2_Z1 g60707 ( .a(n_243), .b(n_4626), .o(n_431) );
BUF_X2 newInst_1490 ( .a(newNet_1489), .o(newNet_1490) );
BUF_X2 newInst_1443 ( .a(newNet_1442), .o(newNet_1443) );
INV_X2 newInst_798 ( .a(newNet_797), .o(newNet_798) );
BUF_X2 newInst_985 ( .a(newNet_984), .o(newNet_985) );
fflopd GPR_reg_17__7_ ( .CK(newNet_1378), .D(n_3162), .Q(GPR_17__7_) );
BUF_X2 newInst_1458 ( .a(newNet_1457), .o(newNet_1458) );
NOR3_Z1 g60121 ( .a(n_42), .b(n_489), .c(pmem_d_9), .o(n_1006) );
NAND2_Z01 final_adder_mux_R16_278_6_g401 ( .a(final_adder_mux_R16_278_6_n_46), .b(final_adder_mux_R16_278_6_n_10), .o(final_adder_mux_R16_278_6_n_48) );
BUF_X2 newInst_1501 ( .a(newNet_1500), .o(newNet_1501) );
NAND2_Z01 g34615 ( .a(n_3897), .b(n_3509), .o(n_3945) );
BUF_X2 newInst_1089 ( .a(newNet_1088), .o(newNet_1089) );
NOR3_Z1 g57849 ( .a(n_1419), .b(n_2994), .c(n_1905), .o(n_3063) );
BUF_X2 newInst_2 ( .a(newNet_1), .o(newNet_2) );
NAND2_Z01 g34113 ( .a(io_do_7), .b(n_4177), .o(n_4386) );
NAND3_Z1 g58702 ( .a(n_4644), .b(n_2151), .c(n_4682), .o(n_2442) );
NAND2_Z01 g58282 ( .a(n_2713), .b(n_1158), .o(n_2788) );
NAND2_Z01 g59319 ( .a(n_4), .b(n_4553), .o(n_1794) );
BUF_X2 newInst_1184 ( .a(newNet_1183), .o(newNet_1184) );
BUF_X2 newInst_294 ( .a(newNet_293), .o(newNet_294) );
AND2_X1 g57994 ( .a(n_2940), .b(n_2214), .o(n_2977) );
INV_X1 g35094 ( .a(n_4569), .o(n_3498) );
NAND2_Z01 g34303 ( .a(n_4166), .b(n_4543), .o(n_4231) );
BUF_X2 newInst_527 ( .a(newNet_526), .o(newNet_527) );
NOR2_Z1 g35115 ( .a(n_3202), .b(pmem_d_3), .o(n_4472) );
NOR3_Z1 g34494 ( .a(n_4007), .b(n_3981), .c(n_4019), .o(n_4050) );
INV_X1 g34984 ( .a(n_3561), .o(n_4602) );
AND2_X1 g58250 ( .a(n_2752), .b(n_2159), .o(n_2817) );
BUF_X2 newInst_156 ( .a(newNet_155), .o(newNet_156) );
INV_X1 g59778 ( .a(n_1343), .o(n_1344) );
NAND2_Z02 g58958 ( .a(n_2115), .b(n_1213), .o(n_2158) );
BUF_X2 newInst_1747 ( .a(newNet_1746), .o(newNet_1747) );
BUF_X2 newInst_737 ( .a(newNet_736), .o(newNet_737) );
AND2_X1 g60583 ( .a(n_61), .b(n_459), .o(n_529) );
NAND2_Z01 g58494 ( .a(n_2571), .b(n_1838), .o(n_2603) );
NAND2_Z01 g58325 ( .a(n_2669), .b(n_2319), .o(n_2740) );
NOR2_Z1 g34609 ( .a(n_3692), .b(n_3660), .o(n_3951) );
BUF_X2 newInst_1200 ( .a(newNet_1199), .o(newNet_1200) );
NOR2_Z1 g60975 ( .a(n_4439), .b(n_4423), .o(n_193) );
AND2_X1 g60630 ( .a(n_459), .b(n_199), .o(n_581) );
NAND2_Z01 g57702 ( .a(n_3140), .b(n_2185), .o(n_3167) );
INV_X2 newInst_563 ( .a(newNet_562), .o(newNet_563) );
NAND2_Z01 g59225 ( .a(n_1851), .b(n_166), .o(n_1897) );
BUF_X2 newInst_1257 ( .a(newNet_1256), .o(newNet_1257) );
BUF_X2 newInst_1173 ( .a(newNet_1172), .o(newNet_1173) );
BUF_X2 newInst_1836 ( .a(newNet_888), .o(newNet_1836) );
NOR2_Z1 g60588 ( .a(n_332), .b(n_181), .o(n_525) );
INV_X1 g35466 ( .a(pZ_9_), .o(n_3258) );
BUF_X2 newInst_1091 ( .a(newNet_1090), .o(newNet_1091) );
NAND2_Z01 g34705 ( .a(n_3631), .b(GPR_11__6_), .o(n_3860) );
NAND2_Z01 g58586 ( .a(n_2462), .b(pY_13_), .o(n_2512) );
BUF_X2 newInst_142 ( .a(newNet_3), .o(newNet_142) );
NAND2_Z01 g59633 ( .a(n_1422), .b(SP_1_), .o(n_1496) );
INV_X1 g61035 ( .a(PC_1_), .o(n_117) );
BUF_X2 newInst_1667 ( .a(newNet_1666), .o(newNet_1667) );
BUF_X2 newInst_1571 ( .a(newNet_1570), .o(newNet_1571) );
NOR2_Z1 g60932 ( .a(n_32), .b(pmem_d_12), .o(n_257) );
NAND2_Z01 g35273 ( .a(n_3289), .b(pY_13_), .o(n_3402) );
NAND2_Z01 g59925 ( .a(n_178), .b(n_1049), .o(n_1192) );
AND2_X1 g58260 ( .a(n_2752), .b(n_2210), .o(n_2807) );
NAND2_Z01 g58695 ( .a(n_2210), .b(GPR_1__2_), .o(n_2411) );
NAND2_Z01 g58129 ( .a(n_2849), .b(n_24), .o(n_2908) );
NAND4_Z1 g60150 ( .a(n_635), .b(n_737), .c(n_560), .d(n_691), .o(n_983) );
NAND2_Z01 g34893 ( .a(n_3590), .b(pY_12_), .o(n_3670) );
AND2_X1 g57751 ( .a(n_3115), .b(n_2200), .o(n_3120) );
NOR2_Z1 g35117 ( .a(n_3205), .b(pmem_d_2), .o(n_4473) );
BUF_X2 newInst_868 ( .a(newNet_867), .o(newNet_868) );
BUF_X2 newInst_134 ( .a(newNet_30), .o(newNet_134) );
NOR4_Z1 g59803 ( .a(n_1221), .b(n_1006), .c(n_4556), .d(n_1005), .o(n_1325) );
NAND2_Z01 g34941 ( .a(n_3552), .b(GPR_0__6_), .o(n_3621) );
NAND3_Z1 g57650 ( .a(n_2562), .b(n_3175), .c(n_2149), .o(n_3192) );
BUF_X2 newInst_1464 ( .a(newNet_1463), .o(newNet_1464) );
NAND2_Z01 g59946 ( .a(n_1018), .b(n_223), .o(n_1180) );
BUF_X2 newInst_231 ( .a(newNet_230), .o(newNet_231) );
BUF_X2 newInst_513 ( .a(newNet_512), .o(newNet_513) );
BUF_X2 newInst_181 ( .a(newNet_180), .o(newNet_181) );
NAND2_Z01 g34847 ( .a(n_3627), .b(GPR_15__1_), .o(n_3716) );
BUF_X2 newInst_1231 ( .a(newNet_1230), .o(newNet_1231) );
BUF_X2 newInst_605 ( .a(newNet_604), .o(newNet_605) );
BUF_X2 newInst_300 ( .a(newNet_299), .o(newNet_300) );
BUF_X2 newInst_1404 ( .a(newNet_1403), .o(newNet_1404) );
BUF_X2 newInst_361 ( .a(newNet_360), .o(newNet_361) );
NAND2_Z01 g58867 ( .a(n_2157), .b(GPR_13__7_), .o(n_2240) );
BUF_X2 newInst_1843 ( .a(newNet_1842), .o(newNet_1843) );
NAND2_Z01 g58154 ( .a(n_2811), .b(n_2415), .o(n_2859) );
NAND3_Z1 g58565 ( .a(n_1785), .b(n_2489), .c(n_1087), .o(n_2533) );
NOR4_Z1 g59772 ( .a(n_510), .b(n_294), .c(n_1153), .d(n_470), .o(n_1357) );
BUF_X2 newInst_1049 ( .a(newNet_1048), .o(newNet_1049) );
NAND2_Z01 g58684 ( .a(n_2211), .b(GPR_19__0_), .o(n_2422) );
NOR3_Z1 g59186 ( .a(n_1818), .b(n_1408), .c(n_793), .o(n_1921) );
NAND2_Z01 g60323 ( .a(n_597), .b(pX_14_), .o(n_804) );
NAND2_Z01 g57658 ( .a(n_3172), .b(n_2298), .o(n_3184) );
NAND2_Z01 g34220 ( .a(n_4294), .b(SP_11_), .o(n_4307) );
BUF_X2 newInst_463 ( .a(newNet_462), .o(newNet_463) );
NOR2_Z1 g60644 ( .a(n_460), .b(n_199), .o(n_574) );
NAND2_Z01 g58876 ( .a(n_2153), .b(GPR_8__2_), .o(n_2231) );
BUF_X2 newInst_1505 ( .a(newNet_953), .o(newNet_1505) );
INV_X1 g60536 ( .a(n_592), .o(n_593) );
NAND2_Z01 g58806 ( .a(n_2197), .b(U_4_), .o(n_2294) );
NAND2_Z01 g58784 ( .a(n_2199), .b(GPR_0__0_), .o(n_2316) );
NAND2_Z01 final_adder_mux_R16_278_6_g422 ( .a(n_4447), .b(n_4431), .o(final_adder_mux_R16_278_6_n_26) );
NOR2_Z1 g59958 ( .a(n_987), .b(n_1017), .o(n_1174) );
BUF_X1 drc_bufs61250 ( .a(n_2170), .o(n_1) );
NOR2_Z1 g34285 ( .a(n_4163), .b(n_3225), .o(n_4248) );
NOR2_Z1 g59691 ( .a(n_1373), .b(n_1022), .o(n_1445) );
INV_X1 g61068 ( .a(PC_9_), .o(n_84) );
NAND2_Z01 g61015 ( .a(n_87), .b(n_48), .o(n_167) );
NAND2_Z01 g34670 ( .a(n_3600), .b(n_3612), .o(n_3895) );
XNOR2_X1 g59812 ( .a(n_1159), .b(pmem_d_9), .o(n_1317) );
BUF_X2 newInst_666 ( .a(newNet_56), .o(newNet_666) );
NAND2_Z01 g60749 ( .a(n_203), .b(SP_1_), .o(n_393) );
XOR2_X1 g60159 ( .a(n_576), .b(n_64), .o(n_1025) );
INV_X2 newInst_1080 ( .a(newNet_1079), .o(newNet_1080) );
XOR2_X1 final_adder_mux_R16_278_6_g415 ( .a(n_4436), .b(n_4420), .o(final_adder_mux_R16_278_6_n_34) );
NAND2_Z01 g60425 ( .a(n_368), .b(GPR_13__2_), .o(n_721) );
NOR3_Z1 g59660 ( .a(n_988), .b(n_1319), .c(n_956), .o(n_1466) );
AND2_X1 g35303 ( .a(n_4561), .b(n_3227), .o(n_3413) );
BUF_X2 newInst_129 ( .a(newNet_128), .o(newNet_129) );
BUF_X2 newInst_343 ( .a(newNet_196), .o(newNet_343) );
XOR2_X1 g60784 ( .a(PC_3_), .b(pmem_d_6), .o(n_319) );
NAND2_Z01 g60939 ( .a(io_do_1), .b(n_35), .o(n_212) );
NAND4_Z1 g58178 ( .a(n_2732), .b(n_2716), .c(n_2174), .d(n_1404), .o(n_2835) );
BUF_X2 newInst_805 ( .a(newNet_804), .o(newNet_805) );
NAND3_Z1 g58484 ( .a(n_480), .b(n_2569), .c(n_4485), .o(n_2612) );
fflopd GPR_reg_21__7_ ( .CK(newNet_1113), .D(n_3155), .Q(GPR_21__7_) );
NAND2_Z01 g58465 ( .a(n_2422), .b(n_2592), .o(n_2631) );
NOR2_Z1 g60882 ( .a(n_57), .b(n_35), .o(n_243) );
NAND2_Z01 g35317 ( .a(n_3289), .b(pY_5_), .o(n_3361) );
NAND2_Z01 g58620 ( .a(n_2354), .b(pX_1_), .o(n_2477) );
BUF_X2 newInst_53 ( .a(newNet_52), .o(newNet_53) );
BUF_X2 newInst_114 ( .a(newNet_113), .o(newNet_114) );
NAND2_Z01 g60474 ( .a(n_371), .b(GPR_21__3_), .o(n_672) );
NAND4_Z1 g59993 ( .a(n_924), .b(n_889), .c(n_936), .d(n_930), .o(n_1136) );
BUF_X2 newInst_1602 ( .a(newNet_1601), .o(newNet_1602) );
BUF_X2 newInst_680 ( .a(newNet_679), .o(newNet_680) );
NAND3_Z1 g60657 ( .a(n_238), .b(n_137), .c(n_4641), .o(n_569) );
NOR2_Z1 g34268 ( .a(n_4163), .b(n_3244), .o(n_4265) );
NAND2_Z01 g58333 ( .a(n_929), .b(n_2690), .o(n_2756) );
NAND4_Z1 g58934 ( .a(n_1691), .b(n_1794), .c(n_2121), .d(n_1643), .o(n_2173) );
NAND2_Z01 g59076 ( .a(n_1896), .b(n_4527), .o(n_2031) );
fflopd GPR_reg_19__4_ ( .CK(newNet_1295), .D(n_2936), .Q(GPR_19__4_) );
NAND2_Z01 g34161 ( .a(n_4317), .b(pmem_d_3), .o(n_4347) );
NAND2_Z01 g59070 ( .a(n_1871), .b(n_4603), .o(n_2037) );
BUF_X2 newInst_674 ( .a(newNet_673), .o(newNet_674) );
NOR2_Z1 g34992 ( .a(n_3535), .b(n_3484), .o(n_3590) );
NAND4_Z1 g60376 ( .a(n_442), .b(n_440), .c(n_428), .d(n_439), .o(n_768) );
NOR2_Z1 g35008 ( .a(n_3510), .b(n_3535), .o(n_3568) );
XNOR2_X1 g58990 ( .a(n_2060), .b(n_1880), .o(n_2118) );
NOR2_Z1 g60357 ( .a(n_602), .b(PC_4_), .o(n_851) );
BUF_X2 newInst_551 ( .a(newNet_550), .o(newNet_551) );
NAND2_Z01 g58240 ( .a(n_2753), .b(n_2193), .o(n_2827) );
fflopd pZ_reg_8_ ( .CK(newNet_47), .D(n_2723), .Q(pZ_8_) );
NAND2_Z01 g58636 ( .a(n_2360), .b(pY_3_), .o(n_2466) );
NAND2_Z01 g58963 ( .a(n_2084), .b(n_1209), .o(n_2142) );
NAND2_Z01 g60710 ( .a(n_198), .b(GPR_20__1_), .o(n_428) );
NAND2_Z01 g58761 ( .a(n_2203), .b(GPR_4__5_), .o(n_2339) );
BUF_X2 newInst_1754 ( .a(newNet_1753), .o(newNet_1754) );
BUF_X2 newInst_1125 ( .a(newNet_1124), .o(newNet_1125) );
NAND4_Z1 g34570 ( .a(n_3682), .b(n_3836), .c(n_3665), .d(n_3837), .o(n_3990) );
NAND3_Z1 g58829 ( .a(n_1793), .b(n_2171), .c(n_1091), .o(n_2278) );
NAND2_Z01 g59624 ( .a(n_1413), .b(io_sp_5_), .o(n_1503) );
INV_X2 g61108 ( .a(pmem_d_2), .o(n_44) );
BUF_X2 newInst_1146 ( .a(newNet_1145), .o(newNet_1146) );
fflopd pY_reg_15_ ( .CK(newNet_166), .D(n_3191), .Q(pY_15_) );
NAND2_Z01 g60786 ( .a(n_192), .b(n_265), .o(n_379) );
BUF_X2 newInst_318 ( .a(newNet_317), .o(newNet_318) );
NAND3_Z1 g59987 ( .a(n_142), .b(n_790), .c(n_163), .o(n_1142) );
NAND2_Z01 g58893 ( .a(n_2140), .b(GPR_9__7_), .o(n_2189) );
NOR4_Z1 g58936 ( .a(n_1757), .b(n_1783), .c(n_1992), .d(n_1642), .o(n_2171) );
INV_X1 drc_bufs61134 ( .a(n_1415), .o(n_16) );
BUF_X2 newInst_1699 ( .a(newNet_127), .o(newNet_1699) );
BUF_X2 newInst_1308 ( .a(newNet_1307), .o(newNet_1308) );
NAND2_Z01 g35135 ( .a(Rd_1_), .b(n_3232), .o(n_3482) );
NAND2_Z01 g34746 ( .a(n_3628), .b(GPR_19__1_), .o(n_3819) );
NAND2_Z01 g34649 ( .a(n_3768), .b(n_4547), .o(n_3911) );
NAND2_Z01 g58548 ( .a(n_2523), .b(pY_12_), .o(n_2549) );
NAND2_Z01 g59823 ( .a(n_1171), .b(dmem_di_3), .o(n_1301) );
NAND2_Z01 g34522 ( .a(n_3663), .b(n_3946), .o(n_4021) );
BUF_X2 newInst_477 ( .a(newNet_476), .o(newNet_477) );
BUF_X2 newInst_381 ( .a(newNet_380), .o(newNet_381) );
NAND2_Z01 g34958 ( .a(n_3552), .b(GPR_11__0_), .o(n_3604) );
NAND2_Z01 g58627 ( .a(n_2362), .b(n_1682), .o(n_2471) );
AND3_X1 g59041 ( .a(n_49), .b(n_1982), .c(pZ_11_), .o(n_2068) );
INV_X1 g59382 ( .a(n_1733), .o(n_1734) );
BUF_X2 newInst_544 ( .a(newNet_70), .o(newNet_544) );
NAND4_Z1 g59539 ( .a(n_1184), .b(n_1515), .c(n_1514), .d(n_1236), .o(n_1589) );
NAND2_Z01 g60290 ( .a(R16_8_), .b(n_14), .o(n_834) );
BUF_X2 newInst_506 ( .a(newNet_505), .o(newNet_506) );
fflopd GPR_reg_21__6_ ( .CK(newNet_1118), .D(n_3075), .Q(GPR_21__6_) );
NOR2_Z1 g59868 ( .a(n_1219), .b(n_458), .o(n_1259) );
NAND2_Z01 g34203 ( .a(io_do_6), .b(n_4177), .o(n_4323) );
NAND2_Z01 g34729 ( .a(n_3592), .b(GPR_22__5_), .o(n_3836) );
INV_X1 g60095 ( .a(n_1027), .o(n_1028) );
BUF_X2 newInst_645 ( .a(newNet_644), .o(newNet_645) );
NAND2_Z01 g60234 ( .a(n_596), .b(GPR_3__0_), .o(n_911) );
NAND2_Z01 g60619 ( .a(n_155), .b(n_383), .o(n_508) );
INV_X1 g60172 ( .a(n_961), .o(n_960) );
NAND2_Z01 g60022 ( .a(n_932), .b(n_917), .o(n_1105) );
BUF_X2 newInst_789 ( .a(newNet_788), .o(newNet_789) );
BUF_X2 newInst_556 ( .a(newNet_118), .o(newNet_556) );
INV_X1 g58615 ( .a(n_2478), .o(n_2479) );
INV_X1 g58745 ( .a(n_2361), .o(n_2360) );
BUF_X2 newInst_63 ( .a(newNet_62), .o(newNet_63) );
NAND2_Z01 final_adder_mux_R16_278_6_g429 ( .a(n_4451), .b(n_4435), .o(final_adder_mux_R16_278_6_n_28) );
INV_X1 g60947 ( .a(n_204), .o(n_203) );
INV_X1 g59556 ( .a(n_1568), .o(n_1569) );
XOR2_X1 g34463 ( .a(n_4056), .b(pY_9_), .o(n_4079) );
AND2_X1 g59689 ( .a(n_1349), .b(n_112), .o(n_1446) );
BUF_X2 newInst_929 ( .a(newNet_928), .o(newNet_929) );
BUF_X2 newInst_922 ( .a(newNet_921), .o(newNet_922) );
AND3_X1 g35240 ( .a(n_4668), .b(n_4684), .c(n_3292), .o(n_4667) );
NOR2_Z1 g35164 ( .a(n_3425), .b(pmem_d_3), .o(n_3465) );
NAND2_Z01 g34691 ( .a(n_3591), .b(U_15_), .o(n_3874) );
NAND4_Z1 g59448 ( .a(n_777), .b(n_1477), .c(n_1612), .d(n_1359), .o(n_1674) );
NAND2_Z01 g60494 ( .a(n_349), .b(U_5_), .o(n_652) );
XOR2_X1 g35144 ( .a(n_3427), .b(pY_4_), .o(n_3475) );
NAND2_Z01 g58718 ( .a(n_2208), .b(GPR_21__7_), .o(n_2389) );
NAND2_Z01 g34097 ( .a(n_4369), .b(n_4368), .o(n_4439) );
NOR2_Z1 g60622 ( .a(n_365), .b(S), .o(n_506) );
NAND2_Z01 g60433 ( .a(n_358), .b(GPR_0__2_), .o(n_713) );
NAND2_Z01 g60482 ( .a(Rd_0_), .b(n_340), .o(n_664) );
BUF_X2 newInst_1482 ( .a(newNet_1481), .o(newNet_1482) );
BUF_X2 newInst_992 ( .a(newNet_801), .o(newNet_992) );
NAND4_Z1 g57911 ( .a(n_2070), .b(n_2549), .c(n_2989), .d(n_2050), .o(n_3028) );
BUF_X2 newInst_962 ( .a(newNet_961), .o(newNet_962) );
BUF_X2 newInst_401 ( .a(newNet_400), .o(newNet_401) );
NAND2_Z01 g58997 ( .a(n_1978), .b(n_4635), .o(n_2110) );
XOR2_X1 g60164 ( .a(n_618), .b(n_298), .o(n_972) );
INV_X1 g59281 ( .a(n_1832), .o(n_1833) );
NOR2_Z1 g60794 ( .a(n_248), .b(n_250), .o(n_372) );
NAND2_Z01 g34817 ( .a(n_3627), .b(GPR_15__2_), .o(n_3746) );
BUF_X2 newInst_1782 ( .a(newNet_1149), .o(newNet_1782) );
NAND2_Z01 g59831 ( .a(n_1216), .b(n_157), .o(n_1294) );
NAND2_Z01 g60350 ( .a(n_576), .b(n_64), .o(n_859) );
NOR4_Z1 g34459 ( .a(n_3846), .b(n_3965), .c(n_4046), .d(n_3702), .o(n_4083) );
AND2_X1 g59428 ( .a(n_1646), .b(n_4553), .o(n_1691) );
INV_X1 g34799 ( .a(n_4598), .o(n_3764) );
BUF_X2 newInst_423 ( .a(newNet_422), .o(newNet_423) );
BUF_X2 newInst_202 ( .a(newNet_126), .o(newNet_202) );
NOR2_Z1 g60958 ( .a(n_4626), .b(n_62), .o(n_159) );
BUF_X2 newInst_635 ( .a(newNet_634), .o(newNet_635) );
NAND2_Z01 g60755 ( .a(io_do_0), .b(n_261), .o(n_464) );
NAND2_Z01 final_adder_mux_R16_278_6_g383 ( .a(final_adder_mux_R16_278_6_n_65), .b(final_adder_mux_R16_278_6_n_2), .o(final_adder_mux_R16_278_6_n_66) );
BUF_X2 newInst_30 ( .a(newNet_29), .o(newNet_30) );
NOR4_Z1 g34241 ( .a(n_4023), .b(n_4034), .c(n_4169), .d(n_3869), .o(n_4292) );
BUF_X2 newInst_1040 ( .a(newNet_1039), .o(newNet_1040) );
NAND2_Z01 g34703 ( .a(n_3581), .b(GPR_16__7_), .o(n_3862) );
NAND2_Z01 g58732 ( .a(n_2206), .b(GPR_23__5_), .o(n_2375) );
NAND2_Z01 g59156 ( .a(n_1896), .b(n_1205), .o(n_1982) );
NAND2_Z01 g58577 ( .a(n_2471), .b(n_1710), .o(n_2526) );
BUF_X2 newInst_846 ( .a(newNet_845), .o(newNet_846) );
NOR2_Z1 g34312 ( .a(n_16064_BAR), .b(n_3532), .o(n_4221) );
BUF_X2 newInst_1427 ( .a(newNet_1426), .o(newNet_1427) );
BUF_X2 newInst_1415 ( .a(newNet_1414), .o(newNet_1415) );
NOR2_Z3 g34209 ( .a(n_4556), .b(pmem_d_8), .o(n_4317) );
BUF_X2 newInst_1274 ( .a(newNet_1273), .o(newNet_1274) );
BUF_X2 newInst_1333 ( .a(newNet_1332), .o(newNet_1333) );
BUF_X2 newInst_1381 ( .a(newNet_874), .o(newNet_1381) );
NAND2_Z01 g60752 ( .a(SP_8_), .b(n_180), .o(n_390) );
NAND2_Z01 g59786 ( .a(n_1268), .b(n_1046), .o(n_1338) );
NOR2_Z1 g35000 ( .a(n_3490), .b(n_3548), .o(n_3581) );
BUF_X2 newInst_720 ( .a(newNet_719), .o(newNet_720) );
AND2_X1 g58397 ( .a(n_2657), .b(n_2201), .o(n_2671) );
BUF_X2 newInst_1051 ( .a(newNet_1050), .o(newNet_1051) );
BUF_X2 newInst_439 ( .a(newNet_438), .o(newNet_439) );
NAND2_Z01 g58862 ( .a(n_2156), .b(GPR_15__0_), .o(n_2245) );
NAND2_Z01 final_adder_mux_R16_278_6_g433 ( .a(n_4450), .b(n_4434), .o(final_adder_mux_R16_278_6_n_16) );
NAND2_Z01 g35333 ( .a(pZ_7_), .b(n_3199), .o(n_3337) );
NAND2_Z01 g58755 ( .a(n_2204), .b(GPR_3__7_), .o(n_2345) );
NAND2_Z01 final_adder_mux_R16_278_6_g380 ( .a(final_adder_mux_R16_278_6_n_68), .b(final_adder_mux_R16_278_6_n_3), .o(final_adder_mux_R16_278_6_n_69) );
BUF_X2 newInst_209 ( .a(newNet_208), .o(newNet_209) );
INV_X1 drc_bufs61147 ( .a(n_1619), .o(n_27) );
NAND2_Z01 g59055 ( .a(n_1902), .b(n_4586), .o(n_2052) );
NOR2_Z1 g34341 ( .a(n_4178), .b(n_4078), .o(n_4193) );
NAND2_Z01 g59700 ( .a(io_do_2), .b(n_1384), .o(n_1430) );
fflopd GPR_reg_13__2_ ( .CK(newNet_1607), .D(n_2780), .Q(GPR_13__2_) );
NAND2_Z01 g58881 ( .a(n_2156), .b(GPR_15__4_), .o(n_2226) );
NAND2_Z01 g59747 ( .a(n_1306), .b(n_234), .o(n_1375) );
BUF_X2 newInst_1489 ( .a(newNet_1488), .o(newNet_1489) );
NAND2_Z01 g58166 ( .a(n_2800), .b(n_2341), .o(n_2844) );
AND2_X1 g58387 ( .a(n_2656), .b(n_2206), .o(n_2681) );
BUF_X2 newInst_1237 ( .a(newNet_1236), .o(newNet_1237) );
NAND4_Z2 g35191 ( .a(n_3339), .b(n_3375), .c(n_3366), .d(n_3392), .o(n_4625) );
AND3_X1 g60848 ( .a(pmem_d_3), .b(n_4651), .c(pmem_d_2), .o(n_338) );
NOR2_Z1 g60733 ( .a(n_217), .b(n_42), .o(n_406) );
BUF_X2 newInst_1556 ( .a(newNet_1555), .o(newNet_1556) );
BUF_X2 newInst_273 ( .a(newNet_246), .o(newNet_273) );
NAND2_Z01 g58740 ( .a(n_2205), .b(GPR_2__5_), .o(n_2367) );
AND2_X1 g58115 ( .a(n_2850), .b(n_2209), .o(n_2897) );
BUF_X2 newInst_1773 ( .a(newNet_1772), .o(newNet_1773) );
NAND4_Z1 g59551 ( .a(n_1149), .b(n_1370), .c(n_1492), .d(n_1054), .o(n_1577) );
NAND2_Z01 g57881 ( .a(n_3010), .b(n_2216), .o(n_3058) );
NAND2_Z01 g61006 ( .a(n_83), .b(n_59), .o(n_133) );
BUF_X2 newInst_51 ( .a(newNet_50), .o(newNet_51) );
NAND2_Z01 g35283 ( .a(U_9_), .b(n_3275), .o(n_3392) );
BUF_X2 newInst_329 ( .a(newNet_328), .o(newNet_329) );
NOR3_Z1 g60667 ( .a(n_277), .b(n_4556), .c(n_32), .o(n_566) );
AND2_X1 g35369 ( .a(n_3301), .b(n_3272), .o(n_3321) );
NAND2_Z01 g34951 ( .a(n_3549), .b(U_4_), .o(n_3611) );
NAND2_Z01 g35027 ( .a(n_3528), .b(n_3281), .o(n_3542) );
NAND2_Z01 g58729 ( .a(n_2206), .b(GPR_23__2_), .o(n_2378) );
NAND2_Z01 g34261 ( .a(n_4176), .b(pX_12_), .o(n_4272) );
NAND2_Z01 g34835 ( .a(n_3581), .b(GPR_16__1_), .o(n_3728) );
NAND2_Z01 g34841 ( .a(n_3597), .b(GPR_17__1_), .o(n_3722) );
XOR2_X1 g59900 ( .a(n_1048), .b(io_do_6), .o(n_1266) );
NOR2_Z1 g35252 ( .a(n_3316), .b(pY_10_), .o(n_4518) );
NAND2_Z01 g58054 ( .a(n_2890), .b(n_2340), .o(n_2928) );
NAND2_Z01 g58167 ( .a(n_2799), .b(n_2333), .o(n_2843) );
INV_X2 newInst_1550 ( .a(newNet_948), .o(newNet_1550) );
BUF_X2 newInst_741 ( .a(newNet_740), .o(newNet_741) );
NAND2_Z01 g59616 ( .a(n_17), .b(V), .o(n_1511) );
BUF_X2 newInst_1848 ( .a(newNet_1847), .o(newNet_1848) );
BUF_X2 newInst_655 ( .a(newNet_654), .o(newNet_655) );
INV_X1 g35491 ( .a(U_3_), .o(n_3234) );
fflopd GPR_reg_1__7_ ( .CK(newNet_1214), .D(n_3159), .Q(GPR_1__7_) );
NOR2_Z1 g59271 ( .a(n_1777), .b(n_1653), .o(n_1841) );
NOR2_Z1 g60990 ( .a(n_4437), .b(n_4421), .o(n_181) );
NOR2_Z1 g34840 ( .a(n_3583), .b(n_4401), .o(n_3723) );
NAND2_Z01 g58274 ( .a(n_2729), .b(n_25), .o(n_2793) );
BUF_X2 newInst_703 ( .a(newNet_702), .o(newNet_703) );
NOR2_Z1 g60346 ( .a(n_747), .b(n_534), .o(n_785) );
NAND2_Z01 g60459 ( .a(n_371), .b(GPR_21__2_), .o(n_687) );
NAND2_Z01 final_adder_mux_R16_278_6_g389 ( .a(final_adder_mux_R16_278_6_n_59), .b(final_adder_mux_R16_278_6_n_7), .o(final_adder_mux_R16_278_6_n_60) );
AND2_X1 g58541 ( .a(n_2536), .b(n_1188), .o(n_2557) );
NOR3_Z1 g59592 ( .a(n_839), .b(n_1491), .c(n_205), .o(n_1546) );
NOR2_Z1 g60592 ( .a(n_373), .b(pX_13_), .o(n_606) );
AND2_X1 g57886 ( .a(n_3009), .b(n_2139), .o(n_3052) );
NAND3_Z1 g34547 ( .a(n_3873), .b(n_3875), .c(n_3874), .o(n_4011) );
AND2_X1 g58356 ( .a(n_2657), .b(n_2159), .o(n_2715) );
AND2_X1 g34654 ( .a(n_3641), .b(state_2_), .o(n_3906) );
BUF_X2 newInst_1789 ( .a(newNet_1788), .o(newNet_1789) );
NAND2_Z01 g60210 ( .a(n_596), .b(GPR_3__3_), .o(n_935) );
INV_X1 g35423 ( .a(n_3287), .o(n_4653) );
NAND4_Z1 g34596 ( .a(n_3674), .b(n_3698), .c(n_3647), .d(n_3699), .o(n_3964) );
NOR2_Z1 g60256 ( .a(n_583), .b(n_92), .o(n_890) );
INV_X1 g35024 ( .a(n_3549), .o(n_3548) );
BUF_X2 newInst_144 ( .a(newNet_143), .o(newNet_144) );
NAND2_Z01 g35454 ( .a(n_4597), .b(n_3261), .o(n_3276) );
NAND2_Z01 g34874 ( .a(n_3572), .b(GPR_4__7_), .o(n_3689) );
BUF_X2 newInst_911 ( .a(newNet_910), .o(newNet_911) );
NAND2_Z01 g58320 ( .a(n_2675), .b(n_2342), .o(n_2745) );
AND2_X1 g59883 ( .a(n_1157), .b(n_1169), .o(n_1244) );
INV_X1 g61089 ( .a(io_do_2), .o(n_63) );
NOR2_Z1 g59344 ( .a(io_do_0), .b(n_1695), .o(n_1800) );
BUF_X2 newInst_987 ( .a(newNet_986), .o(newNet_987) );
NAND2_Z01 g34867 ( .a(n_3629), .b(GPR_3__0_), .o(n_3696) );
NAND2_Z01 g58247 ( .a(n_2754), .b(n_2198), .o(n_2820) );
XOR2_X1 g35051 ( .a(n_3506), .b(n_3210), .o(n_4590) );
NOR2_Z1 g60637 ( .a(n_458), .b(n_197), .o(n_578) );
XOR2_X1 g34480 ( .a(n_4037), .b(pZ_8_), .o(n_4062) );
XOR2_X1 g59905 ( .a(n_1110), .b(io_do_6), .o(n_1265) );
NAND2_Z01 g60209 ( .a(n_591), .b(GPR_22__2_), .o(n_936) );
AND3_X1 g59543 ( .a(n_1335), .b(n_1573), .c(n_309), .o(n_1585) );
BUF_X2 newInst_200 ( .a(newNet_199), .o(newNet_200) );
NAND2_Z01 g60524 ( .a(n_20), .b(Rd_r_4_), .o(n_622) );
NAND2_Z01 g58855 ( .a(n_2157), .b(GPR_13__3_), .o(n_2252) );
NAND2_Z01 g60489 ( .a(n_353), .b(GPR_10__4_), .o(n_657) );
AND2_X1 g35312 ( .a(n_4637), .b(n_3262), .o(n_3412) );
NAND2_Z01 g35217 ( .a(n_4526), .b(pZ_11_), .o(n_4527) );
XOR2_X1 g58570 ( .a(n_2482), .b(n_1770), .o(n_2528) );
NAND2_Z01 g59090 ( .a(n_1875), .b(n_4562), .o(n_2017) );
BUF_X2 newInst_1566 ( .a(newNet_1565), .o(newNet_1566) );
NAND2_Z01 g34387 ( .a(n_4085), .b(Rd_0_), .o(n_4150) );
NAND2_Z01 g60569 ( .a(n_468), .b(pY_3_), .o(n_615) );
INV_X1 g60284 ( .a(n_845), .o(n_846) );
NAND2_Z01 g59144 ( .a(n_1894), .b(n_1180), .o(n_1955) );
BUF_X2 newInst_249 ( .a(newNet_248), .o(newNet_249) );
NAND3_Z1 g34442 ( .a(n_3649), .b(n_4048), .c(n_3743), .o(n_4097) );
NAND2_Z01 g60181 ( .a(n_672), .b(n_675), .o(n_959) );
BUF_X2 newInst_1032 ( .a(newNet_1031), .o(newNet_1032) );
BUF_X2 newInst_492 ( .a(newNet_491), .o(newNet_492) );
NAND2_Z01 g34791 ( .a(n_3625), .b(GPR_1__3_), .o(n_3774) );
XOR2_X1 g34658 ( .a(n_3595), .b(pZ_10_), .o(n_3928) );
NOR4_Z1 g35071 ( .a(n_3444), .b(n_3417), .c(n_3456), .d(n_3347), .o(n_3516) );
NAND4_Z1 g58822 ( .a(n_1717), .b(n_1790), .c(n_2168), .d(n_1639), .o(n_2283) );
BUF_X2 newInst_834 ( .a(newNet_346), .o(newNet_834) );
INV_X1 g35507 ( .a(pmem_d_13), .o(n_3220) );
NAND2_Z01 g57942 ( .a(n_2965), .b(n_2331), .o(n_3000) );
XOR2_X1 g60385 ( .a(n_281), .b(n_131), .o(n_761) );
NOR2_Z1 g35036 ( .a(n_3522), .b(n_3350), .o(n_3544) );
NAND2_Z01 g59407 ( .a(io_do_7), .b(n_1661), .o(n_1735) );
XOR2_X1 final_adder_mux_R16_278_6_g407 ( .a(n_4444), .b(n_4428), .o(final_adder_mux_R16_278_6_n_42) );
NAND2_Z01 g58550 ( .a(n_2522), .b(pZ_12_), .o(n_2547) );
NAND2_Z01 g57984 ( .a(n_2941), .b(n_2216), .o(n_2988) );
XOR2_X1 g35103 ( .a(n_4618), .b(n_3251), .o(n_4465) );
NAND4_Z1 g59441 ( .a(n_812), .b(n_810), .c(n_1599), .d(n_921), .o(n_1679) );
BUF_X2 newInst_1709 ( .a(newNet_1708), .o(newNet_1709) );
BUF_X2 newInst_261 ( .a(newNet_260), .o(newNet_261) );
NAND4_Z1 g60138 ( .a(n_536), .b(n_732), .c(n_734), .d(n_705), .o(n_994) );
NOR2_Z1 g60029 ( .a(n_838), .b(n_344), .o(n_1100) );
BUF_X2 newInst_1347 ( .a(newNet_1346), .o(newNet_1347) );
INV_X1 g35129 ( .a(n_3477), .o(n_4570) );
INV_X1 g61115 ( .a(n_4625), .o(n_37) );
INV_X2 newInst_657 ( .a(newNet_656), .o(newNet_657) );
INV_X1 g60955 ( .a(n_173), .o(n_174) );
NAND4_Z2 g35187 ( .a(n_3404), .b(n_3403), .c(n_3402), .d(n_3411), .o(n_4617) );
NAND2_Z01 g59438 ( .a(n_64), .b(n_1650), .o(n_1682) );
BUF_X2 newInst_1353 ( .a(newNet_1352), .o(newNet_1353) );
BUF_X2 newInst_1506 ( .a(newNet_1505), .o(newNet_1506) );
NOR2_Z1 g34431 ( .a(n_4088), .b(n_3453), .o(n_4106) );
BUF_X2 newInst_873 ( .a(newNet_872), .o(newNet_873) );
AND2_X1 g60612 ( .a(n_359), .b(SP_3_), .o(n_592) );
NAND2_Z01 g59123 ( .a(io_do_5), .b(n_1877), .o(n_1988) );
BUF_X2 newInst_1065 ( .a(newNet_1064), .o(newNet_1065) );
BUF_X2 newInst_767 ( .a(newNet_766), .o(newNet_767) );
NAND4_Z1 g34585 ( .a(n_3750), .b(n_3752), .c(n_3753), .d(n_3749), .o(n_3975) );
NOR4_Z1 g34926 ( .a(n_3449), .b(n_3523), .c(n_4648), .d(n_3231), .o(n_3639) );
AND2_X1 g34352 ( .a(n_4180), .b(n_4534), .o(n_4230) );
NAND2_Z01 g59918 ( .a(n_1020), .b(n_375), .o(n_1195) );
INV_X1 g61028 ( .a(pY_4_), .o(n_124) );
fflopd GPR_reg_0__6_ ( .CK(newNet_1774), .D(n_3064), .Q(GPR_0__6_) );
BUF_X2 newInst_590 ( .a(newNet_502), .o(newNet_590) );
NOR2_Z1 g60416 ( .a(n_436), .b(n_4474), .o(n_730) );
NOR2_Z1 g34413 ( .a(n_4090), .b(n_3991), .o(n_4124) );
NAND2_Z01 g60038 ( .a(n_856), .b(n_4635), .o(n_1092) );
AND2_X1 g59025 ( .a(n_1983), .b(pY_8_), .o(n_2077) );
NAND2_Z01 g57723 ( .a(n_830), .b(n_3131), .o(n_3158) );
NOR2_Z1 final_adder_mux_R16_278_6_g444 ( .a(n_4450), .b(n_4434), .o(final_adder_mux_R16_278_6_n_5) );
NAND4_Z1 g34072 ( .a(n_4197), .b(n_4390), .c(n_4384), .d(n_4198), .o(dmem_do_0) );
BUF_X2 newInst_396 ( .a(newNet_395), .o(newNet_396) );
NAND2_Z01 g60041 ( .a(n_856), .b(n_4606), .o(n_1089) );
NAND2_Z01 g60911 ( .a(PC_6_), .b(pmem_d_6), .o(n_230) );
BUF_X2 newInst_1138 ( .a(newNet_1137), .o(newNet_1138) );
BUF_X2 newInst_246 ( .a(newNet_245), .o(newNet_246) );
BUF_X2 newInst_1742 ( .a(newNet_1741), .o(newNet_1742) );
NAND2_Z01 g60464 ( .a(n_341), .b(pY_0_), .o(n_682) );
BUF_X2 newInst_337 ( .a(newNet_336), .o(newNet_337) );
BUF_X2 newInst_678 ( .a(newNet_677), .o(newNet_678) );
NAND2_Z01 g34853 ( .a(n_3582), .b(GPR_0__0_), .o(n_3710) );
NAND2_Z01 g34938 ( .a(n_3542), .b(n_3307), .o(n_3637) );
NOR4_Z1 g34217 ( .a(n_4210), .b(n_4212), .c(n_4287), .d(n_4115), .o(n_4309) );
NAND2_Z01 g60192 ( .a(n_741), .b(n_642), .o(n_953) );
NAND2_Z01 g34856 ( .a(n_3581), .b(GPR_16__0_), .o(n_3707) );
XOR2_X1 g60675 ( .a(n_259), .b(n_63), .o(n_474) );
BUF_X2 newInst_474 ( .a(newNet_473), .o(newNet_474) );
NAND2_Z01 g34836 ( .a(n_3567), .b(GPR_6__1_), .o(n_3727) );
NOR2_Z1 g58449 ( .a(n_2614), .b(n_1702), .o(n_2644) );
NOR2_Z1 g59109 ( .a(n_1891), .b(n_117), .o(n_2000) );
NOR2_Z1 g35400 ( .a(n_3210), .b(n_3223), .o(n_4522) );
NAND2_Z01 g35448 ( .a(n_3247), .b(n_3220), .o(n_3270) );
NOR2_Z1 g35253 ( .a(n_3317), .b(pX_10_), .o(n_4516) );
BUF_X2 newInst_661 ( .a(newNet_77), .o(newNet_661) );
fflopd GPR_reg_8__7_ ( .CK(newNet_692), .D(n_3146), .Q(GPR_8__7_) );
BUF_X2 newInst_1592 ( .a(newNet_1255), .o(newNet_1592) );
NAND2_Z01 g34732 ( .a(n_3594), .b(GPR_6__5_), .o(n_3833) );
BUF_X2 newInst_541 ( .a(newNet_540), .o(newNet_541) );
AND2_X1 g34317 ( .a(n_4154), .b(n_4088), .o(n_4216) );
BUF_X2 newInst_869 ( .a(newNet_868), .o(newNet_869) );
INV_X1 g59500 ( .a(n_1623), .o(n_1624) );
fflopd GPR_reg_19__7_ ( .CK(newNet_1269), .D(n_3160), .Q(GPR_19__7_) );
NAND2_Z01 g34786 ( .a(n_3635), .b(GPR_14__3_), .o(n_3779) );
AND2_X1 g35058 ( .a(n_4629), .b(n_3238), .o(n_3524) );
AND2_X1 g59851 ( .a(n_1199), .b(io_do_7), .o(n_1276) );
NAND2_Z01 g60695 ( .a(GPR_1__1_), .b(n_183), .o(n_443) );
NAND2_Z01 g34735 ( .a(n_3630), .b(pX_13_), .o(n_3830) );
AND2_X1 g59155 ( .a(n_1893), .b(n_4596), .o(n_1944) );
NAND2_Z01 g35270 ( .a(pZ_13_), .b(n_3199), .o(n_3404) );
INV_X1 g60089 ( .a(n_1044), .o(n_1045) );
BUF_X2 newInst_1628 ( .a(newNet_1627), .o(newNet_1628) );
NOR2_Z1 g60768 ( .a(n_197), .b(n_160), .o(n_457) );
NAND2_Z01 g35416 ( .a(pZ_2_), .b(pmem_d_2), .o(n_3290) );
NAND2_Z01 g35432 ( .a(n_3236), .b(pmem_d_3), .o(n_4488) );
NOR2_Z1 g34419 ( .a(n_4610), .b(n_3519), .o(n_4118) );
BUF_X2 newInst_103 ( .a(newNet_9), .o(newNet_103) );
NOR3_Z1 g59251 ( .a(n_1553), .b(n_1744), .c(n_1621), .o(n_1861) );
NAND2_Z01 final_adder_mux_R16_278_6_g396 ( .a(final_adder_mux_R16_278_6_n_51), .b(final_adder_mux_R16_278_6_n_25), .o(final_adder_mux_R16_278_6_n_53) );
BUF_X2 newInst_1497 ( .a(newNet_1496), .o(newNet_1497) );
NAND4_Z1 g57914 ( .a(n_1951), .b(n_2455), .c(n_2991), .d(n_2016), .o(n_3025) );
BUF_X2 newInst_731 ( .a(newNet_730), .o(newNet_731) );
NAND2_Z01 g35366 ( .a(n_3282), .b(n_3308), .o(n_3323) );
NOR2_Z1 g59522 ( .a(n_576), .b(n_1547), .o(n_1606) );
BUF_X2 newInst_1287 ( .a(newNet_1286), .o(newNet_1287) );
XOR2_X1 g60390 ( .a(n_285), .b(n_151), .o(n_756) );
NAND2_Z01 g59103 ( .a(n_1894), .b(n_1114), .o(n_2006) );
AND2_X1 g35088 ( .a(n_3485), .b(pX_6_), .o(n_3507) );
NAND2_Z01 g34434 ( .a(n_4100), .b(n_4533), .o(n_4126) );
NAND3_Z1 g59495 ( .a(n_1542), .b(n_1417), .c(n_308), .o(n_1633) );
BUF_X2 newInst_579 ( .a(newNet_578), .o(newNet_579) );
NOR2_Z1 g34904 ( .a(n_3562), .b(n_3266), .o(n_3659) );
BUF_X2 newInst_854 ( .a(newNet_752), .o(newNet_854) );
BUF_X2 newInst_823 ( .a(newNet_822), .o(newNet_823) );
BUF_X2 newInst_498 ( .a(newNet_497), .o(newNet_498) );
BUF_X2 newInst_1594 ( .a(newNet_1593), .o(newNet_1594) );
BUF_X2 newInst_221 ( .a(newNet_220), .o(newNet_221) );
NAND2_Z01 g60735 ( .a(n_203), .b(SP_6_), .o(n_404) );
NAND2_Z01 g59069 ( .a(n_1902), .b(n_4591), .o(n_2038) );
BUF_X2 newInst_1212 ( .a(newNet_1211), .o(newNet_1212) );
BUF_X2 newInst_1577 ( .a(newNet_1576), .o(newNet_1577) );
AND2_X1 g57900 ( .a(n_3009), .b(n_2205), .o(n_3038) );
BUF_X2 newInst_13 ( .a(newNet_12), .o(newNet_13) );
NAND2_Z01 g58481 ( .a(n_834), .b(n_2588), .o(n_2621) );
NAND2_Z01 g34818 ( .a(n_3631), .b(GPR_11__2_), .o(n_3745) );
BUF_X2 newInst_1690 ( .a(newNet_1689), .o(newNet_1690) );
BUF_X2 newInst_642 ( .a(newNet_641), .o(newNet_642) );
NAND3_Z1 g59421 ( .a(n_1591), .b(n_66), .c(n_4641), .o(n_1703) );
fflopd pZ_reg_14_ ( .CK(newNet_88), .D(n_3137), .Q(pZ_14_) );
NAND2_Z01 g34388 ( .a(n_4100), .b(SP_4_), .o(n_4151) );
INV_X1 g60535 ( .a(n_594), .o(n_595) );
NAND3_Z1 g59725 ( .a(n_848), .b(n_1272), .c(n_787), .o(n_1402) );
BUF_X2 newInst_889 ( .a(newNet_224), .o(newNet_889) );
NAND2_Z01 g58717 ( .a(n_2208), .b(GPR_21__6_), .o(n_2390) );
NAND2_Z01 g60976 ( .a(n_84), .b(n_59), .o(n_192) );
NOR2_Z1 g60928 ( .a(n_45), .b(pmem_d_11), .o(n_217) );
NOR2_Z1 g59845 ( .a(n_1141), .b(n_1134), .o(n_1281) );
INV_X1 g35422 ( .a(n_3289), .o(n_3288) );
NAND2_Z01 g34715 ( .a(n_3594), .b(GPR_7__6_), .o(n_3850) );
BUF_X2 newInst_413 ( .a(newNet_412), .o(newNet_413) );
NAND2_Z01 g60923 ( .a(PC_3_), .b(pmem_d_3), .o(n_220) );
NAND2_Z01 g34889 ( .a(n_3630), .b(pX_8_), .o(n_3674) );
BUF_X2 newInst_283 ( .a(newNet_282), .o(newNet_283) );
NAND2_Z01 g60414 ( .a(n_360), .b(GPR_3__4_), .o(n_732) );
NOR2_Z1 g34546 ( .a(n_3918), .b(n_3346), .o(n_4012) );
NAND2_Z01 g59644 ( .a(io_do_4), .b(n_1418), .o(n_1477) );
BUF_X2 newInst_1395 ( .a(newNet_1394), .o(newNet_1395) );
BUF_X2 newInst_1003 ( .a(newNet_104), .o(newNet_1003) );
BUF_X2 newInst_1437 ( .a(newNet_1436), .o(newNet_1437) );
NAND2_Z01 g34527 ( .a(n_3756), .b(n_3942), .o(n_4017) );
AND2_X1 g58649 ( .a(n_2362), .b(n_1620), .o(n_2452) );
AND2_X1 g57890 ( .a(n_3009), .b(n_2156), .o(n_3048) );
INV_X1 g35128 ( .a(n_3478), .o(n_4628) );
NAND2_Z01 g60721 ( .a(n_198), .b(GPR_23__2_), .o(n_417) );
NOR2_Z1 g34181 ( .a(n_4324), .b(n_4615), .o(n_4420) );
NAND2_Z01 g34899 ( .a(n_3577), .b(pY_6_), .o(n_3664) );
INV_X1 g34974 ( .a(n_3596), .o(n_3597) );
NAND4_Z1 g60137 ( .a(n_658), .b(n_646), .c(n_625), .d(n_738), .o(n_995) );
NOR2_Z1 g59653 ( .a(n_1403), .b(n_950), .o(n_1472) );
NAND2_Z01 g60293 ( .a(n_596), .b(GPR_3__5_), .o(n_831) );
NAND2_Z01 g58840 ( .a(n_2159), .b(GPR_10__6_), .o(n_2267) );
NOR3_Z1 g58946 ( .a(n_67), .b(n_1943), .c(n_70), .o(n_2151) );
BUF_X2 newInst_1767 ( .a(newNet_1766), .o(newNet_1767) );
BUF_X2 newInst_1405 ( .a(newNet_1404), .o(newNet_1405) );
NAND2_Z01 g35407 ( .a(pY_1_), .b(pmem_d_1), .o(n_3296) );
BUF_X2 newInst_480 ( .a(newNet_258), .o(newNet_480) );
NOR2_Z1 g59878 ( .a(n_1155), .b(n_1166), .o(n_1249) );
NAND2_Z01 g58316 ( .a(n_2679), .b(n_2370), .o(n_2749) );
NAND2_Z01 g58816 ( .a(n_2176), .b(io_do_7), .o(n_2285) );
INV_X1 g35470 ( .a(pmem_d_10), .o(n_3254) );
NAND2_Z01 g35430 ( .a(n_3236), .b(pmem_d_12), .o(n_4482) );
NAND2_Z01 g60434 ( .a(n_342), .b(GPR_17__6_), .o(n_712) );
AND2_X1 g59572 ( .a(n_1468), .b(pmem_d_1), .o(n_1556) );
NAND2_Z01 g34760 ( .a(n_3635), .b(GPR_14__4_), .o(n_3805) );
BUF_X2 newInst_1673 ( .a(newNet_1672), .o(newNet_1673) );
NAND2_Z01 g34400 ( .a(n_3208), .b(pZ_4_), .o(n_4138) );
NAND2_Z01 g34397 ( .a(n_3208), .b(pZ_7_), .o(n_4141) );
INV_X1 g34559 ( .a(n_3985), .o(n_4000) );
BUF_X2 newInst_1297 ( .a(newNet_1296), .o(newNet_1297) );
fflopd GPR_reg_7__7_ ( .CK(newNet_739), .D(n_3147), .Q(GPR_7__7_) );
BUF_X2 newInst_1478 ( .a(newNet_1477), .o(newNet_1478) );
AND4_X1 g34066 ( .a(n_4142), .b(n_4232), .c(n_4395), .d(n_4128), .o(dmem_a_9) );
BUF_X2 newInst_599 ( .a(newNet_598), .o(newNet_599) );
AND2_X1 g34919 ( .a(n_3593), .b(pY_10_), .o(n_3644) );
XNOR2_X1 g35018 ( .a(n_3527), .b(PC_8_), .o(n_4539) );
NAND2_Z01 g60918 ( .a(n_95), .b(pX_6_), .o(n_224) );
BUF_X2 newInst_24 ( .a(newNet_23), .o(newNet_24) );
NOR2_Z1 g34990 ( .a(n_3535), .b(n_3482), .o(n_3592) );
BUF_X1 mybuffer1 ( .o(io_a_1), .a(pmem_d_1) );
NAND2_Z01 g59124 ( .a(n_1896), .b(n_1287), .o(n_1987) );
NAND2_Z01 g60550 ( .a(n_360), .b(GPR_1__2_), .o(n_556) );
XOR2_X1 g59032 ( .a(io_do_5), .b(n_1877), .o(n_2087) );
AND2_X1 g60985 ( .a(PC_4_), .b(pmem_d_7), .o(n_185) );
NAND2_Z01 g58767 ( .a(n_2202), .b(GPR_5__3_), .o(n_2333) );
fflopd GPR_reg_14__6_ ( .CK(newNet_1537), .D(n_3086), .Q(GPR_14__6_) );
NAND2_Z01 g34096 ( .a(n_4371), .b(n_4370), .o(n_4438) );
BUF_X2 newInst_1398 ( .a(newNet_1397), .o(newNet_1398) );
BUF_X2 newInst_449 ( .a(newNet_448), .o(newNet_449) );
NAND2_Z01 g35358 ( .a(n_3200), .b(n_3233), .o(n_4660) );
AND2_X1 g35290 ( .a(n_3260), .b(n_3298), .o(n_3385) );
NAND2_Z01 g60403 ( .a(n_372), .b(U_14_), .o(n_743) );
INV_X2 newInst_1174 ( .a(newNet_1173), .o(newNet_1174) );
NOR2_Z1 g60808 ( .a(n_182), .b(n_258), .o(n_361) );
INV_X1 g35065 ( .a(n_3521), .o(n_4591) );
BUF_X2 newInst_1312 ( .a(newNet_1311), .o(newNet_1312) );
NAND2_Z01 g35083 ( .a(n_3491), .b(n_3469), .o(n_3511) );
NOR2_Z1 g34997 ( .a(n_3550), .b(n_3484), .o(n_3585) );
INV_X1 g60285 ( .a(n_844), .o(n_843) );
AND3_X1 g60666 ( .a(n_4631), .b(n_346), .c(n_4483), .o(n_480) );
NAND4_Z1 g59044 ( .a(n_1507), .b(n_1675), .c(n_1886), .d(n_1506), .o(n_2065) );
fflopd GPR_reg_11__5_ ( .CK(newNet_1688), .D(n_3020), .Q(GPR_11__5_) );
BUF_X2 newInst_1302 ( .a(newNet_1301), .o(newNet_1302) );
AND2_X1 g59472 ( .a(n_1600), .b(n_850), .o(n_1652) );
AND3_X1 g59194 ( .a(n_1112), .b(n_1895), .c(pZ_6_), .o(n_1915) );
BUF_X2 newInst_1052 ( .a(newNet_1051), .o(newNet_1052) );
BUF_X2 newInst_1008 ( .a(newNet_1007), .o(newNet_1008) );
NAND3_Z1 g34085 ( .a(n_4377), .b(n_4322), .c(n_4219), .o(dmem_do_4) );
NAND2_Z01 g60493 ( .a(n_347), .b(GPR_9__3_), .o(n_653) );
NAND2_Z01 g60050 ( .a(n_867), .b(pY_5_), .o(n_1114) );
INV_X1 g34631 ( .a(n_4587), .o(n_3929) );
BUF_X2 newInst_96 ( .a(newNet_95), .o(newNet_96) );
NAND2_Z01 g57713 ( .a(n_3127), .b(n_2381), .o(n_3154) );
BUF_X2 newInst_1549 ( .a(newNet_1548), .o(newNet_1549) );
NAND2_Z01 g60427 ( .a(n_357), .b(pY_10_), .o(n_719) );
AND2_X1 g58513 ( .a(n_2567), .b(n_2203), .o(n_2583) );
AND2_X1 g58503 ( .a(n_2567), .b(n_2213), .o(n_2594) );
BUF_X2 newInst_132 ( .a(newNet_131), .o(newNet_132) );
NAND2_Z01 g60899 ( .a(C), .b(pmem_d_0), .o(n_271) );
BUF_X2 newInst_1163 ( .a(newNet_1162), .o(newNet_1163) );
INV_X1 g61077 ( .a(GPR_14__6_), .o(n_75) );
NAND4_Z1 g57731 ( .a(n_2079), .b(n_2540), .c(n_3103), .d(n_1971), .o(n_3141) );
NAND2_Z01 g60186 ( .a(n_664), .b(n_711), .o(n_968) );
NAND2_Z01 g59606 ( .a(n_1415), .b(N), .o(n_1520) );
NAND2_Z01 g60690 ( .a(GPR_0__1_), .b(n_183), .o(n_448) );
NAND2_Z01 g60326 ( .a(n_519), .b(n_464), .o(n_863) );
BUF_X2 newInst_1759 ( .a(newNet_1758), .o(newNet_1759) );
NAND2_Z01 g60460 ( .a(n_371), .b(GPR_21__0_), .o(n_686) );
NAND2_Z01 g59641 ( .a(io_do_1), .b(n_1418), .o(n_1480) );
BUF_X2 newInst_1011 ( .a(newNet_1010), .o(newNet_1011) );
BUF_X2 newInst_880 ( .a(newNet_879), .o(newNet_880) );
NAND2_Z01 g60102 ( .a(n_867), .b(n_103), .o(n_1018) );
NAND2_Z01 g60206 ( .a(n_582), .b(GPR_11__3_), .o(n_939) );
AND2_X1 g59873 ( .a(n_1168), .b(n_286), .o(n_1254) );
AND2_X1 g59372 ( .a(n_1679), .b(n_1136), .o(n_1766) );
BUF_X2 newInst_1828 ( .a(newNet_321), .o(newNet_1828) );
INV_X1 g35233 ( .a(n_4572), .o(n_3421) );
INV_X1 g61040 ( .a(pY_13_), .o(n_112) );
fflopd GPR_reg_22__4_ ( .CK(newNet_1085), .D(n_2932), .Q(GPR_22__4_) );
BUF_X2 newInst_25 ( .a(newNet_24), .o(newNet_25) );
AND2_X1 g58401 ( .a(n_2657), .b(n_2153), .o(n_2667) );
BUF_X2 newInst_444 ( .a(newNet_443), .o(newNet_444) );
NOR2_Z1 g34360 ( .a(n_4126), .b(n_3250), .o(n_4179) );
NAND2_Z01 g58145 ( .a(n_2821), .b(n_2297), .o(n_2868) );
NAND2_Z01 g58460 ( .a(n_2598), .b(n_2254), .o(n_2636) );
NAND2_Z01 g60578 ( .a(io_do_1), .b(n_377), .o(n_533) );
AND2_X1 g58273 ( .a(n_2752), .b(n_2199), .o(n_2794) );
NAND2_Z01 g34626 ( .a(n_3644), .b(pY_11_), .o(n_3934) );
NAND2_Z01 g58174 ( .a(n_2834), .b(n_928), .o(n_2851) );
NAND2_Z01 g34742 ( .a(n_3585), .b(GPR_13__5_), .o(n_3823) );
NAND2_Z01 g34083 ( .a(n_4164), .b(GPR_Rd_r_0_), .o(n_4390) );
XOR2_X1 g34927 ( .a(n_3546), .b(pZ_9_), .o(n_3767) );
NOR2_Z1 g34335 ( .a(n_16064_BAR), .b(n_3420), .o(n_4199) );
NAND4_Z1 g34590 ( .a(n_3726), .b(n_3727), .c(n_3729), .d(n_3728), .o(n_3970) );
BUF_X2 newInst_1693 ( .a(newNet_1692), .o(newNet_1693) );
BUF_X2 newInst_1183 ( .a(newNet_1182), .o(newNet_1183) );
NOR2_Z1 g34999 ( .a(n_3553), .b(n_3490), .o(n_3582) );
NOR2_Z1 g59332 ( .a(n_1704), .b(n_1386), .o(n_1805) );
NAND2_Z01 g60318 ( .a(n_600), .b(pX_6_), .o(n_808) );
BUF_X2 newInst_1135 ( .a(newNet_1134), .o(newNet_1135) );
BUF_X2 newInst_371 ( .a(newNet_370), .o(newNet_371) );
NAND2_Z01 g58308 ( .a(n_2685), .b(n_2394), .o(n_2762) );
NAND2_Z01 g34337 ( .a(n_4166), .b(n_4555), .o(n_4197) );
BUF_X2 newInst_1807 ( .a(newNet_1806), .o(newNet_1807) );
BUF_X2 newInst_1083 ( .a(newNet_1082), .o(newNet_1083) );
NAND2_Z01 g58736 ( .a(n_2205), .b(GPR_2__1_), .o(n_2371) );
BUF_X2 newInst_782 ( .a(newNet_781), .o(newNet_782) );
NAND4_Z1 g58134 ( .a(n_2071), .b(n_2546), .c(n_2826), .d(n_2053), .o(n_2879) );
AND2_X1 g60600 ( .a(n_460), .b(n_250), .o(n_599) );
NAND2_Z01 g35395 ( .a(pmem_d_15), .b(pmem_d_2), .o(n_4636) );
XOR2_X1 g34930 ( .a(n_3538), .b(n_3226), .o(n_4598) );
NAND2_Z01 g59313 ( .a(n_1726), .b(n_264), .o(n_1807) );
NAND2_Z01 g59461 ( .a(n_1596), .b(SP_6_), .o(n_1660) );
AND2_X1 g34421 ( .a(n_4088), .b(n_4030), .o(n_4116) );
NOR2_Z4 g58177 ( .a(n_2791), .b(n_1587), .o(n_2850) );
BUF_X2 newInst_1850 ( .a(newNet_1214), .o(newNet_1850) );
BUF_X2 newInst_193 ( .a(newNet_192), .o(newNet_193) );
BUF_X2 newInst_238 ( .a(newNet_237), .o(newNet_238) );
NAND2_Z01 g35004 ( .a(n_3509), .b(n_3549), .o(n_3574) );
NAND2_X2 g58906 ( .a(n_2141), .b(n_2090), .o(n_2216) );
BUF_X2 newInst_311 ( .a(newNet_310), .o(newNet_311) );
NAND4_Z1 g58983 ( .a(io_do_0), .b(n_1420), .c(n_1861), .d(n_41), .o(n_2124) );
fflopd pY_reg_6_ ( .CK(newNet_137), .D(n_3113), .Q(pY_6_) );
XOR2_X1 g59413 ( .a(n_1489), .b(n_1602), .o(n_1730) );
BUF_X2 newInst_1761 ( .a(newNet_1760), .o(newNet_1761) );
NOR2_Z1 g34424 ( .a(n_4097), .b(n_3973), .o(n_4113) );
INV_Z1 g16799 ( .a(n_4643), .o(n_4418) );
NAND2_Z01 g58103 ( .a(n_2836), .b(n_495), .o(n_2910) );
NAND2_Z01 g60237 ( .a(n_574), .b(GPR_10__6_), .o(n_908) );
NAND2_Z01 g57947 ( .a(n_2960), .b(n_2305), .o(n_2995) );
fflopd GPR_reg_2__3_ ( .CK(newNet_1002), .D(n_2846), .Q(GPR_2__3_) );
NAND2_Z01 g59134 ( .a(n_1872), .b(n_1052), .o(n_1964) );
BUF_X2 newInst_172 ( .a(newNet_82), .o(newNet_172) );
INV_X1 g61116 ( .a(pmem_d_10), .o(n_36) );
NAND4_Z1 g34227 ( .a(n_4110), .b(n_4200), .c(n_4242), .d(n_4137), .o(n_4304) );
AND2_X1 g57909 ( .a(n_3009), .b(n_2199), .o(n_3030) );
NAND2_Z01 g57705 ( .a(n_3136), .b(n_2186), .o(n_3164) );
BUF_X2 newInst_626 ( .a(newNet_625), .o(newNet_626) );
AND2_X1 g59849 ( .a(n_1158), .b(rst), .o(n_1277) );
NAND3_Z1 g59185 ( .a(n_1815), .b(n_1865), .c(n_795), .o(n_1922) );
NAND2_Z01 g35344 ( .a(n_4486), .b(pmem_d_12), .o(n_4683) );
AND2_X1 g58365 ( .a(n_2656), .b(n_2214), .o(n_2706) );
NAND2_Z01 g58775 ( .a(n_2201), .b(GPR_6__3_), .o(n_2325) );
NAND2_Z01 g59362 ( .a(n_852), .b(n_15), .o(n_1751) );
BUF_X2 newInst_1319 ( .a(newNet_1318), .o(newNet_1319) );
NAND4_Z1 g57773 ( .a(n_1680), .b(n_1524), .c(n_3063), .d(n_1081), .o(n_3108) );
BUF_X2 newInst_1603 ( .a(newNet_1602), .o(newNet_1603) );
BUF_X2 newInst_290 ( .a(newNet_289), .o(newNet_290) );
XOR2_X1 g59379 ( .a(n_1662), .b(SP_14_), .o(n_1739) );
NAND2_Z01 g58728 ( .a(n_2206), .b(GPR_23__1_), .o(n_2379) );
XOR2_X1 g59813 ( .a(n_1186), .b(n_54), .o(n_1316) );
XOR2_X1 g59598 ( .a(n_1453), .b(PC_5_), .o(n_1531) );
NAND2_Z01 g59832 ( .a(n_1206), .b(io_do_3), .o(n_1293) );
BUF_X2 newInst_1281 ( .a(newNet_1280), .o(newNet_1281) );
NAND2_Z01 g57949 ( .a(n_2985), .b(n_836), .o(n_3010) );
BUF_X2 newInst_330 ( .a(newNet_329), .o(newNet_330) );
NAND2_Z01 g60397 ( .a(n_417), .b(n_455), .o(n_749) );
NAND2_Z01 g34538 ( .a(n_3915), .b(n_3926), .o(pmem_a_8) );
NAND4_Z1 g58014 ( .a(n_1918), .b(n_2508), .c(n_2916), .d(n_2055), .o(n_2958) );
NOR2_Z1 g34292 ( .a(n_4163), .b(n_3236), .o(n_4241) );
BUF_X2 newInst_212 ( .a(newNet_211), .o(newNet_212) );
AND3_X1 g59994 ( .a(n_111), .b(n_1112), .c(pZ_7_), .o(n_1135) );
BUF_X2 newInst_351 ( .a(newNet_350), .o(newNet_351) );
BUF_X2 newInst_1370 ( .a(newNet_1369), .o(newNet_1370) );
INV_X1 g60012 ( .a(n_1116), .o(n_1117) );
NAND2_Z01 g60301 ( .a(n_586), .b(n_274), .o(n_823) );
fflopd GPR_reg_17__0_ ( .CK(newNet_1417), .D(n_2639), .Q(GPR_17__0_) );
BUF_X2 newInst_832 ( .a(newNet_831), .o(newNet_832) );
NAND2_Z01 g60890 ( .a(n_4486), .b(n_32), .o(n_276) );
AND2_X1 g58498 ( .a(n_2567), .b(n_2158), .o(n_2599) );
BUF_X2 newInst_957 ( .a(newNet_956), .o(newNet_957) );
INV_X1 g34558 ( .a(n_3998), .o(n_4001) );
BUF_X2 newInst_726 ( .a(newNet_493), .o(newNet_726) );
NAND2_Z01 g34118 ( .a(io_do_1), .b(n_4177), .o(n_4385) );
NAND2_Z01 g35391 ( .a(SP_8_), .b(SP_9_), .o(n_4534) );
NAND4_Z1 g34063 ( .a(n_4279), .b(n_4243), .c(n_4398), .d(n_4144), .o(dmem_a_11) );
NAND2_Z01 g58712 ( .a(n_2208), .b(GPR_21__1_), .o(n_2395) );
AND2_X1 g59171 ( .a(n_1895), .b(pZ_14_), .o(n_1976) );
AND2_X1 g34513 ( .a(n_3984), .b(n_3983), .o(n_4032) );
BUF_X2 newInst_904 ( .a(newNet_903), .o(newNet_904) );
BUF_X2 newInst_184 ( .a(newNet_183), .o(newNet_184) );
NAND3_Z1 g59302 ( .a(n_1681), .b(n_1652), .c(n_798), .o(n_1812) );
NOR2_Z1 g60986 ( .a(PC_1_), .b(pmem_d_1), .o(n_144) );
BUF_X2 newInst_1638 ( .a(newNet_1637), .o(newNet_1638) );
NAND3_Z1 g59247 ( .a(n_24), .b(n_1773), .c(n_41), .o(n_1869) );
AND2_X1 g57752 ( .a(n_3115), .b(n_2153), .o(n_3119) );
BUF_X2 newInst_1075 ( .a(newNet_50), .o(newNet_1075) );
NAND2_Z01 g34669 ( .a(n_3609), .b(n_3610), .o(n_3896) );
NAND2_Z01 g58155 ( .a(n_2810), .b(n_2365), .o(n_2858) );
NOR2_Z1 g34903 ( .a(n_3578), .b(n_3210), .o(n_3660) );
NAND2_Z02 g58962 ( .a(n_2115), .b(n_1215), .o(n_2155) );
BUF_X2 newInst_1725 ( .a(newNet_1724), .o(newNet_1725) );
NAND2_Z01 g60304 ( .a(n_617), .b(n_129), .o(n_820) );
BUF_X2 newInst_1720 ( .a(newNet_1719), .o(newNet_1720) );
AND2_X1 g59230 ( .a(n_1833), .b(n_1036), .o(n_1882) );
NAND2_Z01 g60522 ( .a(n_374), .b(GPR_12__2_), .o(n_624) );
NAND2_Z02 g58974 ( .a(n_2088), .b(n_1209), .o(n_2139) );
BUF_X2 newInst_851 ( .a(newNet_850), .o(newNet_851) );
NAND2_Z01 g59326 ( .a(n_4), .b(n_4539), .o(n_1787) );
INV_X1 g34801 ( .a(n_4585), .o(n_3762) );
NOR2_Z1 g34358 ( .a(n_4148), .b(n_3648), .o(n_4173) );
NAND3_Z1 g35188 ( .a(n_3383), .b(n_3441), .c(n_3407), .o(n_4619) );
XNOR2_X1 g60851 ( .a(n_4444), .b(n_4428), .o(n_290) );
INV_X1 g35323 ( .a(n_3347), .o(n_3346) );
BUF_X2 newInst_1588 ( .a(newNet_1587), .o(newNet_1588) );
AND2_X1 g57745 ( .a(n_3115), .b(n_2206), .o(n_3126) );
BUF_X2 newInst_1227 ( .a(newNet_1226), .o(newNet_1227) );
BUF_X2 newInst_943 ( .a(newNet_942), .o(newNet_943) );
NAND2_Z01 g34956 ( .a(n_3552), .b(GPR_3__1_), .o(n_3606) );
NAND2_Z01 g58675 ( .a(n_2214), .b(GPR_16__0_), .o(n_2431) );
NAND2_Z01 final_adder_mux_R16_278_6_g378 ( .a(final_adder_mux_R16_278_6_n_69), .b(final_adder_mux_R16_278_6_n_21), .o(final_adder_mux_R16_278_6_n_71) );
BUF_X2 newInst_1153 ( .a(newNet_1152), .o(newNet_1153) );
BUF_X2 newInst_713 ( .a(newNet_712), .o(newNet_713) );
NAND2_Z01 g60554 ( .a(n_404), .b(n_394), .o(n_552) );
NAND2_Z01 g34108 ( .a(n_4338), .b(n_4353), .o(n_4448) );
NAND2_Z01 g60076 ( .a(io_do_7), .b(n_841), .o(n_1059) );
BUF_X2 newInst_1684 ( .a(newNet_1041), .o(newNet_1684) );
INV_X1 g61073 ( .a(GPR_14__2_), .o(n_79) );
NAND2_Z01 g58591 ( .a(n_2461), .b(pX_4_), .o(n_2507) );
NAND2_Z01 g57836 ( .a(n_3040), .b(n_2382), .o(n_3074) );
AND2_X1 g58927 ( .a(n_2138), .b(pmem_d_11), .o(n_2176) );
NOR2_Z1 g59013 ( .a(n_1980), .b(n_101), .o(n_2095) );
INV_X1 g61036 ( .a(state_0_), .o(n_116) );
INV_X1 g61103 ( .a(n_4526), .o(n_49) );
NAND2_Z01 g59516 ( .a(n_1549), .b(n_65), .o(n_1623) );
INV_X1 g58659 ( .a(n_2442), .o(n_2443) );
BUF_X2 newInst_1615 ( .a(newNet_1614), .o(newNet_1615) );
BUF_X2 newInst_120 ( .a(newNet_119), .o(newNet_120) );
fflopd GPR_reg_9__2_ ( .CK(newNet_681), .D(n_2736), .Q(GPR_9__2_) );
BUF_X2 newInst_1027 ( .a(newNet_1026), .o(newNet_1027) );
XOR2_X1 g60391 ( .a(n_283), .b(n_143), .o(n_755) );
NOR2_Z1 g60837 ( .a(n_4482), .b(n_252), .o(n_296) );
AND2_X1 g34365 ( .a(n_4124), .b(Rd_0_), .o(n_4170) );
NAND2_Z01 g34614 ( .a(n_3898), .b(n_3491), .o(n_3946) );
NOR2_Z1 g60819 ( .a(n_4561), .b(n_175), .o(n_307) );
NOR4_Z1 g57952 ( .a(n_2558), .b(n_2837), .c(n_2920), .d(n_1407), .o(n_2993) );
NAND2_Z02 g58914 ( .a(n_2160), .b(n_1204), .o(n_2208) );
NAND2_Z01 g59322 ( .a(n_4), .b(n_4547), .o(n_1791) );
NAND4_Z1 g60142 ( .a(n_718), .b(n_687), .c(n_721), .d(n_719), .o(n_990) );
NAND2_Z01 g60332 ( .a(n_577), .b(pmem_d_10), .o(n_862) );
NAND4_Z1 g58487 ( .a(n_1521), .b(n_2445), .c(n_2555), .d(n_1235), .o(n_2609) );
NOR3_Z1 g60122 ( .a(n_199), .b(n_511), .c(n_42), .o(n_1005) );
NAND2_Z01 g58457 ( .a(n_2432), .b(n_2594), .o(n_2639) );
BUF_X2 newInst_1444 ( .a(newNet_1443), .o(newNet_1444) );
BUF_X2 newInst_872 ( .a(newNet_553), .o(newNet_872) );
NAND2_Z01 g34666 ( .a(n_3615), .b(n_3616), .o(n_3899) );
XOR2_X1 g59369 ( .a(io_do_7), .b(n_1661), .o(n_1769) );
NAND2_Z03 g34223 ( .a(n_4291), .b(n_4000), .o(io_do_4) );
NOR3_Z1 g59199 ( .a(n_1768), .b(n_1853), .c(n_579), .o(n_1911) );
NAND2_Z02 g60623 ( .a(n_66), .b(n_366), .o(n_587) );
fflopd GPR_reg_9__3_ ( .CK(newNet_678), .D(n_2839), .Q(GPR_9__3_) );
NOR2_Z1 g58977 ( .a(n_1036), .b(n_2087), .o(n_2130) );
NAND2_Z01 g34277 ( .a(n_4160), .b(n_4586), .o(n_4256) );
NAND2_Z01 g59507 ( .a(n_1574), .b(n_133), .o(n_1628) );
INV_X1 g35518 ( .a(pY_7_), .o(n_3210) );
INV_X1 g61059 ( .a(SP_14_), .o(n_93) );
NAND4_Z1 g34562 ( .a(n_3886), .b(n_3885), .c(n_3887), .d(n_3883), .o(n_3998) );
NAND2_Z01 g59296 ( .a(n_852), .b(n_1764), .o(n_1815) );
INV_X1 g60874 ( .a(n_252), .o(n_251) );
NOR2_Z1 g59165 ( .a(n_1701), .b(n_1855), .o(n_1937) );
NAND2_Z01 g34724 ( .a(n_3597), .b(GPR_16__5_), .o(n_3841) );
INV_X1 g35067 ( .a(n_3519), .o(n_4604) );
BUF_X2 newInst_816 ( .a(newNet_815), .o(newNet_816) );
BUF_X2 newInst_582 ( .a(newNet_581), .o(newNet_582) );
NAND2_Z01 final_adder_mux_R16_278_6_g363 ( .a(final_adder_mux_R16_278_6_n_84), .b(final_adder_mux_R16_278_6_n_23), .o(final_adder_mux_R16_278_6_n_86) );
NAND2_Z01 g58801 ( .a(n_2195), .b(U_14_), .o(n_2299) );
NAND2_Z01 g58287 ( .a(n_2710), .b(n_2259), .o(n_2783) );
fflopd GPR_reg_9__0_ ( .CK(newNet_688), .D(n_2615), .Q(GPR_9__0_) );
AND2_X1 g35299 ( .a(n_3224), .b(n_3298), .o(n_3376) );
NAND2_Z01 g58713 ( .a(n_2208), .b(GPR_21__2_), .o(n_2394) );
BUF_X2 newInst_1036 ( .a(newNet_618), .o(newNet_1036) );
NOR2_Z1 g34969 ( .a(n_3553), .b(n_3482), .o(n_3629) );
BUF_X2 newInst_1642 ( .a(newNet_1641), .o(newNet_1642) );
NAND2_Z01 g34745 ( .a(n_3590), .b(pY_13_), .o(n_3820) );
AND2_X1 g59976 ( .a(n_350), .b(n_1031), .o(n_1149) );
BUF_X2 newInst_632 ( .a(newNet_631), .o(newNet_632) );
AND2_X1 g60965 ( .a(n_4630), .b(n_59), .o(n_155) );
NAND2_Z01 g34718 ( .a(n_3590), .b(pY_14_), .o(n_3847) );
BUF_X2 newInst_309 ( .a(newNet_32), .o(newNet_309) );
NAND2_Z01 g34103 ( .a(n_4356), .b(n_4350), .o(n_4450) );
AND2_X1 g58378 ( .a(n_2656), .b(n_2210), .o(n_2693) );
BUF_X2 newInst_572 ( .a(newNet_571), .o(newNet_572) );
fflopd GPR_reg_11__6_ ( .CK(newNet_1683), .D(n_3089), .Q(GPR_11__6_) );
AND2_X1 g35227 ( .a(n_3355), .b(pZ_3_), .o(n_3442) );
NOR2_Z4 g58065 ( .a(n_2883), .b(n_1583), .o(n_2940) );
BUF_X2 newInst_228 ( .a(newNet_227), .o(newNet_228) );
XOR2_X1 g60866 ( .a(n_4437), .b(n_4421), .o(n_282) );
BUF_X2 newInst_293 ( .a(newNet_292), .o(newNet_293) );
NAND2_Z01 g34894 ( .a(n_3577), .b(pY_3_), .o(n_3669) );
NAND2_Z01 g58326 ( .a(n_2668), .b(n_2318), .o(n_2739) );
BUF_X2 newInst_973 ( .a(newNet_972), .o(newNet_973) );
fflopd PC_reg_10_ ( .CK(newNet_651), .D(n_2610), .Q(PC_10_) );
BUF_X2 newInst_538 ( .a(newNet_537), .o(newNet_538) );
INV_X1 g34373 ( .a(n_4159), .o(n_4158) );
fflopd GPR_Rd_r_reg_7_ ( .CK(newNet_1835), .D(io_do_7), .Q(GPR_Rd_r_7_) );
BUF_X2 newInst_391 ( .a(newNet_390), .o(newNet_391) );
AND2_X1 g58375 ( .a(n_2656), .b(n_2211), .o(n_2696) );
BUF_X2 newInst_191 ( .a(newNet_190), .o(newNet_191) );
BUF_X2 newInst_1623 ( .a(newNet_1622), .o(newNet_1623) );
NAND2_Z01 g58724 ( .a(n_2207), .b(GPR_22__5_), .o(n_2383) );
NAND2_Z01 g59116 ( .a(n_1856), .b(io_do_3), .o(n_1993) );
BUF_X2 newInst_253 ( .a(newNet_252), .o(newNet_253) );
NOR2_Z1 g35013 ( .a(n_3511), .b(n_3535), .o(n_3563) );
NOR2_Z2 g59215 ( .a(n_1829), .b(n_16064_BAR), .o(n_1902) );
BUF_X2 newInst_1703 ( .a(newNet_1124), .o(newNet_1703) );
INV_X1 g35228 ( .a(n_3431), .o(n_3432) );
BUF_X2 newInst_1652 ( .a(newNet_1651), .o(newNet_1652) );
NAND3_Z1 g34450 ( .a(n_3838), .b(n_4051), .c(n_3839), .o(n_4090) );
NAND4_Z1 g59732 ( .a(n_945), .b(n_869), .c(n_1281), .d(n_942), .o(n_1398) );
BUF_X2 newInst_1656 ( .a(newNet_1655), .o(newNet_1656) );
BUF_X2 newInst_1240 ( .a(newNet_1239), .o(newNet_1240) );
NAND2_Z01 g60725 ( .a(n_200), .b(GPR_8__4_), .o(n_413) );
NAND2_Z01 g59180 ( .a(n_1872), .b(n_1670), .o(n_1927) );
NAND2_Z01 g59858 ( .a(n_1163), .b(n_101), .o(n_1306) );
BUF_X2 newInst_1293 ( .a(newNet_1292), .o(newNet_1293) );
NOR2_Z1 g59964 ( .a(n_1044), .b(n_969), .o(n_1172) );
BUF_X2 newInst_1648 ( .a(newNet_1647), .o(newNet_1648) );
AND2_X1 g58408 ( .a(n_2655), .b(n_1733), .o(n_2660) );
NAND4_Z1 g59889 ( .a(n_483), .b(n_898), .c(n_975), .d(n_356), .o(n_1238) );
NAND2_Z01 g60027 ( .a(n_4603), .b(n_856), .o(n_1102) );
BUF_X2 newInst_230 ( .a(newNet_229), .o(newNet_230) );
NAND2_Z01 g34912 ( .a(n_3563), .b(pZ_2_), .o(n_3651) );
NAND2_Z01 g34100 ( .a(n_4363), .b(n_4362), .o(n_4442) );
XOR2_X1 g58533 ( .a(n_2550), .b(n_2087), .o(n_2564) );
AND2_X1 g58004 ( .a(n_2940), .b(n_2204), .o(n_2967) );
AND2_X1 g57737 ( .a(n_3115), .b(n_2214), .o(n_3135) );
NAND2_Z01 g34948 ( .a(n_3552), .b(GPR_10__5_), .o(n_3614) );
NAND2_Z01 g58097 ( .a(n_2851), .b(n_2194), .o(n_2916) );

endmodule
