module INV_X1 ();
  output o;
  input a;
endmodule

module INV_X2 ();
  output o;
  input a;
endmodule

module INV_X3 ();
  output o;
  input a;
endmodule

module INV_X4 ();
  output o;
  input a;
endmodule

module INV_X6 ();
  output o;
  input a;
endmodule

module INV_X8 ();
  output o;
  input a;
endmodule

module INV_X10 ();
  output o;
  input a;
endmodule

module INV_X20 ();
  output o;
  input a;
endmodule

module INV_X40 ();
  output o;
  input a;
endmodule

module INV_X80 ();
  output o;
  input a;
endmodule

module INV_Y1 ();
  output o;
  input a;
endmodule

module INV_Y2 ();
  output o;
  input a;
endmodule

module INV_Y3 ();
  output o;
  input a;
endmodule

module INV_Y4 ();
  output o;
  input a;
endmodule

module INV_Y6 ();
  output o;
  input a;
endmodule

module INV_Y8 ();
  output o;
  input a;
endmodule

module INV_Y10 ();
  output o;
  input a;
endmodule

module INV_Y20 ();
  output o;
  input a;
endmodule

module INV_Y40 ();
  output o;
  input a;
endmodule

module INV_Y80 ();
  output o;
  input a;
endmodule

module INV_Z1 ();
  output o;
  input a;
endmodule

module INV_Z2 ();
  output o;
  input a;
endmodule

module INV_Z3 ();
  output o;
  input a;
endmodule

module INV_Z4 ();
  output o;
  input a;
endmodule

module INV_Z6 ();
  output o;
  input a;
endmodule

module INV_Z8 ();
  output o;
  input a;
endmodule

module INV_Z10 ();
  output o;
  input a;
endmodule

module INV_Z20 ();
  output o;
  input a;
endmodule

module INV_Z40 ();
  output o;
  input a;
endmodule

module INV_Z80 ();
  output o;
  input a;
endmodule

module NAND2_X1 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X2 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X3 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X4 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X6 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X8 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X10 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X20 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X40 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_X80 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y01 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y02 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y03 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y04 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y06 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y08 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y10 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y20 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y40 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Y80 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z01 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z02 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z03 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z04 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z06 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z08 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z10 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z20 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z40 ();
  output o;
  input a;
  input b;
endmodule

module NAND2_Z80 ();
  output o;
  input a;
  input b;
endmodule

module NAND3_X1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X2 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X3 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X4 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X6 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X8 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_X80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y2 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y3 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y4 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y6 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y8 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Y80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z2 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z3 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z4 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z6 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z8 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND3_Z80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NAND4_X1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X2 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X3 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X4 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X6 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X8 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_X80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y2 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y3 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y4 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y6 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y8 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Y80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z2 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z3 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z4 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z6 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z8 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NAND4_Z80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR2_X1 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X2 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X3 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X4 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X6 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X8 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X10 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X20 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X40 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_X80 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y1 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y2 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y3 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y4 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y6 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y8 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y10 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y20 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y40 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Y80 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z1 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z2 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z3 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z4 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z6 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z8 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z10 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z20 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z40 ();
  output o;
  input a;
  input b;
endmodule

module NOR2_Z80 ();
  output o;
  input a;
  input b;
endmodule

module NOR3_X1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X2 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X3 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X4 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X6 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X8 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_X80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y2 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y3 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y4 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y6 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y8 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Y80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z2 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z3 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z4 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z6 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z8 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z10 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z20 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z40 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR3_Z80 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module NOR4_X1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X2 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X3 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X4 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X6 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X8 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_X80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y2 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y3 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y4 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y6 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y8 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Y80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z2 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z3 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z4 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z6 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z8 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z10 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z20 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z40 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module NOR4_Z80 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module DFF_X80 ();
  output q;
  input ck;
  input d;
endmodule

module BUF_X1 ();
  output o;
  input a;
endmodule

module BUF_X2 ();
  output o;
  input a;
endmodule

module BUF_X3 ();
  output o;
  input a;
endmodule

module BUF_X4 ();
  output o;
  input a;
endmodule

module BUF_X6 ();
  output o;
  input a;
endmodule

module BUF_X8 ();
  output o;
  input a;
endmodule

module BUF_X10 ();
  output o;
  input a;
endmodule

module BUF_X20 ();
  output o;
  input a;
endmodule

module BUF_X40 ();
  output o;
  input a;
endmodule

module BUF_X80 ();
  output o;
  input a;
endmodule

module DFF_X160 ();
  output q;
  input ck;
  input d;
endmodule

module DFFN_X80 ();
  output q;
  input ckn;
  input d;
endmodule

module DFFN_X160 ();
  output q;
  input ckn;
  input d;
endmodule

module OR2_X1 ();
  output o;
  input a;
  input b;
endmodule

module OR3_X1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module OR4_X1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module AND2_X1 ();
  output o;
  input a;
  input b;
endmodule

module AND3_X1 ();
  output o;
  input a;
  input b;
  input c;
endmodule

module AND4_X1 ();
  output o;
  input a;
  input b;
  input c;
  input d;
endmodule

module XOR2_X1 ();
  output o;
  input a;
  input b;
endmodule

module XNOR2_X1 ();
  output o;
  input a;
  input b;
endmodule

module fflopd ();
  input D;
  input CK;
  output Q;
endmodule

module fflopd_2 ();
  input D;
  input CK;
  output Q;
endmodule

module fflopd_3 ();
  input D;
  input CK;
  output Q;
endmodule

module fflopd_ckn ();
  input D;
  input CKN;
  output Q;
endmodule

module fflopd_ckn_2 ();
  input D;
  input CKN;
  output Q;
endmodule

module fflopd_ckn_3 ();
  input D;
  input CKN;
  output Q;
endmodule

