module top;

// Start PIs
input d_6;
input d_0;
input d_5;
input d_1;
input d_8;
input d_15;
input d_12;
input d_3;
input d_13;
input tau_clk;
input d_2;
input d_14;
input d_11;
input d_10;
input d_7;
input d_4;
input d_9;

// Start POs
output crc32N_2;
output crc32N_31;
output crc32N_29;
output crc32N_30;
output crc32N_3;
output crc32N_1;
output crc32N_11;
output crc32N_13;
output crc32N_9;
output crc32N_14;
output crc32N_8;
output crc32N_28;
output crc32N_5;
output crc32N_27;
output crc32N_10;
output crc32N_17;
output crc32N_21;
output crc32N_6;
output crc32N_18;
output crc32N_4;
output crc32N_24;
output crc32N_16;
output crc32N_23;
output crc32N_7;
output crc32N_22;
output crc32N_25;
output crc32N_20;
output crc32N_19;
output crc32N_0;
output crc32N_15;
output crc32N_26;
output crc32N_12;

// Start wires
wire newNet_120;
wire make_crc32d16_n_132;
wire newNet_199;
wire newNet_134;
wire newNet_110;
wire crc32N_2;
wire newNet_10;
wire make_crc32d16_n_272;
wire newNet_166;
wire make_crc32d16_n_73;
wire newNet_191;
wire newNet_130;
wire make_crc32d16_n_53;
wire make_crc32d16_n_186;
wire newNet_24;
wire make_crc32d16_n_38;
wire make_crc32d16_n_41;
wire newNet_7;
wire newNet_170;
wire newNet_79;
wire make_crc32d16_n_153;
wire make_crc32d16_n_87;
wire d_12;
wire newNet_178;
wire make_crc32d16_n_131;
wire newNet_117;
wire newNet_73;
wire newNet_63;
wire crc32_27_;
wire newNet_193;
wire newNet_2;
wire newNet_25;
wire newNet_80;
wire make_crc32d16_n_47;
wire newNet_16;
wire make_crc32d16_n_94;
wire make_crc32d16_n_136;
wire make_crc32d16_n_61;
wire make_crc32d16_n_164;
wire newNet_145;
wire newNet_38;
wire newNet_61;
wire make_crc32d16_n_81;
wire newNet_162;
wire make_crc32d16_n_110;
wire crc32N_23;
wire newNet_155;
wire make_crc32d16_n_4;
wire newNet_124;
wire newNet_149;
wire newNet_101;
wire crc32_26_;
wire d_2;
wire newNet_83;
wire make_crc32d16_n_175;
wire crc32_4_;
wire crc32_8_;
wire make_crc32d16_n_204;
wire newNet_189;
wire newNet_160;
wire make_crc32d16_n_68;
wire newNet_113;
wire crc32_7_;
wire newNet_88;
wire newNet_53;
wire make_crc32d16_n_26;
wire make_crc32d16_n_78;
wire make_crc32d16_n_178;
wire make_crc32d16_n_166;
wire crc32_20_;
wire newNet_92;
wire make_crc32d16_n_98;
wire newNet_19;
wire make_crc32d16_n_64;
wire newNet_57;
wire newNet_26;
wire make_crc32d16_n_105;
wire newNet_76;
wire make_crc32d16_n_189;
wire d_13;
wire make_crc32d16_n_116;
wire newNet_95;
wire newNet_46;
wire crc32N_8;
wire make_crc32d16_n_181;
wire d_10;
wire make_crc32d16_n_42;
wire crc32N_27;
wire newNet_62;
wire newNet_183;
wire newNet_30;
wire newNet_157;
wire newNet_21;
wire newNet_139;
wire make_crc32d16_n_107;
wire make_crc32d16_n_146;
wire newNet_140;
wire make_crc32d16_n_21;
wire newNet_174;
wire crc32_1_;
wire d_6;
wire newNet_13;
wire newNet_99;
wire make_crc32d16_n_15;
wire d_8;
wire crc32N_16;
wire make_crc32d16_n_58;
wire make_crc32d16_n_159;
wire d_15;
wire crc32N_7;
wire make_crc32d16_n_2;
wire make_crc32d16_n_194;
wire crc32N_22;
wire newNet_108;
wire newNet_11;
wire newNet_195;
wire newNet_150;
wire make_crc32d16_n_100;
wire make_crc32d16_n_190;
wire make_crc32d16_n_161;
wire crc32_23_;
wire make_crc32d16_n_28;
wire newNet_123;
wire newNet_67;
wire make_crc32d16_n_172;
wire make_crc32d16_n_7;
wire make_crc32d16_n_91;
wire make_crc32d16_n_152;
wire make_crc32d16_n_257;
wire crc32N_29;
wire newNet_171;
wire crc32_9_;
wire newNet_119;
wire crc32N_3;
wire make_crc32d16_n_79;
wire d_1;
wire newNet_196;
wire make_crc32d16_n_130;
wire make_crc32d16_n_271;
wire make_crc32d16_n_142;
wire newNet_3;
wire make_crc32d16_n_80;
wire newNet_158;
wire make_crc32d16_n_35;
wire make_crc32d16_n_169;
wire make_crc32d16_n_40;
wire make_crc32d16_n_69;
wire newNet_28;
wire make_crc32d16_n_203;
wire newNet_70;
wire make_crc32d16_n_86;
wire newNet_144;
wire newNet_185;
wire make_crc32d16_n_60;
wire newNet_188;
wire newNet_8;
wire make_crc32d16_n_197;
wire make_crc32d16_n_171;
wire newNet_29;
wire make_crc32d16_n_25;
wire make_crc32d16_n_215;
wire newNet_116;
wire make_crc32d16_n_174;
wire newNet_51;
wire newNet_5;
wire newNet_154;
wire newNet_190;
wire newNet_74;
wire newNet_23;
wire d_3;
wire newNet_47;
wire newNet_18;
wire crc32_14_;
wire make_crc32d16_n_65;
wire make_crc32d16_n_134;
wire make_crc32d16_n_206;
wire make_crc32d16_n_137;
wire newNet_41;
wire make_crc32d16_n_230;
wire make_crc32d16_n_156;
wire make_crc32d16_n_11;
wire newNet_15;
wire crc32_16_;
wire newNet_77;
wire newNet_66;
wire newNet_121;
wire newNet_34;
wire make_crc32d16_n_104;
wire make_crc32d16_n_72;
wire make_crc32d16_n_19;
wire newNet_109;
wire newNet_90;
wire newNet_12;
wire newNet_0;
wire make_crc32d16_n_179;
wire newNet_126;
wire newNet_14;
wire make_crc32d16_n_45;
wire newNet_50;
wire make_crc32d16_n_32;
wire newNet_115;
wire newNet_146;
wire tau_clk;
wire newNet_56;
wire crc32N_9;
wire make_crc32d16_n_111;
wire newNet_133;
wire newNet_112;
wire newNet_169;
wire newNet_163;
wire newNet_138;
wire newNet_98;
wire make_crc32d16_n_210;
wire make_crc32d16_n_71;
wire make_crc32d16_n_20;
wire crc32_24_;
wire newNet_137;
wire make_crc32d16_n_128;
wire newNet_165;
wire newNet_27;
wire crc32N_17;
wire crc32N_21;
wire make_crc32d16_n_183;
wire make_crc32d16_n_214;
wire crc32N_4;
wire newNet_184;
wire make_crc32d16_n_36;
wire make_crc32d16_n_57;
wire make_crc32d16_n_198;
wire make_crc32d16_n_18;
wire make_crc32d16_n_112;
wire make_crc32d16_n_138;
wire make_crc32d16_n_160;
wire make_crc32d16_n_209;
wire crc32_15_;
wire make_crc32d16_n_145;
wire newNet_105;
wire newNet_31;
wire make_crc32d16_n_188;
wire newNet_177;
wire newNet_39;
wire newNet_153;
wire crc32_0_;
wire make_crc32d16_n_1;
wire newNet_94;
wire make_crc32d16_n_219;
wire newNet_40;
wire make_crc32d16_n_95;
wire d_7;
wire crc32N_0;
wire newNet_122;
wire make_crc32d16_n_14;
wire crc32N_26;
wire newNet_85;
wire make_crc32d16_n_8;
wire make_crc32d16_n_135;
wire newNet_181;
wire d_0;
wire make_crc32d16_n_63;
wire newNet_6;
wire make_crc32d16_n_177;
wire make_crc32d16_n_168;
wire make_crc32d16_n_217;
wire crc32N_11;
wire newNet_129;
wire newNet_197;
wire newNet_71;
wire make_crc32d16_n_157;
wire make_crc32d16_n_162;
wire crc32N_13;
wire make_crc32d16_n_92;
wire newNet_65;
wire newNet_103;
wire make_crc32d16_n_6;
wire newNet_48;
wire newNet_42;
wire make_crc32d16_n_216;
wire crc32N_28;
wire make_crc32d16_n_221;
wire make_crc32d16_n_76;
wire newNet_36;
wire make_crc32d16_n_201;
wire newNet_182;
wire newNet_161;
wire newNet_4;
wire crc32N_5;
wire newNet_32;
wire d_4;
wire make_crc32d16_n_273;
wire make_crc32d16_n_211;
wire newNet_143;
wire d_9;
wire newNet_107;
wire newNet_172;
wire crc32_29_;
wire make_crc32d16_n_123;
wire newNet_69;
wire make_crc32d16_n_85;
wire make_crc32d16_n_155;
wire make_crc32d16_n_192;
wire crc32_3_;
wire newNet_52;
wire make_crc32d16_n_43;
wire newNet_81;
wire newNet_89;
wire newNet_1;
wire make_crc32d16_n_31;
wire make_crc32d16_n_170;
wire make_crc32d16_n_82;
wire d_14;
wire newNet_9;
wire crc32_30_;
wire newNet_159;
wire make_crc32d16_n_149;
wire make_crc32d16_n_187;
wire make_crc32d16_n_67;
wire make_crc32d16_n_17;
wire newNet_75;
wire make_crc32d16_n_165;
wire crc32N_30;
wire newNet_55;
wire newNet_17;
wire make_crc32d16_n_103;
wire crc32N_1;
wire newNet_147;
wire make_crc32d16_n_75;
wire crc32_18_;
wire newNet_164;
wire newNet_192;
wire make_crc32d16_n_56;
wire make_crc32d16_n_89;
wire make_crc32d16_n_151;
wire crc32_10_;
wire newNet_136;
wire make_crc32d16_n_44;
wire crc32N_10;
wire newNet_102;
wire newNet_168;
wire crc32N_18;
wire newNet_125;
wire crc32_2_;
wire make_crc32d16_n_270;
wire make_crc32d16_n_113;
wire make_crc32d16_n_96;
wire make_crc32d16_n_99;
wire newNet_93;
wire make_crc32d16_n_184;
wire crc32_25_;
wire make_crc32d16_n_127;
wire newNet_127;
wire make_crc32d16_n_182;
wire make_crc32d16_n_102;
wire newNet_82;
wire make_crc32d16_n_266;
wire newNet_132;
wire make_crc32d16_n_140;
wire newNet_33;
wire crc32N_25;
wire make_crc32d16_n_208;
wire make_crc32d16_n_54;
wire crc32N_20;
wire newNet_118;
wire newNet_106;
wire make_crc32d16_n_34;
wire make_crc32d16_n_109;
wire newNet_20;
wire make_crc32d16_n_50;
wire newNet_176;
wire make_crc32d16_n_144;
wire newNet_152;
wire newNet_111;
wire newNet_114;
wire newNet_142;
wire newNet_104;
wire make_crc32d16_n_0;
wire make_crc32d16_n_207;
wire make_crc32d16_n_93;
wire make_crc32d16_n_27;
wire newNet_167;
wire make_crc32d16_n_195;
wire newNet_179;
wire make_crc32d16_n_256;
wire make_crc32d16_n_218;
wire make_crc32d16_n_200;
wire make_crc32d16_n_141;
wire make_crc32d16_n_148;
wire make_crc32d16_n_52;
wire make_crc32d16_n_13;
wire crc32_12_;
wire make_crc32d16_n_122;
wire make_crc32d16_n_205;
wire newNet_198;
wire make_crc32d16_n_9;
wire newNet_135;
wire newNet_35;
wire crc32N_14;
wire make_crc32d16_n_133;
wire make_crc32d16_n_46;
wire make_crc32d16_n_139;
wire make_crc32d16_n_62;
wire crc32_21_;
wire make_crc32d16_n_213;
wire newNet_86;
wire newNet_60;
wire newNet_131;
wire newNet_100;
wire newNet_44;
wire make_crc32d16_n_108;
wire make_crc32d16_n_48;
wire newNet_72;
wire make_crc32d16_n_66;
wire newNet_97;
wire newNet_128;
wire d_5;
wire make_crc32d16_n_10;
wire newNet_186;
wire make_crc32d16_n_154;
wire make_crc32d16_n_83;
wire newNet_45;
wire newNet_37;
wire newNet_173;
wire make_crc32d16_n_70;
wire crc32_19_;
wire newNet_64;
wire crc32_17_;
wire newNet_54;
wire make_crc32d16_n_269;
wire make_crc32d16_n_143;
wire crc32N_19;
wire newNet_78;
wire make_crc32d16_n_51;
wire newNet_49;
wire newNet_180;
wire make_crc32d16_n_39;
wire make_crc32d16_n_274;
wire make_crc32d16_n_55;
wire newNet_43;
wire crc32_28_;
wire crc32N_31;
wire newNet_96;
wire make_crc32d16_n_115;
wire make_crc32d16_n_191;
wire newNet_58;
wire crc32_31_;
wire make_crc32d16_n_59;
wire newNet_91;
wire make_crc32d16_n_129;
wire make_crc32d16_n_97;
wire newNet_148;
wire newNet_22;
wire make_crc32d16_n_150;
wire crc32_22_;
wire newNet_141;
wire d_11;
wire crc32_6_;
wire make_crc32d16_n_106;
wire make_crc32d16_n_30;
wire crc32_5_;
wire make_crc32d16_n_84;
wire make_crc32d16_n_101;
wire make_crc32d16_n_74;
wire make_crc32d16_n_180;
wire make_crc32d16_n_114;
wire make_crc32d16_n_173;
wire newNet_84;
wire make_crc32d16_n_147;
wire crc32N_6;
wire make_crc32d16_n_125;
wire newNet_156;
wire newNet_194;
wire newNet_87;
wire crc32N_24;
wire crc32_13_;
wire make_crc32d16_n_126;
wire newNet_59;
wire make_crc32d16_n_29;
wire newNet_175;
wire make_crc32d16_n_5;
wire make_crc32d16_n_185;
wire make_crc32d16_n_3;
wire make_crc32d16_n_88;
wire newNet_187;
wire make_crc32d16_n_90;
wire make_crc32d16_n_77;
wire make_crc32d16_n_176;
wire make_crc32d16_n_12;
wire make_crc32d16_n_158;
wire crc32_11_;
wire make_crc32d16_n_163;
wire newNet_68;
wire make_crc32d16_n_16;
wire crc32N_15;
wire newNet_151;
wire make_crc32d16_n_167;
wire crc32N_12;

// Start cells
XOR2_X1 make_crc32d16_g2182 ( .a(make_crc32d16_n_3), .b(make_crc32d16_n_70), .o(make_crc32d16_n_90) );
fflopd make_crc32d16_crc_reg_11_ ( .CK(newNet_150), .D(make_crc32d16_n_183), .Q(crc32_11_) );
XOR2_X1 make_crc32d16_g2165 ( .a(make_crc32d16_n_71), .b(make_crc32d16_n_92), .o(make_crc32d16_n_104) );
XOR2_X1 make_crc32d16_g2060 ( .a(make_crc32d16_n_136), .b(make_crc32d16_n_273), .o(make_crc32d16_n_148) );
BUF_X2 newInst_54 ( .a(newNet_53), .o(newNet_54) );
XOR2_X1 make_crc32d16_g2036 ( .a(make_crc32d16_n_162), .b(make_crc32d16_n_139), .o(make_crc32d16_n_174) );
XOR2_X1 make_crc32d16_g2093 ( .a(d_10), .b(d_9), .o(make_crc32d16_n_208) );
XOR2_X1 make_crc32d16_g2079 ( .a(make_crc32d16_n_127), .b(make_crc32d16_n_269), .o(make_crc32d16_n_133) );
INV_Z1 g33 ( .a(crc32_0_), .o(crc32N_31) );
XOR2_X1 make_crc32d16_g2040 ( .a(make_crc32d16_n_157), .b(make_crc32d16_n_126), .o(make_crc32d16_n_173) );
XOR2_X1 make_crc32d16_g2116 ( .a(crc32_29_), .b(crc32_28_), .o(make_crc32d16_n_195) );
BUF_X2 newInst_138 ( .a(newNet_137), .o(newNet_138) );
XOR2_X1 make_crc32d16_g2024 ( .a(make_crc32d16_n_173), .b(make_crc32d16_n_147), .o(make_crc32d16_n_181) );
XOR2_X1 make_crc32d16_g2231 ( .a(make_crc32d16_n_204), .b(crc32_19_), .o(make_crc32d16_n_39) );
INV_Z1 g57 ( .a(crc32_26_), .o(crc32N_5) );
BUF_X2 newInst_3 ( .a(newNet_2), .o(newNet_3) );
INV_Z1 g37 ( .a(crc32_15_), .o(crc32N_16) );
BUF_X2 newInst_74 ( .a(newNet_73), .o(newNet_74) );
INV_X2 newInst_187 ( .a(newNet_186), .o(newNet_187) );
BUF_X2 newInst_68 ( .a(newNet_67), .o(newNet_68) );
XOR2_X1 make_crc32d16_g2189 ( .a(make_crc32d16_n_72), .b(make_crc32d16_n_56), .o(make_crc32d16_n_83) );
XOR2_X1 make_crc32d16_g2084 ( .a(crc32_22_), .b(crc32_20_), .o(make_crc32d16_n_204) );
BUF_X2 newInst_32 ( .a(newNet_31), .o(newNet_32) );
BUF_X2 newInst_79 ( .a(newNet_78), .o(newNet_79) );
XOR2_X1 make_crc32d16_g2055 ( .a(make_crc32d16_n_144), .b(make_crc32d16_n_130), .o(make_crc32d16_n_153) );
BUF_X2 newInst_85 ( .a(newNet_84), .o(newNet_85) );
XOR2_X1 make_crc32d16_g2223 ( .a(d_10), .b(d_6), .o(make_crc32d16_n_46) );
XOR2_X1 make_crc32d16_g2251 ( .a(crc32_20_), .b(d_7), .o(make_crc32d16_n_25) );
XOR2_X1 make_crc32d16_g2065 ( .a(make_crc32d16_n_133), .b(make_crc32d16_n_126), .o(make_crc32d16_n_149) );
BUF_X2 newInst_143 ( .a(newNet_142), .o(newNet_143) );
BUF_X2 newInst_116 ( .a(newNet_45), .o(newNet_116) );
BUF_X2 newInst_2 ( .a(newNet_1), .o(newNet_2) );
BUF_X2 newInst_60 ( .a(newNet_59), .o(newNet_60) );
XOR2_X1 make_crc32d16_g2087 ( .a(d_5), .b(d_2), .o(make_crc32d16_n_266) );
XOR2_X1 make_crc32d16_g2248 ( .a(make_crc32d16_n_206), .b(d_9), .o(make_crc32d16_n_19) );
BUF_X2 newInst_196 ( .a(newNet_195), .o(newNet_196) );
fflopd make_crc32d16_crc_reg_16_ ( .CK(newNet_71), .D(make_crc32d16_n_100), .Q(crc32_16_) );
BUF_X2 newInst_186 ( .a(newNet_185), .o(newNet_186) );
BUF_X2 newInst_36 ( .a(newNet_35), .o(newNet_36) );
XOR2_X1 make_crc32d16_g2121 ( .a(crc32_16_), .b(d_15), .o(make_crc32d16_n_197) );
XOR2_X1 make_crc32d16_g2034 ( .a(make_crc32d16_n_164), .b(make_crc32d16_n_153), .o(make_crc32d16_n_176) );
BUF_X2 newInst_103 ( .a(newNet_102), .o(newNet_103) );
XOR2_X1 make_crc32d16_g2222 ( .a(make_crc32d16_n_219), .b(d_6), .o(make_crc32d16_n_50) );
XOR2_X1 make_crc32d16_g2190 ( .a(make_crc32d16_n_55), .b(make_crc32d16_n_1), .o(make_crc32d16_n_82) );
BUF_X2 newInst_156 ( .a(newNet_155), .o(newNet_156) );
XOR2_X1 make_crc32d16_g2022 ( .a(make_crc32d16_n_173), .b(make_crc32d16_n_144), .o(make_crc32d16_n_183) );
fflopd make_crc32d16_crc_reg_3_ ( .CK(newNet_188), .D(make_crc32d16_n_191), .Q(crc32_3_) );
BUF_X2 newInst_7 ( .a(newNet_6), .o(newNet_7) );
BUF_X2 newInst_159 ( .a(newNet_158), .o(newNet_159) );
XOR2_X1 make_crc32d16_g2256 ( .a(crc32_4_), .b(d_11), .o(make_crc32d16_n_13) );
XOR2_X1 make_crc32d16_g2209 ( .a(make_crc32d16_n_36), .b(make_crc32d16_n_48), .o(make_crc32d16_n_63) );
INV_Z1 g43 ( .a(crc32_4_), .o(crc32N_27) );
XOR2_X1 make_crc32d16_g2230 ( .a(crc32_24_), .b(crc32_9_), .o(make_crc32d16_n_40) );
fflopd make_crc32d16_crc_reg_6_ ( .CK(newNet_196), .D(make_crc32d16_n_190), .Q(crc32_6_) );
BUF_X2 newInst_173 ( .a(newNet_172), .o(newNet_173) );
XOR2_X1 make_crc32d16_g2066 ( .a(make_crc32d16_n_129), .b(make_crc32d16_n_130), .o(make_crc32d16_n_143) );
BUF_X2 newInst_108 ( .a(newNet_107), .o(newNet_108) );
XOR2_X1 make_crc32d16_g2076 ( .a(make_crc32d16_n_128), .b(d_1), .o(make_crc32d16_n_230) );
INV_Z1 g60 ( .a(crc32_27_), .o(crc32N_4) );
BUF_X2 newInst_58 ( .a(newNet_57), .o(newNet_58) );
BUF_X2 newInst_43 ( .a(newNet_42), .o(newNet_43) );
BUF_X2 newInst_73 ( .a(newNet_38), .o(newNet_73) );
BUF_X2 newInst_26 ( .a(newNet_25), .o(newNet_26) );
XOR2_X1 make_crc32d16_g2194 ( .a(make_crc32d16_n_43), .b(make_crc32d16_n_16), .o(make_crc32d16_n_78) );
XOR2_X1 make_crc32d16_g2247 ( .a(d_13), .b(d_12), .o(make_crc32d16_n_20) );
XOR2_X1 make_crc32d16_g2080 ( .a(make_crc32d16_n_273), .b(make_crc32d16_n_122), .o(make_crc32d16_n_135) );
BUF_X2 newInst_16 ( .a(newNet_6), .o(newNet_16) );
XOR2_X1 make_crc32d16_g2187 ( .a(make_crc32d16_n_8), .b(make_crc32d16_n_58), .o(make_crc32d16_n_85) );
XOR2_X1 make_crc32d16_g2098 ( .a(d_6), .b(d_2), .o(make_crc32d16_n_128) );
INV_Z1 g54 ( .a(crc32_24_), .o(crc32N_7) );
BUF_X2 newInst_65 ( .a(newNet_64), .o(newNet_65) );
BUF_X2 newInst_169 ( .a(newNet_168), .o(newNet_169) );
BUF_X2 newInst_131 ( .a(newNet_130), .o(newNet_131) );
XOR2_X1 make_crc32d16_g2243 ( .a(make_crc32d16_n_205), .b(d_9), .o(make_crc32d16_n_28) );
fflopd make_crc32d16_crc_reg_12_ ( .CK(newNet_159), .D(make_crc32d16_n_181), .Q(crc32_12_) );
BUF_X2 newInst_13 ( .a(newNet_12), .o(newNet_13) );
BUF_X2 newInst_150 ( .a(newNet_149), .o(newNet_150) );
XOR2_X1 make_crc32d16_g2145 ( .a(make_crc32d16_n_108), .b(make_crc32d16_n_57), .o(make_crc32d16_n_113) );
BUF_X2 newInst_142 ( .a(newNet_141), .o(newNet_142) );
BUF_X2 newInst_37 ( .a(newNet_36), .o(newNet_37) );
BUF_X2 newInst_146 ( .a(newNet_145), .o(newNet_146) );
fflopd make_crc32d16_crc_reg_29_ ( .CK(newNet_41), .D(make_crc32d16_n_99), .Q(crc32_29_) );
fflopd make_crc32d16_crc_reg_19_ ( .CK(newNet_111), .D(make_crc32d16_n_114), .Q(crc32_19_) );
BUF_X2 newInst_12 ( .a(newNet_11), .o(newNet_12) );
BUF_X2 newInst_88 ( .a(newNet_87), .o(newNet_88) );
XOR2_X1 make_crc32d16_g2105 ( .a(crc32_21_), .b(d_10), .o(make_crc32d16_n_125) );
fflopd make_crc32d16_crc_reg_26_ ( .CK(newNet_62), .D(make_crc32d16_n_104), .Q(crc32_26_) );
XOR2_X1 make_crc32d16_g2163 ( .a(make_crc32d16_n_95), .b(make_crc32d16_n_12), .o(make_crc32d16_n_106) );
BUF_X2 newInst_134 ( .a(newNet_108), .o(newNet_134) );
XOR2_X1 make_crc32d16_g2272 ( .a(make_crc32d16_n_266), .b(crc32_5_), .o(make_crc32d16_n_0) );
XOR2_X1 make_crc32d16_g2152 ( .a(make_crc32d16_n_101), .b(d_10), .o(make_crc32d16_n_108) );
XOR2_X1 make_crc32d16_g2070 ( .a(make_crc32d16_n_269), .b(make_crc32d16_n_272), .o(make_crc32d16_n_144) );
XOR2_X1 make_crc32d16_g2205 ( .a(make_crc32d16_n_35), .b(make_crc32d16_n_5), .o(make_crc32d16_n_67) );
XOR2_X1 make_crc32d16_g2101 ( .a(crc32_23_), .b(d_8), .o(make_crc32d16_n_129) );
XOR2_X1 make_crc32d16_g2166 ( .a(make_crc32d16_n_91), .b(make_crc32d16_n_48), .o(make_crc32d16_n_103) );
INV_Z1 g47 ( .a(crc32_10_), .o(crc32N_21) );
BUF_X2 newInst_17 ( .a(newNet_16), .o(newNet_17) );
BUF_X2 newInst_104 ( .a(newNet_103), .o(newNet_104) );
BUF_X2 newInst_21 ( .a(newNet_20), .o(newNet_21) );
XOR2_X1 make_crc32d16_g2045 ( .a(make_crc32d16_n_156), .b(make_crc32d16_n_273), .o(make_crc32d16_n_166) );
BUF_X2 newInst_177 ( .a(newNet_176), .o(newNet_177) );
XOR2_X1 make_crc32d16_g2268 ( .a(make_crc32d16_n_221), .b(crc32_2_), .o(make_crc32d16_n_3) );
BUF_X2 newInst_111 ( .a(newNet_110), .o(newNet_111) );
XOR2_X1 make_crc32d16_g2052 ( .a(make_crc32d16_n_151), .b(make_crc32d16_n_139), .o(make_crc32d16_n_157) );
BUF_X2 newInst_49 ( .a(newNet_48), .o(newNet_49) );
XOR2_X1 make_crc32d16_g2058 ( .a(make_crc32d16_n_139), .b(make_crc32d16_n_129), .o(make_crc32d16_n_152) );
BUF_X2 newInst_149 ( .a(newNet_148), .o(newNet_149) );
XOR2_X1 make_crc32d16_g2203 ( .a(make_crc32d16_n_271), .b(crc32_10_), .o(make_crc32d16_n_69) );
BUF_X2 newInst_181 ( .a(newNet_180), .o(newNet_181) );
BUF_X2 newInst_83 ( .a(newNet_82), .o(newNet_83) );
fflopd make_crc32d16_crc_reg_27_ ( .CK(newNet_88), .D(make_crc32d16_n_110), .Q(crc32_27_) );
XOR2_X1 make_crc32d16_g2017 ( .a(make_crc32d16_n_177), .b(make_crc32d16_n_143), .o(make_crc32d16_n_188) );
BUF_X2 newInst_80 ( .a(newNet_79), .o(newNet_80) );
XOR2_X1 make_crc32d16_g2271 ( .a(crc32_16_), .b(d_15), .o(make_crc32d16_n_21) );
BUF_X2 newInst_20 ( .a(newNet_19), .o(newNet_20) );
XOR2_X1 make_crc32d16_g2204 ( .a(make_crc32d16_n_6), .b(make_crc32d16_n_274), .o(make_crc32d16_n_68) );
XOR2_X1 make_crc32d16_g2114 ( .a(crc32_28_), .b(crc32_27_), .o(make_crc32d16_n_200) );
XOR2_X1 make_crc32d16_g2083 ( .a(crc32_22_), .b(crc32_21_), .o(make_crc32d16_n_205) );
BUF_X2 newInst_124 ( .a(newNet_123), .o(newNet_124) );
XOR2_X1 make_crc32d16_g2244 ( .a(crc32_23_), .b(d_8), .o(make_crc32d16_n_47) );
INV_Z1 g49 ( .a(crc32_22_), .o(crc32N_9) );
BUF_X2 newInst_97 ( .a(newNet_96), .o(newNet_97) );
fflopd make_crc32d16_crc_reg_4_ ( .CK(newNet_124), .D(make_crc32d16_n_171), .Q(crc32_4_) );
XOR2_X1 make_crc32d16_g2109 ( .a(d_14), .b(d_13), .o(make_crc32d16_n_214) );
XOR2_X1 make_crc32d16_g2035 ( .a(make_crc32d16_n_165), .b(make_crc32d16_n_166), .o(make_crc32d16_n_175) );
XOR2_X1 make_crc32d16_g2162 ( .a(make_crc32d16_n_90), .b(make_crc32d16_n_74), .o(make_crc32d16_n_107) );
XOR2_X1 make_crc32d16_g2011 ( .a(make_crc32d16_n_182), .b(make_crc32d16_n_125), .o(make_crc32d16_n_189) );
BUF_X2 newInst_165 ( .a(newNet_164), .o(newNet_165) );
BUF_X2 newInst_29 ( .a(newNet_28), .o(newNet_29) );
fflopd make_crc32d16_crc_reg_24_ ( .CK(newNet_72), .D(make_crc32d16_n_105), .Q(crc32_24_) );
XOR2_X1 make_crc32d16_g2075 ( .a(make_crc32d16_n_125), .b(make_crc32d16_n_131), .o(make_crc32d16_n_137) );
XOR2_X1 make_crc32d16_g2019 ( .a(make_crc32d16_n_179), .b(make_crc32d16_n_272), .o(make_crc32d16_n_186) );
BUF_X2 newInst_110 ( .a(newNet_109), .o(newNet_110) );
INV_Z1 g41 ( .a(crc32_17_), .o(crc32N_14) );
BUF_X2 newInst_137 ( .a(newNet_136), .o(newNet_137) );
XOR2_X1 make_crc32d16_g2232 ( .a(crc32_31_), .b(d_8), .o(make_crc32d16_n_38) );
XOR2_X1 make_crc32d16_g2226 ( .a(crc32_25_), .b(crc32_30_), .o(make_crc32d16_n_44) );
INV_Z1 g51 ( .a(crc32_5_), .o(crc32N_26) );
BUF_X2 newInst_24 ( .a(newNet_23), .o(newNet_24) );
BUF_X2 newInst_86 ( .a(newNet_85), .o(newNet_86) );
XOR2_X1 make_crc32d16_g2171 ( .a(make_crc32d16_n_85), .b(make_crc32d16_n_59), .o(make_crc32d16_n_98) );
BUF_X2 newInst_117 ( .a(newNet_63), .o(newNet_117) );
fflopd make_crc32d16_crc_reg_23_ ( .CK(newNet_9), .D(make_crc32d16_n_112), .Q(crc32_23_) );
fflopd make_crc32d16_crc_reg_2_ ( .CK(newNet_179), .D(make_crc32d16_n_192), .Q(crc32_2_) );
XOR2_X1 make_crc32d16_g2039 ( .a(make_crc32d16_n_161), .b(make_crc32d16_n_122), .o(make_crc32d16_n_170) );
XOR2_X1 make_crc32d16_g2164 ( .a(make_crc32d16_n_94), .b(make_crc32d16_n_76), .o(make_crc32d16_n_105) );
XOR2_X1 make_crc32d16_g2023 ( .a(make_crc32d16_n_179), .b(make_crc32d16_n_145), .o(make_crc32d16_n_182) );
BUF_X2 newInst_59 ( .a(newNet_58), .o(newNet_59) );
BUF_X2 newInst_69 ( .a(newNet_68), .o(newNet_69) );
BUF_X2 newInst_48 ( .a(newNet_20), .o(newNet_48) );
BUF_X2 newInst_10 ( .a(newNet_8), .o(newNet_10) );
fflopd make_crc32d16_crc_reg_0_ ( .CK(newNet_15), .D(make_crc32d16_n_88), .Q(crc32_0_) );
BUF_X2 newInst_168 ( .a(newNet_167), .o(newNet_168) );
XOR2_X1 make_crc32d16_g2255 ( .a(make_crc32d16_n_200), .b(crc32_6_), .o(make_crc32d16_n_14) );
XOR2_X1 make_crc32d16_g2249 ( .a(make_crc32d16_n_203), .b(d_12), .o(make_crc32d16_n_18) );
BUF_X2 newInst_171 ( .a(newNet_170), .o(newNet_171) );
XOR2_X1 make_crc32d16_g2191 ( .a(make_crc32d16_n_14), .b(make_crc32d16_n_80), .o(make_crc32d16_n_81) );
XOR2_X1 make_crc32d16_g2008 ( .a(make_crc32d16_n_187), .b(make_crc32d16_n_142), .o(make_crc32d16_n_192) );
BUF_X2 newInst_129 ( .a(newNet_128), .o(newNet_129) );
fflopd make_crc32d16_crc_reg_17_ ( .CK(newNet_61), .D(make_crc32d16_n_97), .Q(crc32_17_) );
BUF_X2 newInst_28 ( .a(newNet_27), .o(newNet_28) );
INV_Z1 g40 ( .a(crc32_8_), .o(crc32N_23) );
XOR2_X1 make_crc32d16_g2056 ( .a(make_crc32d16_n_145), .b(make_crc32d16_n_132), .o(make_crc32d16_n_156) );
XOR2_X1 make_crc32d16_g2229 ( .a(make_crc32d16_n_198), .b(crc32_30_), .o(make_crc32d16_n_41) );
BUF_X2 newInst_55 ( .a(newNet_54), .o(newNet_55) );
BUF_X2 newInst_6 ( .a(newNet_5), .o(newNet_6) );
XOR2_X1 make_crc32d16_g2021 ( .a(make_crc32d16_n_172), .b(make_crc32d16_n_125), .o(make_crc32d16_n_184) );
fflopd make_crc32d16_crc_reg_8_ ( .CK(newNet_133), .D(make_crc32d16_n_178), .Q(crc32_8_) );
XOR2_X1 make_crc32d16_g2033 ( .a(make_crc32d16_n_167), .b(make_crc32d16_n_125), .o(make_crc32d16_n_177) );
XOR2_X1 make_crc32d16_g2224 ( .a(d_6), .b(d_4), .o(make_crc32d16_n_45) );
XOR2_X1 make_crc32d16_g2054 ( .a(make_crc32d16_n_150), .b(make_crc32d16_n_137), .o(make_crc32d16_n_161) );
BUF_X2 newInst_170 ( .a(newNet_29), .o(newNet_170) );
BUF_X2 newInst_53 ( .a(newNet_52), .o(newNet_53) );
BUF_X2 newInst_33 ( .a(newNet_32), .o(newNet_33) );
XOR2_X1 make_crc32d16_g2199 ( .a(make_crc32d16_n_40), .b(make_crc32d16_n_20), .o(make_crc32d16_n_73) );
BUF_X2 newInst_114 ( .a(newNet_113), .o(newNet_114) );
BUF_X2 newInst_19 ( .a(newNet_18), .o(newNet_19) );
XOR2_X1 make_crc32d16_g2208 ( .a(make_crc32d16_n_274), .b(crc32_12_), .o(make_crc32d16_n_64) );
BUF_X2 newInst_162 ( .a(newNet_161), .o(newNet_162) );
XOR2_X1 make_crc32d16_g2097 ( .a(d_2), .b(d_0), .o(make_crc32d16_n_256) );
XOR2_X1 make_crc32d16_g2236 ( .a(crc32_21_), .b(d_7), .o(make_crc32d16_n_34) );
XOR2_X1 make_crc32d16_g2181 ( .a(make_crc32d16_n_67), .b(make_crc32d16_n_273), .o(make_crc32d16_n_91) );
BUF_X2 newInst_96 ( .a(newNet_95), .o(newNet_96) );
XOR2_X1 make_crc32d16_g2240 ( .a(make_crc32d16_n_218), .b(crc32_21_), .o(make_crc32d16_n_48) );
XOR2_X1 make_crc32d16_g2220 ( .a(make_crc32d16_n_28), .b(make_crc32d16_n_44), .o(make_crc32d16_n_52) );
XOR2_X1 make_crc32d16_g2049 ( .a(make_crc32d16_n_149), .b(make_crc32d16_n_151), .o(make_crc32d16_n_160) );
BUF_X2 newInst_157 ( .a(newNet_156), .o(newNet_157) );
XOR2_X1 make_crc32d16_g2221 ( .a(crc32_29_), .b(d_6), .o(make_crc32d16_n_51) );
BUF_X2 newInst_197 ( .a(newNet_153), .o(newNet_197) );
XOR2_X1 make_crc32d16_g2067 ( .a(make_crc32d16_n_127), .b(make_crc32d16_n_131), .o(make_crc32d16_n_142) );
BUF_X2 newInst_132 ( .a(newNet_131), .o(newNet_132) );
XOR2_X1 make_crc32d16_g2215 ( .a(make_crc32d16_n_50), .b(make_crc32d16_n_30), .o(make_crc32d16_n_57) );
BUF_X2 newInst_145 ( .a(newNet_144), .o(newNet_145) );
INV_X2 newInst_93 ( .a(newNet_92), .o(newNet_93) );
XOR2_X1 make_crc32d16_g2196 ( .a(make_crc32d16_n_272), .b(make_crc32d16_n_42), .o(make_crc32d16_n_76) );
XOR2_X1 make_crc32d16_g2259 ( .a(crc32_7_), .b(d_15), .o(make_crc32d16_n_10) );
BUF_X2 newInst_122 ( .a(newNet_121), .o(newNet_122) );
BUF_X2 newInst_84 ( .a(newNet_18), .o(newNet_84) );
XOR2_X1 make_crc32d16_g2195 ( .a(make_crc32d16_n_9), .b(crc32_31_), .o(make_crc32d16_n_77) );
XOR2_X1 make_crc32d16_g2150 ( .a(make_crc32d16_n_103), .b(make_crc32d16_n_47), .o(make_crc32d16_n_110) );
BUF_X2 newInst_176 ( .a(newNet_175), .o(newNet_176) );
BUF_X2 newInst_109 ( .a(newNet_108), .o(newNet_109) );
XOR2_X1 make_crc32d16_g2062 ( .a(make_crc32d16_n_137), .b(make_crc32d16_n_136), .o(make_crc32d16_n_147) );
BUF_X2 newInst_128 ( .a(newNet_127), .o(newNet_128) );
XOR2_X1 make_crc32d16_g2018 ( .a(make_crc32d16_n_174), .b(make_crc32d16_n_197), .o(make_crc32d16_n_187) );
BUF_X2 newInst_125 ( .a(newNet_102), .o(newNet_125) );
INV_Z1 g46 ( .a(crc32_20_), .o(crc32N_11) );
BUF_X2 newInst_25 ( .a(newNet_24), .o(newNet_25) );
fflopd make_crc32d16_crc_reg_28_ ( .CK(newNet_47), .D(make_crc32d16_n_102), .Q(crc32_28_) );
BUF_X2 newInst_42 ( .a(newNet_22), .o(newNet_42) );
BUF_X2 newInst_135 ( .a(newNet_134), .o(newNet_135) );
BUF_X2 newInst_4 ( .a(newNet_3), .o(newNet_4) );
XOR2_X1 make_crc32d16_g2263 ( .a(make_crc32d16_n_209), .b(make_crc32d16_n_194), .o(make_crc32d16_n_6) );
INV_Z1 g58 ( .a(crc32_6_), .o(crc32N_25) );
XOR2_X1 make_crc32d16_g2051 ( .a(make_crc32d16_n_155), .b(make_crc32d16_n_135), .o(make_crc32d16_n_158) );
BUF_X2 newInst_52 ( .a(newNet_51), .o(newNet_52) );
BUF_X2 newInst_64 ( .a(newNet_63), .o(newNet_64) );
BUF_X2 newInst_102 ( .a(newNet_71), .o(newNet_102) );
XOR2_X1 make_crc32d16_g2044 ( .a(make_crc32d16_n_149), .b(make_crc32d16_n_138), .o(make_crc32d16_n_167) );
BUF_X2 newInst_105 ( .a(newNet_104), .o(newNet_105) );
XOR2_X1 make_crc32d16_g2235 ( .a(crc32_17_), .b(crc32_20_), .o(make_crc32d16_n_35) );
BUF_X2 newInst_0 ( .a(tau_clk), .o(newNet_0) );
fflopd make_crc32d16_crc_reg_21_ ( .CK(newNet_90), .D(make_crc32d16_n_82), .Q(crc32_21_) );
XOR2_X1 make_crc32d16_g2078 ( .a(make_crc32d16_n_269), .b(make_crc32d16_n_123), .o(make_crc32d16_n_134) );
XOR2_X1 make_crc32d16_g2179 ( .a(make_crc32d16_n_11), .b(make_crc32d16_n_78), .o(make_crc32d16_n_93) );
XOR2_X1 make_crc32d16_g2169 ( .a(make_crc32d16_n_87), .b(crc32_31_), .o(make_crc32d16_n_101) );
XOR2_X1 make_crc32d16_g2102 ( .a(crc32_24_), .b(d_7), .o(make_crc32d16_n_127) );
BUF_X2 newInst_70 ( .a(newNet_69), .o(newNet_70) );
XOR2_X1 make_crc32d16_g2210 ( .a(make_crc32d16_n_4), .b(make_crc32d16_n_31), .o(make_crc32d16_n_62) );
XOR2_X1 make_crc32d16_g2086 ( .a(crc32_22_), .b(crc32_23_), .o(make_crc32d16_n_198) );
XOR2_X1 make_crc32d16_g2092 ( .a(crc32_25_), .b(d_6), .o(make_crc32d16_n_130) );
INV_Z1 g55 ( .a(crc32_12_), .o(crc32N_19) );
XOR2_X1 make_crc32d16_g2276 ( .a(crc32_30_), .b(d_1), .o(make_crc32d16_n_272) );
XOR2_X1 make_crc32d16_g2186 ( .a(make_crc32d16_n_60), .b(make_crc32d16_n_18), .o(make_crc32d16_n_86) );
XOR2_X1 make_crc32d16_g2071 ( .a(make_crc32d16_n_127), .b(make_crc32d16_n_123), .o(make_crc32d16_n_140) );
BUF_X2 newInst_81 ( .a(newNet_80), .o(newNet_81) );
XOR2_X1 make_crc32d16_g2057 ( .a(make_crc32d16_n_139), .b(make_crc32d16_n_274), .o(make_crc32d16_n_155) );
BUF_X2 newInst_87 ( .a(newNet_86), .o(newNet_87) );
BUF_X2 newInst_18 ( .a(newNet_17), .o(newNet_18) );
INV_Z1 g42 ( .a(crc32_18_), .o(crc32N_13) );
XOR2_X1 make_crc32d16_g2239 ( .a(crc32_19_), .b(crc32_22_), .o(make_crc32d16_n_31) );
XOR2_X1 make_crc32d16_g2217 ( .a(make_crc32d16_n_0), .b(make_crc32d16_n_46), .o(make_crc32d16_n_55) );
BUF_X2 newInst_76 ( .a(newNet_75), .o(newNet_76) );
fflopd make_crc32d16_crc_reg_20_ ( .CK(newNet_26), .D(make_crc32d16_n_83), .Q(crc32_20_) );
fflopd make_crc32d16_crc_reg_10_ ( .CK(newNet_116), .D(make_crc32d16_n_176), .Q(crc32_10_) );
XOR2_X1 make_crc32d16_g2082 ( .a(crc32_22_), .b(crc32_24_), .o(make_crc32d16_n_207) );
XOR2_X1 make_crc32d16_g2148 ( .a(make_crc32d16_n_106), .b(make_crc32d16_n_51), .o(make_crc32d16_n_112) );
BUF_X2 newInst_14 ( .a(newNet_13), .o(newNet_14) );
XOR2_X1 make_crc32d16_g2257 ( .a(make_crc32d16_n_209), .b(make_crc32d16_n_210), .o(make_crc32d16_n_12) );
XOR2_X1 make_crc32d16_g2053 ( .a(make_crc32d16_n_146), .b(make_crc32d16_n_272), .o(make_crc32d16_n_162) );
BUF_X2 newInst_11 ( .a(newNet_10), .o(newNet_11) );
BUF_X2 newInst_193 ( .a(newNet_192), .o(newNet_193) );
INV_Z1 g39 ( .a(crc32_16_), .o(crc32N_15) );
BUF_X2 newInst_175 ( .a(newNet_174), .o(newNet_175) );
BUF_X2 newInst_45 ( .a(newNet_44), .o(newNet_45) );
BUF_X2 newInst_63 ( .a(newNet_7), .o(newNet_63) );
INV_Z1 g52 ( .a(crc32_11_), .o(crc32N_20) );
XOR2_X1 make_crc32d16_g2089 ( .a(d_3), .b(d_2), .o(make_crc32d16_n_257) );
XOR2_X1 make_crc32d16_g2108 ( .a(d_5), .b(d_1), .o(make_crc32d16_n_116) );
XOR2_X1 make_crc32d16_g2185 ( .a(make_crc32d16_n_61), .b(d_0), .o(make_crc32d16_n_87) );
XOR2_X1 make_crc32d16_g2273 ( .a(crc32_19_), .b(d_12), .o(make_crc32d16_n_269) );
INV_Z1 g45 ( .a(crc32_19_), .o(crc32N_12) );
XOR2_X1 make_crc32d16_g2173 ( .a(make_crc32d16_n_81), .b(make_crc32d16_n_53), .o(make_crc32d16_n_96) );
XOR2_X1 make_crc32d16_g2168 ( .a(make_crc32d16_n_63), .b(make_crc32d16_n_84), .o(make_crc32d16_n_100) );
BUF_X2 newInst_180 ( .a(newNet_166), .o(newNet_180) );
BUF_X2 newInst_178 ( .a(newNet_177), .o(newNet_178) );
BUF_X2 newInst_164 ( .a(newNet_163), .o(newNet_164) );
BUF_X2 newInst_50 ( .a(newNet_49), .o(newNet_50) );
BUF_X2 newInst_172 ( .a(newNet_171), .o(newNet_172) );
BUF_X2 newInst_167 ( .a(newNet_166), .o(newNet_167) );
INV_Z1 g35 ( .a(crc32_3_), .o(crc32N_28) );
XOR2_X1 make_crc32d16_g2180 ( .a(make_crc32d16_n_69), .b(make_crc32d16_n_19), .o(make_crc32d16_n_92) );
XOR2_X1 make_crc32d16_g2245 ( .a(d_11), .b(d_8), .o(make_crc32d16_n_27) );
XOR2_X1 make_crc32d16_g2009 ( .a(make_crc32d16_n_186), .b(make_crc32d16_n_152), .o(make_crc32d16_n_191) );
BUF_X2 newInst_67 ( .a(newNet_66), .o(newNet_67) );
XOR2_X1 make_crc32d16_g2254 ( .a(crc32_25_), .b(d_3), .o(make_crc32d16_n_15) );
BUF_X2 newInst_34 ( .a(newNet_7), .o(newNet_34) );
BUF_X2 newInst_77 ( .a(newNet_76), .o(newNet_77) );
BUF_X2 newInst_23 ( .a(newNet_22), .o(newNet_23) );
XOR2_X1 make_crc32d16_g2068 ( .a(make_crc32d16_n_127), .b(make_crc32d16_n_273), .o(make_crc32d16_n_141) );
XOR2_X1 make_crc32d16_g2096 ( .a(crc32_25_), .b(crc32_21_), .o(make_crc32d16_n_216) );
XOR2_X1 make_crc32d16_g2246 ( .a(crc32_26_), .b(d_9), .o(make_crc32d16_n_26) );
XOR2_X1 make_crc32d16_g2032 ( .a(make_crc32d16_n_159), .b(make_crc32d16_n_141), .o(make_crc32d16_n_178) );
XOR2_X1 make_crc32d16_g2228 ( .a(crc32_17_), .b(crc32_18_), .o(make_crc32d16_n_42) );
INV_Z1 g59 ( .a(crc32_13_), .o(crc32N_18) );
XOR2_X1 make_crc32d16_g2197 ( .a(make_crc32d16_n_271), .b(make_crc32d16_n_47), .o(make_crc32d16_n_75) );
XOR2_X1 make_crc32d16_g2238 ( .a(make_crc32d16_n_207), .b(crc32_18_), .o(make_crc32d16_n_32) );
BUF_X2 newInst_121 ( .a(newNet_120), .o(newNet_121) );
INV_Z1 g44 ( .a(crc32_9_), .o(crc32N_22) );
XOR2_X1 make_crc32d16_g2091 ( .a(crc32_29_), .b(d_2), .o(make_crc32d16_n_131) );
XOR2_X1 make_crc32d16_g2207 ( .a(make_crc32d16_n_32), .b(make_crc32d16_n_34), .o(make_crc32d16_n_65) );
BUF_X2 newInst_98 ( .a(newNet_97), .o(newNet_98) );
BUF_X2 newInst_30 ( .a(newNet_29), .o(newNet_30) );
BUF_X2 newInst_27 ( .a(tau_clk), .o(newNet_27) );
BUF_X2 newInst_113 ( .a(newNet_112), .o(newNet_113) );
XOR2_X1 make_crc32d16_g2074 ( .a(make_crc32d16_n_122), .b(make_crc32d16_n_274), .o(make_crc32d16_n_138) );
XOR2_X1 make_crc32d16_g2048 ( .a(make_crc32d16_n_149), .b(make_crc32d16_n_270), .o(make_crc32d16_n_163) );
XOR2_X1 make_crc32d16_g2201 ( .a(make_crc32d16_n_39), .b(make_crc32d16_n_21), .o(make_crc32d16_n_71) );
BUF_X2 newInst_56 ( .a(newNet_55), .o(newNet_56) );
XOR2_X1 make_crc32d16_g2010 ( .a(make_crc32d16_n_184), .b(make_crc32d16_n_140), .o(make_crc32d16_n_190) );
XOR2_X1 make_crc32d16_g2095 ( .a(crc32_25_), .b(crc32_23_), .o(make_crc32d16_n_201) );
BUF_X2 newInst_136 ( .a(newNet_135), .o(newNet_136) );
BUF_X2 newInst_39 ( .a(newNet_38), .o(newNet_39) );
XOR2_X1 make_crc32d16_g2107 ( .a(d_11), .b(d_10), .o(make_crc32d16_n_218) );
BUF_X2 newInst_71 ( .a(newNet_70), .o(newNet_71) );
XOR2_X1 make_crc32d16_g2063 ( .a(make_crc32d16_n_136), .b(make_crc32d16_n_129), .o(make_crc32d16_n_146) );
XOR2_X1 make_crc32d16_g2192 ( .a(make_crc32d16_n_272), .b(make_crc32d16_n_21), .o(make_crc32d16_n_80) );
BUF_X2 newInst_158 ( .a(newNet_157), .o(newNet_158) );
BUF_X2 newInst_184 ( .a(newNet_183), .o(newNet_184) );
XOR2_X1 make_crc32d16_g2085 ( .a(crc32_22_), .b(d_9), .o(make_crc32d16_n_132) );
BUF_X2 newInst_90 ( .a(newNet_89), .o(newNet_90) );
fflopd make_crc32d16_crc_reg_7_ ( .CK(newNet_199), .D(make_crc32d16_n_189), .Q(crc32_7_) );
INV_Z1 g62 ( .a(crc32_14_), .o(crc32N_17) );
XOR2_X1 make_crc32d16_g2111 ( .a(crc32_17_), .b(d_14), .o(make_crc32d16_n_123) );
XOR2_X1 make_crc32d16_g2213 ( .a(make_crc32d16_n_25), .b(make_crc32d16_n_27), .o(make_crc32d16_n_59) );
XOR2_X1 make_crc32d16_g2277 ( .a(crc32_27_), .b(d_4), .o(make_crc32d16_n_273) );
XOR2_X1 make_crc32d16_g2072 ( .a(make_crc32d16_n_116), .b(d_0), .o(make_crc32d16_n_221) );
BUF_X2 newInst_153 ( .a(newNet_152), .o(newNet_153) );
XOR2_X1 make_crc32d16_g2103 ( .a(crc32_31_), .b(d_0), .o(make_crc32d16_n_126) );
BUF_X2 newInst_5 ( .a(newNet_4), .o(newNet_5) );
BUF_X2 newInst_8 ( .a(newNet_7), .o(newNet_8) );
XOR2_X1 make_crc32d16_g2120 ( .a(crc32_17_), .b(crc32_16_), .o(make_crc32d16_n_210) );
BUF_X2 newInst_179 ( .a(newNet_178), .o(newNet_179) );
INV_Z1 g34 ( .a(crc32_1_), .o(crc32N_30) );
BUF_X2 newInst_101 ( .a(newNet_100), .o(newNet_101) );
BUF_X2 newInst_62 ( .a(newNet_19), .o(newNet_62) );
XOR2_X1 make_crc32d16_g2200 ( .a(make_crc32d16_n_50), .b(make_crc32d16_n_13), .o(make_crc32d16_n_72) );
XOR2_X1 make_crc32d16_g2214 ( .a(make_crc32d16_n_271), .b(make_crc32d16_n_272), .o(make_crc32d16_n_58) );
BUF_X2 newInst_106 ( .a(newNet_105), .o(newNet_106) );
XOR2_X1 make_crc32d16_g2059 ( .a(make_crc32d16_n_137), .b(make_crc32d16_n_270), .o(make_crc32d16_n_154) );
XOR2_X1 make_crc32d16_g2258 ( .a(make_crc32d16_n_230), .b(crc32_1_), .o(make_crc32d16_n_11) );
BUF_X2 newInst_151 ( .a(newNet_36), .o(newNet_151) );
BUF_X2 newInst_1 ( .a(newNet_0), .o(newNet_1) );
INV_X2 newInst_140 ( .a(newNet_139), .o(newNet_140) );
BUF_X2 newInst_163 ( .a(newNet_162), .o(newNet_163) );
INV_Z1 g63 ( .a(crc32_29_), .o(crc32N_2) );
XOR2_X1 make_crc32d16_g2043 ( .a(make_crc32d16_n_162), .b(make_crc32d16_n_135), .o(make_crc32d16_n_172) );
BUF_X2 newInst_192 ( .a(newNet_191), .o(newNet_192) );
BUF_X2 newInst_89 ( .a(newNet_68), .o(newNet_89) );
XOR2_X1 make_crc32d16_g2261 ( .a(make_crc32d16_n_217), .b(crc32_14_), .o(make_crc32d16_n_8) );
XOR2_X1 make_crc32d16_g2262 ( .a(make_crc32d16_n_214), .b(crc32_8_), .o(make_crc32d16_n_7) );
XOR2_X1 make_crc32d16_g2042 ( .a(make_crc32d16_n_162), .b(make_crc32d16_n_161), .o(make_crc32d16_n_168) );
XOR2_X1 make_crc32d16_g2218 ( .a(make_crc32d16_n_25), .b(make_crc32d16_n_21), .o(make_crc32d16_n_54) );
fflopd make_crc32d16_crc_reg_9_ ( .CK(newNet_115), .D(make_crc32d16_n_169), .Q(crc32_9_) );
XOR2_X1 make_crc32d16_g2211 ( .a(make_crc32d16_n_273), .b(d_7), .o(make_crc32d16_n_61) );
XOR2_X1 make_crc32d16_g2170 ( .a(make_crc32d16_n_62), .b(make_crc32d16_n_86), .o(make_crc32d16_n_99) );
XOR2_X1 make_crc32d16_g2241 ( .a(crc32_21_), .b(crc32_15_), .o(make_crc32d16_n_30) );
XOR2_X1 make_crc32d16_g2038 ( .a(make_crc32d16_n_160), .b(make_crc32d16_n_148), .o(make_crc32d16_n_171) );
XOR2_X1 make_crc32d16_g2151 ( .a(make_crc32d16_n_101), .b(make_crc32d16_n_47), .o(make_crc32d16_n_109) );
XOR2_X1 make_crc32d16_g2143 ( .a(make_crc32d16_n_111), .b(make_crc32d16_n_73), .o(make_crc32d16_n_115) );
XOR2_X1 make_crc32d16_g2178 ( .a(make_crc32d16_n_75), .b(make_crc32d16_n_7), .o(make_crc32d16_n_94) );
INV_Z1 g38 ( .a(crc32_31_), .o(crc32N_0) );
BUF_X2 newInst_75 ( .a(newNet_74), .o(newNet_75) );
BUF_X2 newInst_51 ( .a(newNet_24), .o(newNet_51) );
XOR2_X1 make_crc32d16_g2020 ( .a(make_crc32d16_n_170), .b(make_crc32d16_n_156), .o(make_crc32d16_n_185) );
BUF_X2 newInst_188 ( .a(newNet_187), .o(newNet_188) );
XOR2_X1 make_crc32d16_g2149 ( .a(make_crc32d16_n_101), .b(make_crc32d16_n_213), .o(make_crc32d16_n_111) );
XOR2_X1 make_crc32d16_g2061 ( .a(make_crc32d16_n_138), .b(make_crc32d16_n_197), .o(make_crc32d16_n_151) );
XOR2_X1 make_crc32d16_g2266 ( .a(make_crc32d16_n_201), .b(d_2), .o(make_crc32d16_n_4) );
BUF_X2 newInst_194 ( .a(newNet_193), .o(newNet_194) );
BUF_X2 newInst_112 ( .a(newNet_18), .o(newNet_112) );
BUF_X2 newInst_107 ( .a(newNet_106), .o(newNet_107) );
BUF_X2 newInst_183 ( .a(newNet_182), .o(newNet_183) );
XOR2_X1 make_crc32d16_g2025 ( .a(make_crc32d16_n_172), .b(make_crc32d16_n_149), .o(make_crc32d16_n_180) );
BUF_X2 newInst_161 ( .a(newNet_160), .o(newNet_161) );
BUF_X2 newInst_115 ( .a(newNet_83), .o(newNet_115) );
BUF_X2 newInst_139 ( .a(newNet_138), .o(newNet_139) );
BUF_X2 newInst_120 ( .a(newNet_119), .o(newNet_120) );
XOR2_X1 make_crc32d16_g2188 ( .a(make_crc32d16_n_54), .b(make_crc32d16_n_2), .o(make_crc32d16_n_84) );
XOR2_X1 make_crc32d16_g2104 ( .a(crc32_29_), .b(crc32_26_), .o(make_crc32d16_n_215) );
XOR2_X1 make_crc32d16_g2274 ( .a(crc32_18_), .b(d_13), .o(make_crc32d16_n_270) );
XOR2_X1 make_crc32d16_g2088 ( .a(crc32_25_), .b(crc32_24_), .o(make_crc32d16_n_219) );
XOR2_X1 make_crc32d16_g2219 ( .a(make_crc32d16_n_15), .b(make_crc32d16_n_45), .o(make_crc32d16_n_53) );
INV_Z1 g36 ( .a(crc32_7_), .o(crc32N_24) );
BUF_X2 newInst_148 ( .a(newNet_147), .o(newNet_148) );
fflopd make_crc32d16_crc_reg_30_ ( .CK(newNet_33), .D(make_crc32d16_n_98), .Q(crc32_30_) );
BUF_X2 newInst_22 ( .a(newNet_21), .o(newNet_22) );
BUF_X2 newInst_61 ( .a(newNet_60), .o(newNet_61) );
XOR2_X1 make_crc32d16_g2270 ( .a(make_crc32d16_n_216), .b(make_crc32d16_n_215), .o(make_crc32d16_n_1) );
XOR2_X1 make_crc32d16_g2242 ( .a(crc32_24_), .b(crc32_3_), .o(make_crc32d16_n_29) );
BUF_X2 newInst_95 ( .a(newNet_94), .o(newNet_95) );
BUF_X2 newInst_133 ( .a(newNet_132), .o(newNet_133) );
XOR2_X1 make_crc32d16_g2227 ( .a(crc32_17_), .b(d_10), .o(make_crc32d16_n_43) );
XOR2_X1 make_crc32d16_g2064 ( .a(make_crc32d16_n_134), .b(make_crc32d16_n_271), .o(make_crc32d16_n_150) );
XOR2_X1 make_crc32d16_g2069 ( .a(make_crc32d16_n_129), .b(make_crc32d16_n_197), .o(make_crc32d16_n_145) );
XOR2_X1 make_crc32d16_g2216 ( .a(make_crc32d16_n_25), .b(make_crc32d16_n_274), .o(make_crc32d16_n_56) );
BUF_X2 newInst_127 ( .a(newNet_126), .o(newNet_127) );
fflopd make_crc32d16_crc_reg_31_ ( .CK(newNet_98), .D(make_crc32d16_n_113), .Q(crc32_31_) );
XOR2_X1 make_crc32d16_g2047 ( .a(make_crc32d16_n_154), .b(make_crc32d16_n_197), .o(make_crc32d16_n_164) );
BUF_X2 newInst_144 ( .a(newNet_71), .o(newNet_144) );
fflopd make_crc32d16_crc_reg_25_ ( .CK(newNet_101), .D(make_crc32d16_n_115), .Q(crc32_25_) );
BUF_X2 newInst_41 ( .a(newNet_40), .o(newNet_41) );
BUF_X2 newInst_195 ( .a(newNet_194), .o(newNet_195) );
fflopd make_crc32d16_crc_reg_13_ ( .CK(newNet_125), .D(make_crc32d16_n_168), .Q(crc32_13_) );
XOR2_X1 make_crc32d16_g2112 ( .a(crc32_20_), .b(d_11), .o(make_crc32d16_n_122) );
XOR2_X1 make_crc32d16_g2252 ( .a(crc32_29_), .b(d_14), .o(make_crc32d16_n_16) );
BUF_X2 newInst_38 ( .a(newNet_37), .o(newNet_38) );
XOR2_X1 make_crc32d16_g2077 ( .a(make_crc32d16_n_132), .b(make_crc32d16_n_270), .o(make_crc32d16_n_136) );
XOR2_X1 make_crc32d16_g2234 ( .a(make_crc32d16_n_195), .b(crc32_24_), .o(make_crc32d16_n_36) );
BUF_X2 newInst_190 ( .a(newNet_189), .o(newNet_190) );
BUF_X2 newInst_94 ( .a(newNet_93), .o(newNet_94) );
BUF_X2 newInst_119 ( .a(newNet_118), .o(newNet_119) );
BUF_X2 newInst_35 ( .a(newNet_34), .o(newNet_35) );
fflopd make_crc32d16_crc_reg_15_ ( .CK(newNet_146), .D(make_crc32d16_n_188), .Q(crc32_15_) );
XOR2_X1 make_crc32d16_g2278 ( .a(crc32_28_), .b(d_3), .o(make_crc32d16_n_274) );
XOR2_X1 make_crc32d16_g2275 ( .a(crc32_26_), .b(d_5), .o(make_crc32d16_n_271) );
XOR2_X1 make_crc32d16_g2172 ( .a(make_crc32d16_n_93), .b(make_crc32d16_n_52), .o(make_crc32d16_n_97) );
fflopd make_crc32d16_crc_reg_5_ ( .CK(newNet_143), .D(make_crc32d16_n_185), .Q(crc32_5_) );
BUF_X2 newInst_155 ( .a(newNet_154), .o(newNet_155) );
INV_X2 newInst_46 ( .a(newNet_45), .o(newNet_46) );
XOR2_X1 make_crc32d16_g2090 ( .a(d_14), .b(d_9), .o(make_crc32d16_n_211) );
XOR2_X1 make_crc32d16_g2100 ( .a(crc32_24_), .b(crc32_23_), .o(make_crc32d16_n_217) );
XOR2_X1 make_crc32d16_g2264 ( .a(crc32_11_), .b(d_14), .o(make_crc32d16_n_5) );
BUF_X2 newInst_154 ( .a(newNet_153), .o(newNet_154) );
BUF_X2 newInst_198 ( .a(newNet_197), .o(newNet_198) );
XOR2_X1 make_crc32d16_g2094 ( .a(d_9), .b(d_8), .o(make_crc32d16_n_203) );
BUF_X2 newInst_31 ( .a(newNet_30), .o(newNet_31) );
XOR2_X1 make_crc32d16_g2167 ( .a(make_crc32d16_n_65), .b(make_crc32d16_n_89), .o(make_crc32d16_n_102) );
BUF_X2 newInst_72 ( .a(newNet_44), .o(newNet_72) );
INV_Z1 g48 ( .a(crc32_21_), .o(crc32N_10) );
fflopd make_crc32d16_crc_reg_14_ ( .CK(newNet_169), .D(make_crc32d16_n_180), .Q(crc32_14_) );
BUF_X2 newInst_126 ( .a(newNet_114), .o(newNet_126) );
XOR2_X1 make_crc32d16_g2198 ( .a(make_crc32d16_n_41), .b(make_crc32d16_n_26), .o(make_crc32d16_n_74) );
XOR2_X1 make_crc32d16_g2250 ( .a(make_crc32d16_n_208), .b(d_13), .o(make_crc32d16_n_17) );
XOR2_X1 make_crc32d16_g2212 ( .a(make_crc32d16_n_51), .b(crc32_13_), .o(make_crc32d16_n_60) );
XOR2_X1 make_crc32d16_g2110 ( .a(d_12), .b(d_11), .o(make_crc32d16_n_206) );
BUF_X2 newInst_130 ( .a(newNet_129), .o(newNet_130) );
fflopd make_crc32d16_crc_reg_1_ ( .CK(newNet_114), .D(make_crc32d16_n_175), .Q(crc32_1_) );
BUF_X2 newInst_166 ( .a(newNet_165), .o(newNet_166) );
BUF_X2 newInst_100 ( .a(newNet_99), .o(newNet_100) );
XOR2_X1 make_crc32d16_g2046 ( .a(make_crc32d16_n_155), .b(make_crc32d16_n_131), .o(make_crc32d16_n_165) );
INV_Z1 g53 ( .a(crc32_23_), .o(crc32N_8) );
BUF_X2 newInst_47 ( .a(newNet_46), .o(newNet_47) );
BUF_X2 newInst_147 ( .a(newNet_23), .o(newNet_147) );
BUF_X2 newInst_141 ( .a(newNet_140), .o(newNet_141) );
BUF_X2 newInst_92 ( .a(newNet_91), .o(newNet_92) );
BUF_X2 newInst_57 ( .a(newNet_56), .o(newNet_57) );
XOR2_X1 make_crc32d16_g2099 ( .a(d_9), .b(d_6), .o(make_crc32d16_n_194) );
XOR2_X1 make_crc32d16_g2144 ( .a(make_crc32d16_n_109), .b(make_crc32d16_n_66), .o(make_crc32d16_n_114) );
INV_Z1 g61 ( .a(crc32_28_), .o(crc32N_3) );
XOR2_X1 make_crc32d16_g2202 ( .a(make_crc32d16_n_270), .b(make_crc32d16_n_38), .o(make_crc32d16_n_70) );
fflopd make_crc32d16_crc_reg_22_ ( .CK(newNet_83), .D(make_crc32d16_n_96), .Q(crc32_22_) );
XOR2_X1 make_crc32d16_g2193 ( .a(make_crc32d16_n_197), .b(make_crc32d16_n_271), .o(make_crc32d16_n_79) );
XOR2_X1 make_crc32d16_g2260 ( .a(make_crc32d16_n_211), .b(make_crc32d16_n_256), .o(make_crc32d16_n_9) );
BUF_X2 newInst_199 ( .a(newNet_198), .o(newNet_199) );
XOR2_X1 make_crc32d16_g2041 ( .a(make_crc32d16_n_158), .b(make_crc32d16_n_154), .o(make_crc32d16_n_169) );
XOR2_X1 make_crc32d16_g2118 ( .a(crc32_19_), .b(crc32_18_), .o(make_crc32d16_n_213) );
BUF_X2 newInst_44 ( .a(newNet_43), .o(newNet_44) );
fflopd make_crc32d16_crc_reg_18_ ( .CK(newNet_50), .D(make_crc32d16_n_107), .Q(crc32_18_) );
XOR2_X1 make_crc32d16_g2206 ( .a(make_crc32d16_n_29), .b(make_crc32d16_n_269), .o(make_crc32d16_n_66) );
BUF_X2 newInst_174 ( .a(newNet_173), .o(newNet_174) );
INV_Z1 g64 ( .a(crc32_30_), .o(crc32N_1) );
BUF_X2 newInst_191 ( .a(newNet_190), .o(newNet_191) );
XOR2_X1 make_crc32d16_g2050 ( .a(make_crc32d16_n_151), .b(make_crc32d16_n_150), .o(make_crc32d16_n_159) );
BUF_X2 newInst_66 ( .a(newNet_65), .o(newNet_66) );
XOR2_X1 make_crc32d16_g2037 ( .a(make_crc32d16_n_163), .b(make_crc32d16_n_271), .o(make_crc32d16_n_179) );
XOR2_X1 make_crc32d16_g2184 ( .a(make_crc32d16_n_68), .b(make_crc32d16_n_79), .o(make_crc32d16_n_88) );
BUF_X2 newInst_40 ( .a(newNet_39), .o(newNet_40) );
XOR2_X1 make_crc32d16_g2269 ( .a(make_crc32d16_n_257), .b(crc32_0_), .o(make_crc32d16_n_2) );
BUF_X2 newInst_123 ( .a(newNet_122), .o(newNet_123) );
BUF_X2 newInst_99 ( .a(newNet_53), .o(newNet_99) );
BUF_X2 newInst_82 ( .a(newNet_81), .o(newNet_82) );
BUF_X2 newInst_152 ( .a(newNet_151), .o(newNet_152) );
XOR2_X1 make_crc32d16_g2177 ( .a(make_crc32d16_n_77), .b(make_crc32d16_n_10), .o(make_crc32d16_n_95) );
BUF_X2 newInst_78 ( .a(newNet_77), .o(newNet_78) );
BUF_X2 newInst_91 ( .a(newNet_49), .o(newNet_91) );
BUF_X2 newInst_118 ( .a(newNet_117), .o(newNet_118) );
BUF_X2 newInst_15 ( .a(newNet_14), .o(newNet_15) );
XOR2_X1 make_crc32d16_g2073 ( .a(make_crc32d16_n_130), .b(make_crc32d16_n_123), .o(make_crc32d16_n_139) );
BUF_X2 newInst_9 ( .a(newNet_8), .o(newNet_9) );
XOR2_X1 make_crc32d16_g2183 ( .a(make_crc32d16_n_64), .b(make_crc32d16_n_17), .o(make_crc32d16_n_89) );
BUF_X2 newInst_185 ( .a(newNet_184), .o(newNet_185) );
XOR2_X1 make_crc32d16_g2081 ( .a(crc32_25_), .b(crc32_22_), .o(make_crc32d16_n_209) );
BUF_X2 newInst_160 ( .a(newNet_140), .o(newNet_160) );
BUF_X2 newInst_189 ( .a(newNet_60), .o(newNet_189) );
INV_Z1 g50 ( .a(crc32_2_), .o(crc32N_29) );
BUF_X2 newInst_182 ( .a(newNet_181), .o(newNet_182) );
INV_Z1 g56 ( .a(crc32_25_), .o(crc32N_6) );

endmodule
